
module inputBuffer_1 ( clk, reset, polarity, sendIn, readyIn, dataIn, dataOut, 
        request, outputBufferGrant );
  input [63:0] dataIn;
  output [63:0] dataOut;
  output [1:0] request;
  input [1:0] outputBufferGrant;
  input clk, reset, polarity, sendIn;
  output readyIn;
  wire   n924, n925, evenBufferFull, oddBufferFull, n140, n141, n142, n143,
         n144, n145, n146, n147, n152, n153, n154, n155, n156, n157, n158,
         n159, n169, n177, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n148, n149, n150,
         n151, n160, n161, n162, n163, n164, n165, n166, n167, n168, n170,
         n171, n172, n173, n174, n175, n176, n178, n179, n180, n181, n182,
         n183, n184, n314, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923;
  wire   [63:0] evenBuffer;
  wire   [63:0] oddBuffer;
  wire   [7:1] sub_131_aco_carry;
  wire   [7:1] sub_111_aco_carry;

  DFFSR oddBufferFull_reg ( .D(n801), .CLK(clk), .R(n427), .S(1'b1), .Q(
        oddBufferFull) );
  DFFSR evenBufferFull_reg ( .D(n800), .CLK(clk), .R(n427), .S(1'b1), .Q(
        evenBufferFull) );
  DFFSR oddBuffer_reg_63_ ( .D(n799), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[63]) );
  DFFSR oddBuffer_reg_62_ ( .D(n798), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[62]) );
  DFFSR oddBuffer_reg_61_ ( .D(n797), .CLK(clk), .R(n427), .S(1'b1), .Q(
        oddBuffer[61]) );
  DFFSR oddBuffer_reg_60_ ( .D(n796), .CLK(clk), .R(n427), .S(1'b1), .Q(
        oddBuffer[60]) );
  DFFSR oddBuffer_reg_59_ ( .D(n795), .CLK(clk), .R(n426), .S(1'b1), .Q(
        oddBuffer[59]) );
  DFFSR oddBuffer_reg_58_ ( .D(n794), .CLK(clk), .R(n427), .S(1'b1), .Q(
        oddBuffer[58]) );
  DFFSR oddBuffer_reg_57_ ( .D(n793), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[57]) );
  DFFSR oddBuffer_reg_56_ ( .D(n792), .CLK(clk), .R(n426), .S(1'b1), .Q(
        oddBuffer[56]) );
  DFFSR oddBuffer_reg_55_ ( .D(n791), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[55]) );
  DFFSR oddBuffer_reg_54_ ( .D(n790), .CLK(clk), .R(n427), .S(1'b1), .Q(
        oddBuffer[54]) );
  DFFSR oddBuffer_reg_53_ ( .D(n789), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[53]) );
  DFFSR oddBuffer_reg_52_ ( .D(n788), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[52]) );
  DFFSR oddBuffer_reg_51_ ( .D(n787), .CLK(clk), .R(n426), .S(1'b1), .Q(
        oddBuffer[51]) );
  DFFSR oddBuffer_reg_50_ ( .D(n786), .CLK(clk), .R(n426), .S(1'b1), .Q(
        oddBuffer[50]) );
  DFFSR oddBuffer_reg_49_ ( .D(n785), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[49]) );
  DFFSR oddBuffer_reg_48_ ( .D(n784), .CLK(clk), .R(n426), .S(1'b1), .Q(
        oddBuffer[48]) );
  DFFSR oddBuffer_reg_47_ ( .D(n783), .CLK(clk), .R(n426), .S(1'b1), .Q(
        oddBuffer[47]) );
  DFFSR oddBuffer_reg_46_ ( .D(n782), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[46]) );
  DFFSR oddBuffer_reg_45_ ( .D(n781), .CLK(clk), .R(n427), .S(1'b1), .Q(
        oddBuffer[45]) );
  DFFSR oddBuffer_reg_44_ ( .D(n780), .CLK(clk), .R(n427), .S(1'b1), .Q(
        oddBuffer[44]) );
  DFFSR oddBuffer_reg_43_ ( .D(n779), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[43]) );
  DFFSR oddBuffer_reg_42_ ( .D(n778), .CLK(clk), .R(n427), .S(1'b1), .Q(
        oddBuffer[42]) );
  DFFSR oddBuffer_reg_41_ ( .D(n777), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[41]) );
  DFFSR oddBuffer_reg_40_ ( .D(n776), .CLK(clk), .R(n427), .S(1'b1), .Q(
        oddBuffer[40]) );
  DFFSR oddBuffer_reg_39_ ( .D(n775), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[39]) );
  DFFSR oddBuffer_reg_38_ ( .D(n774), .CLK(clk), .R(n427), .S(1'b1), .Q(
        oddBuffer[38]) );
  DFFSR oddBuffer_reg_37_ ( .D(n773), .CLK(clk), .R(n427), .S(1'b1), .Q(
        oddBuffer[37]) );
  DFFSR oddBuffer_reg_36_ ( .D(n772), .CLK(clk), .R(n427), .S(1'b1), .Q(
        oddBuffer[36]) );
  DFFSR oddBuffer_reg_35_ ( .D(n771), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[35]) );
  DFFSR oddBuffer_reg_34_ ( .D(n770), .CLK(clk), .R(n426), .S(1'b1), .Q(
        oddBuffer[34]) );
  DFFSR oddBuffer_reg_33_ ( .D(n769), .CLK(clk), .R(n427), .S(1'b1), .Q(
        oddBuffer[33]) );
  DFFSR oddBuffer_reg_32_ ( .D(n768), .CLK(clk), .R(n426), .S(1'b1), .Q(
        oddBuffer[32]) );
  DFFSR oddBuffer_reg_31_ ( .D(n767), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[31]) );
  DFFSR oddBuffer_reg_30_ ( .D(n766), .CLK(clk), .R(n427), .S(1'b1), .Q(
        oddBuffer[30]) );
  DFFSR oddBuffer_reg_29_ ( .D(n765), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[29]) );
  DFFSR oddBuffer_reg_28_ ( .D(n764), .CLK(clk), .R(n427), .S(1'b1), .Q(
        oddBuffer[28]) );
  DFFSR oddBuffer_reg_27_ ( .D(n763), .CLK(clk), .R(n426), .S(1'b1), .Q(
        oddBuffer[27]) );
  DFFSR oddBuffer_reg_26_ ( .D(n762), .CLK(clk), .R(n426), .S(1'b1), .Q(
        oddBuffer[26]) );
  DFFSR oddBuffer_reg_25_ ( .D(n761), .CLK(clk), .R(n426), .S(1'b1), .Q(
        oddBuffer[25]) );
  DFFSR oddBuffer_reg_24_ ( .D(n760), .CLK(clk), .R(n426), .S(1'b1), .Q(
        oddBuffer[24]) );
  DFFSR oddBuffer_reg_23_ ( .D(n759), .CLK(clk), .R(n427), .S(1'b1), .Q(
        oddBuffer[23]) );
  DFFSR oddBuffer_reg_22_ ( .D(n758), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[22]) );
  DFFSR oddBuffer_reg_21_ ( .D(n757), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[21]) );
  DFFSR oddBuffer_reg_20_ ( .D(n756), .CLK(clk), .R(n426), .S(1'b1), .Q(
        oddBuffer[20]) );
  DFFSR oddBuffer_reg_19_ ( .D(n755), .CLK(clk), .R(n426), .S(1'b1), .Q(
        oddBuffer[19]) );
  DFFSR oddBuffer_reg_18_ ( .D(n754), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[18]) );
  DFFSR oddBuffer_reg_17_ ( .D(n753), .CLK(clk), .R(n427), .S(1'b1), .Q(
        oddBuffer[17]) );
  DFFSR oddBuffer_reg_16_ ( .D(n752), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[16]) );
  DFFSR oddBuffer_reg_15_ ( .D(n751), .CLK(clk), .R(n426), .S(1'b1), .Q(
        oddBuffer[15]) );
  DFFSR oddBuffer_reg_14_ ( .D(n750), .CLK(clk), .R(n426), .S(1'b1), .Q(
        oddBuffer[14]) );
  DFFSR oddBuffer_reg_13_ ( .D(n749), .CLK(clk), .R(n427), .S(1'b1), .Q(
        oddBuffer[13]) );
  DFFSR oddBuffer_reg_12_ ( .D(n748), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[12]) );
  DFFSR oddBuffer_reg_11_ ( .D(n747), .CLK(clk), .R(n426), .S(1'b1), .Q(
        oddBuffer[11]) );
  DFFSR oddBuffer_reg_10_ ( .D(n746), .CLK(clk), .R(n427), .S(1'b1), .Q(
        oddBuffer[10]) );
  DFFSR oddBuffer_reg_9_ ( .D(n745), .CLK(clk), .R(n427), .S(1'b1), .Q(
        oddBuffer[9]) );
  DFFSR oddBuffer_reg_8_ ( .D(n744), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[8]) );
  DFFSR oddBuffer_reg_7_ ( .D(n743), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[7]) );
  DFFSR oddBuffer_reg_6_ ( .D(n742), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[6]) );
  DFFSR oddBuffer_reg_5_ ( .D(n741), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[5]) );
  DFFSR oddBuffer_reg_4_ ( .D(n740), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[4]) );
  DFFSR oddBuffer_reg_3_ ( .D(n739), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[3]) );
  DFFSR oddBuffer_reg_2_ ( .D(n738), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[2]) );
  DFFSR oddBuffer_reg_1_ ( .D(n737), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[1]) );
  DFFSR oddBuffer_reg_0_ ( .D(n736), .CLK(clk), .R(n428), .S(1'b1), .Q(
        oddBuffer[0]) );
  DFFSR evenBuffer_reg_63_ ( .D(n735), .CLK(clk), .R(n428), .S(1'b1), .Q(
        evenBuffer[63]) );
  DFFSR evenBuffer_reg_62_ ( .D(n734), .CLK(clk), .R(n428), .S(1'b1), .Q(
        evenBuffer[62]) );
  DFFSR evenBuffer_reg_61_ ( .D(n733), .CLK(clk), .R(n428), .S(1'b1), .Q(
        evenBuffer[61]) );
  DFFSR evenBuffer_reg_60_ ( .D(n732), .CLK(clk), .R(n428), .S(1'b1), .Q(
        evenBuffer[60]) );
  DFFSR evenBuffer_reg_59_ ( .D(n731), .CLK(clk), .R(n426), .S(1'b1), .Q(
        evenBuffer[59]) );
  DFFSR evenBuffer_reg_58_ ( .D(n730), .CLK(clk), .R(n427), .S(1'b1), .Q(
        evenBuffer[58]) );
  DFFSR evenBuffer_reg_57_ ( .D(n729), .CLK(clk), .R(n428), .S(1'b1), .Q(
        evenBuffer[57]) );
  DFFSR evenBuffer_reg_56_ ( .D(n728), .CLK(clk), .R(n427), .S(1'b1), .Q(
        evenBuffer[56]) );
  DFFSR evenBuffer_reg_55_ ( .D(n727), .CLK(clk), .R(n428), .S(1'b1), .Q(
        evenBuffer[55]) );
  DFFSR evenBuffer_reg_54_ ( .D(n726), .CLK(clk), .R(n426), .S(1'b1), .Q(
        evenBuffer[54]) );
  DFFSR evenBuffer_reg_53_ ( .D(n725), .CLK(clk), .R(n426), .S(1'b1), .Q(
        evenBuffer[53]) );
  DFFSR evenBuffer_reg_52_ ( .D(n724), .CLK(clk), .R(n427), .S(1'b1), .Q(
        evenBuffer[52]) );
  DFFSR evenBuffer_reg_51_ ( .D(n723), .CLK(clk), .R(n427), .S(1'b1), .Q(
        evenBuffer[51]) );
  DFFSR evenBuffer_reg_50_ ( .D(n722), .CLK(clk), .R(n428), .S(1'b1), .Q(
        evenBuffer[50]) );
  DFFSR evenBuffer_reg_49_ ( .D(n721), .CLK(clk), .R(n426), .S(1'b1), .Q(
        evenBuffer[49]) );
  DFFSR evenBuffer_reg_48_ ( .D(n720), .CLK(clk), .R(n428), .S(1'b1), .Q(
        evenBuffer[48]) );
  DFFSR evenBuffer_reg_47_ ( .D(n719), .CLK(clk), .R(n428), .S(1'b1), .Q(
        evenBuffer[47]) );
  DFFSR evenBuffer_reg_46_ ( .D(n718), .CLK(clk), .R(n426), .S(1'b1), .Q(
        evenBuffer[46]) );
  DFFSR evenBuffer_reg_45_ ( .D(n717), .CLK(clk), .R(n426), .S(1'b1), .Q(
        evenBuffer[45]) );
  DFFSR evenBuffer_reg_44_ ( .D(n716), .CLK(clk), .R(n426), .S(1'b1), .Q(
        evenBuffer[44]) );
  DFFSR evenBuffer_reg_43_ ( .D(n715), .CLK(clk), .R(n427), .S(1'b1), .Q(
        evenBuffer[43]) );
  DFFSR evenBuffer_reg_42_ ( .D(n714), .CLK(clk), .R(n428), .S(1'b1), .Q(
        evenBuffer[42]) );
  DFFSR evenBuffer_reg_41_ ( .D(n713), .CLK(clk), .R(n426), .S(1'b1), .Q(
        evenBuffer[41]) );
  DFFSR evenBuffer_reg_40_ ( .D(n712), .CLK(clk), .R(n426), .S(1'b1), .Q(
        evenBuffer[40]) );
  DFFSR evenBuffer_reg_39_ ( .D(n711), .CLK(clk), .R(n427), .S(1'b1), .Q(
        evenBuffer[39]) );
  DFFSR evenBuffer_reg_38_ ( .D(n710), .CLK(clk), .R(n426), .S(1'b1), .Q(
        evenBuffer[38]) );
  DFFSR evenBuffer_reg_37_ ( .D(n709), .CLK(clk), .R(n428), .S(1'b1), .Q(
        evenBuffer[37]) );
  DFFSR evenBuffer_reg_36_ ( .D(n708), .CLK(clk), .R(n427), .S(1'b1), .Q(
        evenBuffer[36]) );
  DFFSR evenBuffer_reg_35_ ( .D(n707), .CLK(clk), .R(n428), .S(1'b1), .Q(
        evenBuffer[35]) );
  DFFSR evenBuffer_reg_34_ ( .D(n706), .CLK(clk), .R(n426), .S(1'b1), .Q(
        evenBuffer[34]) );
  DFFSR evenBuffer_reg_33_ ( .D(n705), .CLK(clk), .R(n427), .S(1'b1), .Q(
        evenBuffer[33]) );
  DFFSR evenBuffer_reg_32_ ( .D(n704), .CLK(clk), .R(n428), .S(1'b1), .Q(
        evenBuffer[32]) );
  DFFSR evenBuffer_reg_31_ ( .D(n703), .CLK(clk), .R(n426), .S(1'b1), .Q(
        evenBuffer[31]) );
  DFFSR evenBuffer_reg_30_ ( .D(n702), .CLK(clk), .R(n427), .S(1'b1), .Q(
        evenBuffer[30]) );
  DFFSR evenBuffer_reg_29_ ( .D(n701), .CLK(clk), .R(n428), .S(1'b1), .Q(
        evenBuffer[29]) );
  DFFSR evenBuffer_reg_28_ ( .D(n700), .CLK(clk), .R(n426), .S(1'b1), .Q(
        evenBuffer[28]) );
  DFFSR evenBuffer_reg_27_ ( .D(n699), .CLK(clk), .R(n427), .S(1'b1), .Q(
        evenBuffer[27]) );
  DFFSR evenBuffer_reg_26_ ( .D(n698), .CLK(clk), .R(n426), .S(1'b1), .Q(
        evenBuffer[26]) );
  DFFSR evenBuffer_reg_25_ ( .D(n697), .CLK(clk), .R(n427), .S(1'b1), .Q(
        evenBuffer[25]) );
  DFFSR evenBuffer_reg_24_ ( .D(n696), .CLK(clk), .R(n428), .S(1'b1), .Q(
        evenBuffer[24]) );
  DFFSR evenBuffer_reg_23_ ( .D(n695), .CLK(clk), .R(n427), .S(1'b1), .Q(
        evenBuffer[23]) );
  DFFSR evenBuffer_reg_22_ ( .D(n694), .CLK(clk), .R(n427), .S(1'b1), .Q(
        evenBuffer[22]) );
  DFFSR evenBuffer_reg_21_ ( .D(n693), .CLK(clk), .R(n427), .S(1'b1), .Q(
        evenBuffer[21]) );
  DFFSR evenBuffer_reg_20_ ( .D(n692), .CLK(clk), .R(n427), .S(1'b1), .Q(
        evenBuffer[20]) );
  DFFSR evenBuffer_reg_19_ ( .D(n691), .CLK(clk), .R(n427), .S(1'b1), .Q(
        evenBuffer[19]) );
  DFFSR evenBuffer_reg_18_ ( .D(n690), .CLK(clk), .R(n427), .S(1'b1), .Q(
        evenBuffer[18]) );
  DFFSR evenBuffer_reg_17_ ( .D(n689), .CLK(clk), .R(n427), .S(1'b1), .Q(
        evenBuffer[17]) );
  DFFSR evenBuffer_reg_16_ ( .D(n688), .CLK(clk), .R(n427), .S(1'b1), .Q(
        evenBuffer[16]) );
  DFFSR evenBuffer_reg_15_ ( .D(n687), .CLK(clk), .R(n427), .S(1'b1), .Q(
        evenBuffer[15]) );
  DFFSR evenBuffer_reg_14_ ( .D(n686), .CLK(clk), .R(n427), .S(1'b1), .Q(
        evenBuffer[14]) );
  DFFSR evenBuffer_reg_13_ ( .D(n685), .CLK(clk), .R(n427), .S(1'b1), .Q(
        evenBuffer[13]) );
  DFFSR evenBuffer_reg_12_ ( .D(n684), .CLK(clk), .R(n427), .S(1'b1), .Q(
        evenBuffer[12]) );
  DFFSR evenBuffer_reg_11_ ( .D(n683), .CLK(clk), .R(n426), .S(1'b1), .Q(
        evenBuffer[11]) );
  DFFSR evenBuffer_reg_10_ ( .D(n682), .CLK(clk), .R(n426), .S(1'b1), .Q(
        evenBuffer[10]) );
  DFFSR evenBuffer_reg_9_ ( .D(n681), .CLK(clk), .R(n426), .S(1'b1), .Q(
        evenBuffer[9]) );
  DFFSR evenBuffer_reg_8_ ( .D(n680), .CLK(clk), .R(n426), .S(1'b1), .Q(
        evenBuffer[8]) );
  DFFSR evenBuffer_reg_7_ ( .D(n679), .CLK(clk), .R(n426), .S(1'b1), .Q(
        evenBuffer[7]) );
  DFFSR evenBuffer_reg_6_ ( .D(n678), .CLK(clk), .R(n426), .S(1'b1), .Q(
        evenBuffer[6]) );
  DFFSR evenBuffer_reg_5_ ( .D(n677), .CLK(clk), .R(n426), .S(1'b1), .Q(
        evenBuffer[5]) );
  DFFSR evenBuffer_reg_4_ ( .D(n676), .CLK(clk), .R(n426), .S(1'b1), .Q(
        evenBuffer[4]) );
  DFFSR evenBuffer_reg_3_ ( .D(n675), .CLK(clk), .R(n426), .S(1'b1), .Q(
        evenBuffer[3]) );
  DFFSR evenBuffer_reg_2_ ( .D(n674), .CLK(clk), .R(n426), .S(1'b1), .Q(
        evenBuffer[2]) );
  DFFSR evenBuffer_reg_1_ ( .D(n673), .CLK(clk), .R(n426), .S(1'b1), .Q(
        evenBuffer[1]) );
  DFFSR evenBuffer_reg_0_ ( .D(n672), .CLK(clk), .R(n426), .S(1'b1), .Q(
        evenBuffer[0]) );
  NAND3X1 U281 ( .A(n169), .B(n440), .C(n418), .Y(n461) );
  NAND3X1 U282 ( .A(n353), .B(n177), .C(n432), .Y(n460) );
  NAND3X1 U284 ( .A(n179), .B(n441), .C(n418), .Y(n463) );
  NAND3X1 U285 ( .A(n353), .B(n322), .C(n432), .Y(n462) );
  NOR2X1 U286 ( .A(reset), .B(n77), .Y(readyIn) );
  AOI22X1 U287 ( .A(n432), .B(n452), .C(n451), .D(n442), .Y(n464) );
  OAI21X1 U288 ( .A(n465), .B(n922), .C(n337), .Y(n672) );
  OAI21X1 U290 ( .A(n465), .B(n921), .C(n325), .Y(n673) );
  OAI21X1 U292 ( .A(n465), .B(n920), .C(n184), .Y(n674) );
  OAI21X1 U294 ( .A(n465), .B(n919), .C(n171), .Y(n675) );
  OAI21X1 U296 ( .A(n465), .B(n918), .C(n160), .Y(n676) );
  OAI21X1 U298 ( .A(n465), .B(n917), .C(n134), .Y(n677) );
  OAI21X1 U300 ( .A(n465), .B(n916), .C(n124), .Y(n678) );
  OAI21X1 U302 ( .A(n465), .B(n915), .C(n114), .Y(n679) );
  OAI21X1 U304 ( .A(n465), .B(n914), .C(n104), .Y(n680) );
  OAI21X1 U306 ( .A(n465), .B(n913), .C(n95), .Y(n681) );
  OAI21X1 U308 ( .A(n465), .B(n912), .C(n87), .Y(n682) );
  OAI21X1 U310 ( .A(n465), .B(n911), .C(n76), .Y(n683) );
  OAI21X1 U312 ( .A(n465), .B(n910), .C(n336), .Y(n684) );
  OAI21X1 U314 ( .A(n465), .B(n909), .C(n324), .Y(n685) );
  OAI21X1 U316 ( .A(n465), .B(n908), .C(n75), .Y(n686) );
  OAI21X1 U318 ( .A(n465), .B(n907), .C(n183), .Y(n687) );
  OAI21X1 U320 ( .A(n465), .B(n906), .C(n170), .Y(n688) );
  OAI21X1 U322 ( .A(n465), .B(n905), .C(n151), .Y(n689) );
  OAI21X1 U324 ( .A(n465), .B(n904), .C(n133), .Y(n690) );
  OAI21X1 U326 ( .A(n465), .B(n903), .C(n123), .Y(n691) );
  OAI21X1 U328 ( .A(n465), .B(n902), .C(n113), .Y(n692) );
  OAI21X1 U330 ( .A(n465), .B(n901), .C(n103), .Y(n693) );
  OAI21X1 U332 ( .A(n465), .B(n900), .C(n94), .Y(n694) );
  OAI21X1 U334 ( .A(n465), .B(n899), .C(n86), .Y(n695) );
  OAI21X1 U336 ( .A(n465), .B(n898), .C(n74), .Y(n696) );
  OAI21X1 U338 ( .A(n465), .B(n897), .C(n335), .Y(n697) );
  OAI21X1 U340 ( .A(n465), .B(n896), .C(n73), .Y(n698) );
  OAI21X1 U342 ( .A(n465), .B(n895), .C(n182), .Y(n699) );
  OAI21X1 U344 ( .A(n465), .B(n894), .C(n168), .Y(n700) );
  OAI21X1 U346 ( .A(n465), .B(n893), .C(n150), .Y(n701) );
  OAI21X1 U348 ( .A(n465), .B(n892), .C(n132), .Y(n702) );
  OAI21X1 U350 ( .A(n465), .B(n891), .C(n122), .Y(n703) );
  OAI21X1 U352 ( .A(n465), .B(n890), .C(n112), .Y(n704) );
  OAI21X1 U354 ( .A(n465), .B(n889), .C(n102), .Y(n705) );
  OAI21X1 U356 ( .A(n465), .B(n888), .C(n93), .Y(n706) );
  OAI21X1 U358 ( .A(n465), .B(n887), .C(n85), .Y(n707) );
  OAI21X1 U360 ( .A(n465), .B(n886), .C(n72), .Y(n708) );
  OAI21X1 U362 ( .A(n465), .B(n885), .C(n71), .Y(n709) );
  OAI21X1 U364 ( .A(n465), .B(n884), .C(n70), .Y(n710) );
  OAI21X1 U366 ( .A(n465), .B(n883), .C(n181), .Y(n711) );
  OAI21X1 U368 ( .A(n465), .B(n882), .C(n167), .Y(n712) );
  OAI21X1 U370 ( .A(n465), .B(n881), .C(n149), .Y(n713) );
  OAI21X1 U372 ( .A(n465), .B(n880), .C(n131), .Y(n714) );
  OAI21X1 U374 ( .A(n465), .B(n879), .C(n121), .Y(n715) );
  OAI21X1 U376 ( .A(n465), .B(n878), .C(n111), .Y(n716) );
  OAI21X1 U378 ( .A(n465), .B(n877), .C(n101), .Y(n717) );
  OAI21X1 U380 ( .A(n465), .B(n876), .C(n92), .Y(n718) );
  OAI21X1 U382 ( .A(n465), .B(n875), .C(n84), .Y(n719) );
  OAI21X1 U384 ( .A(n465), .B(n874), .C(n343), .Y(n720) );
  OAI21X1 U386 ( .A(n465), .B(n873), .C(n332), .Y(n721) );
  OAI21X1 U388 ( .A(n465), .B(n872), .C(n69), .Y(n722) );
  OAI21X1 U390 ( .A(n465), .B(n871), .C(n68), .Y(n723) );
  OAI21X1 U392 ( .A(n465), .B(n870), .C(n331), .Y(n724) );
  OAI21X1 U394 ( .A(n465), .B(n869), .C(n320), .Y(n725) );
  OAI21X1 U396 ( .A(n465), .B(n868), .C(n148), .Y(n726) );
  OAI21X1 U398 ( .A(n465), .B(n867), .C(n130), .Y(n727) );
  OAI21X1 U400 ( .A(n465), .B(n866), .C(n166), .Y(n728) );
  OAI21X1 U402 ( .A(n465), .B(n865), .C(n120), .Y(n729) );
  OAI21X1 U404 ( .A(n465), .B(n864), .C(n110), .Y(n730) );
  OAI21X1 U406 ( .A(n465), .B(n863), .C(n100), .Y(n731) );
  OAI21X1 U408 ( .A(n465), .B(n862), .C(n91), .Y(n732) );
  OAI21X1 U410 ( .A(n465), .B(n861), .C(n83), .Y(n733) );
  OAI21X1 U412 ( .A(n465), .B(n860), .C(n67), .Y(n734) );
  OAI21X1 U414 ( .A(n465), .B(n859), .C(n66), .Y(n735) );
  OAI21X1 U416 ( .A(n531), .B(n858), .C(n350), .Y(n736) );
  OAI21X1 U418 ( .A(n531), .B(n857), .C(n342), .Y(n737) );
  OAI21X1 U420 ( .A(n531), .B(n856), .C(n330), .Y(n738) );
  OAI21X1 U422 ( .A(n531), .B(n855), .C(n319), .Y(n739) );
  OAI21X1 U424 ( .A(n531), .B(n854), .C(n349), .Y(n740) );
  OAI21X1 U426 ( .A(n531), .B(n853), .C(n176), .Y(n741) );
  OAI21X1 U428 ( .A(n531), .B(n852), .C(n165), .Y(n742) );
  OAI21X1 U430 ( .A(n531), .B(n851), .C(n139), .Y(n743) );
  OAI21X1 U432 ( .A(n531), .B(n850), .C(n129), .Y(n744) );
  OAI21X1 U434 ( .A(n531), .B(n849), .C(n119), .Y(n745) );
  OAI21X1 U436 ( .A(n531), .B(n848), .C(n109), .Y(n746) );
  OAI21X1 U438 ( .A(n531), .B(n847), .C(n99), .Y(n747) );
  OAI21X1 U440 ( .A(n531), .B(n846), .C(n90), .Y(n748) );
  OAI21X1 U442 ( .A(n531), .B(n845), .C(n341), .Y(n749) );
  OAI21X1 U444 ( .A(n531), .B(n844), .C(n65), .Y(n750) );
  OAI21X1 U446 ( .A(n531), .B(n843), .C(n329), .Y(n751) );
  OAI21X1 U448 ( .A(n531), .B(n842), .C(n348), .Y(n752) );
  OAI21X1 U450 ( .A(n531), .B(n841), .C(n318), .Y(n753) );
  OAI21X1 U452 ( .A(n531), .B(n840), .C(n175), .Y(n754) );
  OAI21X1 U454 ( .A(n531), .B(n839), .C(n164), .Y(n755) );
  OAI21X1 U456 ( .A(n531), .B(n838), .C(n138), .Y(n756) );
  OAI21X1 U458 ( .A(n531), .B(n837), .C(n128), .Y(n757) );
  OAI21X1 U460 ( .A(n531), .B(n836), .C(n118), .Y(n758) );
  OAI21X1 U462 ( .A(n531), .B(n835), .C(n108), .Y(n759) );
  OAI21X1 U464 ( .A(n531), .B(n834), .C(n98), .Y(n760) );
  OAI21X1 U466 ( .A(n531), .B(n833), .C(n89), .Y(n761) );
  OAI21X1 U468 ( .A(n531), .B(n832), .C(n64), .Y(n762) );
  OAI21X1 U470 ( .A(n531), .B(n831), .C(n340), .Y(n763) );
  OAI21X1 U472 ( .A(n531), .B(n830), .C(n347), .Y(n764) );
  OAI21X1 U474 ( .A(n531), .B(n829), .C(n328), .Y(n765) );
  OAI21X1 U476 ( .A(n531), .B(n828), .C(n317), .Y(n766) );
  OAI21X1 U478 ( .A(n531), .B(n827), .C(n174), .Y(n767) );
  OAI21X1 U480 ( .A(n531), .B(n826), .C(n163), .Y(n768) );
  OAI21X1 U482 ( .A(n531), .B(n825), .C(n137), .Y(n769) );
  OAI21X1 U484 ( .A(n531), .B(n824), .C(n127), .Y(n770) );
  OAI21X1 U486 ( .A(n531), .B(n823), .C(n117), .Y(n771) );
  OAI21X1 U488 ( .A(n531), .B(n822), .C(n107), .Y(n772) );
  OAI21X1 U490 ( .A(n531), .B(n821), .C(n97), .Y(n773) );
  OAI21X1 U492 ( .A(n531), .B(n820), .C(n88), .Y(n774) );
  OAI21X1 U494 ( .A(n531), .B(n819), .C(n339), .Y(n775) );
  OAI21X1 U496 ( .A(n531), .B(n818), .C(n346), .Y(n776) );
  OAI21X1 U498 ( .A(n531), .B(n817), .C(n327), .Y(n777) );
  OAI21X1 U500 ( .A(n531), .B(n816), .C(n316), .Y(n778) );
  OAI21X1 U502 ( .A(n531), .B(n815), .C(n173), .Y(n779) );
  OAI21X1 U504 ( .A(n531), .B(n814), .C(n162), .Y(n780) );
  OAI21X1 U506 ( .A(n531), .B(n813), .C(n136), .Y(n781) );
  OAI21X1 U508 ( .A(n531), .B(n812), .C(n126), .Y(n782) );
  OAI21X1 U510 ( .A(n531), .B(n811), .C(n116), .Y(n783) );
  OAI21X1 U512 ( .A(n531), .B(n810), .C(n106), .Y(n784) );
  OAI21X1 U514 ( .A(n531), .B(n809), .C(n63), .Y(n785) );
  OAI21X1 U516 ( .A(n531), .B(n808), .C(n82), .Y(n786) );
  OAI21X1 U518 ( .A(n531), .B(n807), .C(n62), .Y(n787) );
  OAI21X1 U520 ( .A(n531), .B(n806), .C(n96), .Y(n788) );
  OAI21X1 U522 ( .A(n531), .B(n805), .C(n326), .Y(n789) );
  OAI21X1 U524 ( .A(n531), .B(n804), .C(n81), .Y(n790) );
  OAI21X1 U526 ( .A(n531), .B(n803), .C(n61), .Y(n791) );
  OAI21X1 U528 ( .A(n531), .B(n802), .C(n338), .Y(n792) );
  OAI21X1 U530 ( .A(n531), .B(n459), .C(n314), .Y(n793) );
  OAI21X1 U532 ( .A(n531), .B(n458), .C(n172), .Y(n794) );
  OAI21X1 U534 ( .A(n531), .B(n457), .C(n161), .Y(n795) );
  OAI21X1 U536 ( .A(n531), .B(n456), .C(n135), .Y(n796) );
  OAI21X1 U538 ( .A(n531), .B(n455), .C(n125), .Y(n797) );
  OAI21X1 U540 ( .A(n531), .B(n454), .C(n115), .Y(n798) );
  OAI21X1 U542 ( .A(n531), .B(n453), .C(n105), .Y(n799) );
  OAI21X1 U544 ( .A(n452), .B(n465), .C(n351), .Y(n800) );
  OAI21X1 U546 ( .A(n432), .B(n78), .C(n359), .Y(n465) );
  OAI21X1 U548 ( .A(n451), .B(n531), .C(n360), .Y(n801) );
  OAI21X1 U550 ( .A(n432), .B(n923), .C(n599), .Y(n531) );
  NOR3X1 U553 ( .A(n323), .B(n344), .C(n422), .Y(n601) );
  NOR3X1 U555 ( .A(n178), .B(n333), .C(n357), .Y(n600) );
  NOR3X1 U558 ( .A(n180), .B(n334), .C(n358), .Y(n605) );
  NOR3X1 U560 ( .A(n321), .B(n345), .C(n423), .Y(n604) );
  OAI21X1 U562 ( .A(n433), .B(n913), .C(n60), .Y(dataOut[9]) );
  OAI21X1 U564 ( .A(n433), .B(n914), .C(n59), .Y(dataOut[8]) );
  OAI21X1 U566 ( .A(n433), .B(n915), .C(n58), .Y(dataOut[7]) );
  OAI21X1 U568 ( .A(n433), .B(n916), .C(n57), .Y(dataOut[6]) );
  OAI21X1 U570 ( .A(n433), .B(n859), .C(n56), .Y(dataOut[63]) );
  OAI21X1 U572 ( .A(n433), .B(n860), .C(n55), .Y(dataOut[62]) );
  OAI21X1 U574 ( .A(n433), .B(n861), .C(n54), .Y(dataOut[61]) );
  OAI21X1 U576 ( .A(n433), .B(n862), .C(n53), .Y(dataOut[60]) );
  OAI21X1 U578 ( .A(n433), .B(n917), .C(n52), .Y(dataOut[5]) );
  OAI21X1 U580 ( .A(n433), .B(n863), .C(n51), .Y(dataOut[59]) );
  OAI21X1 U582 ( .A(n434), .B(n864), .C(n50), .Y(dataOut[58]) );
  OAI21X1 U584 ( .A(n434), .B(n865), .C(n49), .Y(dataOut[57]) );
  OAI21X1 U586 ( .A(n434), .B(n866), .C(n48), .Y(dataOut[56]) );
  AOI22X1 U588 ( .A(n147), .B(n442), .C(n159), .D(n432), .Y(n621) );
  AOI22X1 U589 ( .A(n146), .B(n442), .C(n158), .D(n432), .Y(n622) );
  AOI22X1 U590 ( .A(n145), .B(n442), .C(n157), .D(n432), .Y(n623) );
  AOI22X1 U591 ( .A(n144), .B(n442), .C(n156), .D(n432), .Y(n624) );
  AOI22X1 U592 ( .A(n143), .B(n442), .C(n155), .D(n432), .Y(n625) );
  AOI22X1 U593 ( .A(n142), .B(n442), .C(n154), .D(n432), .Y(n626) );
  OAI21X1 U594 ( .A(n434), .B(n918), .C(n47), .Y(dataOut[4]) );
  AOI22X1 U596 ( .A(n141), .B(n442), .C(n153), .D(n432), .Y(n628) );
  AOI22X1 U597 ( .A(n140), .B(n442), .C(n152), .D(n432), .Y(n629) );
  OAI21X1 U598 ( .A(n434), .B(n875), .C(n46), .Y(dataOut[47]) );
  OAI21X1 U600 ( .A(n435), .B(n876), .C(n45), .Y(dataOut[46]) );
  OAI21X1 U602 ( .A(n435), .B(n877), .C(n44), .Y(dataOut[45]) );
  OAI21X1 U604 ( .A(n434), .B(n878), .C(n43), .Y(dataOut[44]) );
  OAI21X1 U606 ( .A(n435), .B(n879), .C(n42), .Y(dataOut[43]) );
  OAI21X1 U608 ( .A(n435), .B(n880), .C(n41), .Y(dataOut[42]) );
  OAI21X1 U610 ( .A(n435), .B(n881), .C(n40), .Y(dataOut[41]) );
  OAI21X1 U612 ( .A(n435), .B(n882), .C(n39), .Y(dataOut[40]) );
  OAI21X1 U614 ( .A(n435), .B(n919), .C(n38), .Y(dataOut[3]) );
  OAI21X1 U616 ( .A(n435), .B(n883), .C(n37), .Y(dataOut[39]) );
  OAI21X1 U618 ( .A(n436), .B(n884), .C(n36), .Y(dataOut[38]) );
  OAI21X1 U620 ( .A(n436), .B(n885), .C(n35), .Y(dataOut[37]) );
  OAI21X1 U622 ( .A(n435), .B(n886), .C(n34), .Y(dataOut[36]) );
  OAI21X1 U624 ( .A(n436), .B(n887), .C(n33), .Y(dataOut[35]) );
  OAI21X1 U626 ( .A(n436), .B(n888), .C(n32), .Y(dataOut[34]) );
  OAI21X1 U628 ( .A(n436), .B(n889), .C(n31), .Y(dataOut[33]) );
  OAI21X1 U630 ( .A(n436), .B(n890), .C(n30), .Y(dataOut[32]) );
  OAI21X1 U632 ( .A(n436), .B(n891), .C(n29), .Y(dataOut[31]) );
  OAI21X1 U634 ( .A(n436), .B(n892), .C(n28), .Y(dataOut[30]) );
  OAI21X1 U636 ( .A(n437), .B(n920), .C(n27), .Y(dataOut[2]) );
  OAI21X1 U638 ( .A(n437), .B(n893), .C(n26), .Y(dataOut[29]) );
  OAI21X1 U640 ( .A(n436), .B(n894), .C(n25), .Y(dataOut[28]) );
  OAI21X1 U642 ( .A(n437), .B(n895), .C(n24), .Y(dataOut[27]) );
  OAI21X1 U644 ( .A(n435), .B(n896), .C(n23), .Y(dataOut[26]) );
  OAI21X1 U646 ( .A(n437), .B(n897), .C(n22), .Y(dataOut[25]) );
  OAI21X1 U648 ( .A(n436), .B(n898), .C(n21), .Y(dataOut[24]) );
  OAI21X1 U650 ( .A(n436), .B(n899), .C(n20), .Y(dataOut[23]) );
  OAI21X1 U652 ( .A(n435), .B(n900), .C(n19), .Y(dataOut[22]) );
  OAI21X1 U654 ( .A(n436), .B(n901), .C(n18), .Y(dataOut[21]) );
  OAI21X1 U656 ( .A(n435), .B(n902), .C(n17), .Y(dataOut[20]) );
  OAI21X1 U658 ( .A(n436), .B(n921), .C(n16), .Y(dataOut[1]) );
  OAI21X1 U660 ( .A(n435), .B(n903), .C(n15), .Y(dataOut[19]) );
  OAI21X1 U662 ( .A(n434), .B(n904), .C(n14), .Y(dataOut[18]) );
  OAI21X1 U664 ( .A(n434), .B(n905), .C(n13), .Y(dataOut[17]) );
  OAI21X1 U666 ( .A(n434), .B(n906), .C(n12), .Y(dataOut[16]) );
  OAI21X1 U668 ( .A(n434), .B(n907), .C(n11), .Y(dataOut[15]) );
  OAI21X1 U670 ( .A(n434), .B(n908), .C(n10), .Y(dataOut[14]) );
  OAI21X1 U672 ( .A(n434), .B(n909), .C(n9), .Y(dataOut[13]) );
  OAI21X1 U674 ( .A(n433), .B(n910), .C(n8), .Y(dataOut[12]) );
  OAI21X1 U676 ( .A(n434), .B(n911), .C(n7), .Y(dataOut[11]) );
  OAI21X1 U678 ( .A(n433), .B(n912), .C(n6), .Y(dataOut[10]) );
  OAI21X1 U680 ( .A(n433), .B(n922), .C(n5), .Y(dataOut[0]) );
  AND2X1 U4 ( .A(n2), .B(n4), .Y(n924) );
  OR2X1 U5 ( .A(n169), .B(n423), .Y(sub_111_aco_carry[1]) );
  OR2X1 U133 ( .A(n177), .B(n357), .Y(sub_131_aco_carry[1]) );
  OR2X1 U135 ( .A(sub_111_aco_carry[1]), .B(n345), .Y(sub_111_aco_carry[2]) );
  OR2X1 U136 ( .A(sub_131_aco_carry[1]), .B(n333), .Y(sub_131_aco_carry[2]) );
  OR2X1 U137 ( .A(sub_111_aco_carry[2]), .B(n421), .Y(sub_111_aco_carry[3]) );
  OR2X1 U138 ( .A(sub_131_aco_carry[2]), .B(n356), .Y(sub_131_aco_carry[3]) );
  OR2X1 U139 ( .A(sub_111_aco_carry[3]), .B(n420), .Y(sub_111_aco_carry[4]) );
  OR2X1 U140 ( .A(sub_131_aco_carry[3]), .B(n355), .Y(sub_131_aco_carry[4]) );
  OR2X1 U141 ( .A(sub_111_aco_carry[4]), .B(n358), .Y(sub_111_aco_carry[5]) );
  OR2X1 U142 ( .A(sub_131_aco_carry[4]), .B(n422), .Y(sub_131_aco_carry[5]) );
  OR2X1 U143 ( .A(sub_111_aco_carry[5]), .B(n334), .Y(sub_111_aco_carry[6]) );
  OR2X1 U144 ( .A(sub_131_aco_carry[5]), .B(n344), .Y(sub_131_aco_carry[6]) );
  OR2X1 U145 ( .A(sub_111_aco_carry[6]), .B(n419), .Y(sub_111_aco_carry[7]) );
  OR2X1 U146 ( .A(sub_131_aco_carry[6]), .B(n354), .Y(sub_131_aco_carry[7]) );
  AND2X1 U147 ( .A(n1), .B(n3), .Y(n925) );
  OR2X1 U148 ( .A(n442), .B(n78), .Y(n599) );
  BUFX2 U149 ( .A(n462), .Y(n1) );
  BUFX2 U150 ( .A(n460), .Y(n2) );
  BUFX2 U151 ( .A(n463), .Y(n3) );
  BUFX2 U152 ( .A(n461), .Y(n4) );
  AND2X1 U153 ( .A(n416), .B(n438), .Y(n671) );
  INVX1 U154 ( .A(n671), .Y(n5) );
  AND2X1 U155 ( .A(n406), .B(n437), .Y(n670) );
  INVX1 U156 ( .A(n670), .Y(n6) );
  AND2X1 U157 ( .A(n405), .B(n437), .Y(n669) );
  INVX1 U158 ( .A(n669), .Y(n7) );
  AND2X1 U159 ( .A(n404), .B(n437), .Y(n668) );
  INVX1 U160 ( .A(n668), .Y(n8) );
  AND2X1 U161 ( .A(n403), .B(n437), .Y(n667) );
  INVX1 U162 ( .A(n667), .Y(n9) );
  AND2X1 U163 ( .A(n402), .B(n437), .Y(n666) );
  INVX1 U164 ( .A(n666), .Y(n10) );
  AND2X1 U165 ( .A(n401), .B(n437), .Y(n665) );
  INVX1 U166 ( .A(n665), .Y(n11) );
  AND2X1 U167 ( .A(n400), .B(n438), .Y(n664) );
  INVX1 U168 ( .A(n664), .Y(n12) );
  AND2X1 U169 ( .A(n399), .B(n438), .Y(n663) );
  INVX1 U170 ( .A(n663), .Y(n13) );
  AND2X1 U171 ( .A(n398), .B(n437), .Y(n662) );
  INVX1 U172 ( .A(n662), .Y(n14) );
  AND2X1 U173 ( .A(n397), .B(n437), .Y(n661) );
  INVX1 U174 ( .A(n661), .Y(n15) );
  AND2X1 U175 ( .A(n415), .B(n438), .Y(n660) );
  INVX1 U176 ( .A(n660), .Y(n16) );
  AND2X1 U177 ( .A(n396), .B(n437), .Y(n659) );
  INVX1 U178 ( .A(n659), .Y(n17) );
  AND2X1 U179 ( .A(n395), .B(n437), .Y(n658) );
  INVX1 U180 ( .A(n658), .Y(n18) );
  AND2X1 U181 ( .A(n394), .B(n438), .Y(n657) );
  INVX1 U182 ( .A(n657), .Y(n19) );
  AND2X1 U183 ( .A(n393), .B(n437), .Y(n656) );
  INVX1 U184 ( .A(n656), .Y(n20) );
  AND2X1 U185 ( .A(n392), .B(n438), .Y(n655) );
  INVX1 U186 ( .A(n655), .Y(n21) );
  AND2X1 U187 ( .A(n391), .B(n438), .Y(n654) );
  INVX1 U188 ( .A(n654), .Y(n22) );
  AND2X1 U189 ( .A(n390), .B(n438), .Y(n653) );
  INVX1 U190 ( .A(n653), .Y(n23) );
  AND2X1 U191 ( .A(n389), .B(n438), .Y(n652) );
  INVX1 U192 ( .A(n652), .Y(n24) );
  AND2X1 U193 ( .A(n388), .B(n438), .Y(n651) );
  INVX1 U194 ( .A(n651), .Y(n25) );
  AND2X1 U195 ( .A(n387), .B(n438), .Y(n650) );
  INVX1 U196 ( .A(n650), .Y(n26) );
  AND2X1 U197 ( .A(n414), .B(n438), .Y(n649) );
  INVX1 U198 ( .A(n649), .Y(n27) );
  AND2X1 U199 ( .A(n386), .B(n438), .Y(n648) );
  INVX1 U200 ( .A(n648), .Y(n28) );
  AND2X1 U201 ( .A(n385), .B(n438), .Y(n647) );
  INVX1 U202 ( .A(n647), .Y(n29) );
  AND2X1 U203 ( .A(n384), .B(n438), .Y(n646) );
  INVX1 U204 ( .A(n646), .Y(n30) );
  AND2X1 U205 ( .A(n383), .B(n438), .Y(n645) );
  INVX1 U206 ( .A(n645), .Y(n31) );
  AND2X1 U207 ( .A(n382), .B(n438), .Y(n644) );
  INVX1 U208 ( .A(n644), .Y(n32) );
  AND2X1 U209 ( .A(n381), .B(n438), .Y(n643) );
  INVX1 U210 ( .A(n643), .Y(n33) );
  AND2X1 U211 ( .A(n380), .B(n439), .Y(n642) );
  INVX1 U212 ( .A(n642), .Y(n34) );
  AND2X1 U213 ( .A(n379), .B(n439), .Y(n641) );
  INVX1 U214 ( .A(n641), .Y(n35) );
  AND2X1 U215 ( .A(n378), .B(n439), .Y(n640) );
  INVX1 U216 ( .A(n640), .Y(n36) );
  AND2X1 U217 ( .A(n377), .B(n439), .Y(n639) );
  INVX1 U218 ( .A(n639), .Y(n37) );
  AND2X1 U219 ( .A(n413), .B(n439), .Y(n638) );
  INVX1 U220 ( .A(n638), .Y(n38) );
  AND2X1 U221 ( .A(n376), .B(n439), .Y(n637) );
  INVX1 U222 ( .A(n637), .Y(n39) );
  AND2X1 U223 ( .A(n375), .B(n439), .Y(n636) );
  INVX1 U224 ( .A(n636), .Y(n40) );
  AND2X1 U225 ( .A(n374), .B(n439), .Y(n635) );
  INVX1 U226 ( .A(n635), .Y(n41) );
  AND2X1 U227 ( .A(n373), .B(n439), .Y(n634) );
  INVX1 U228 ( .A(n634), .Y(n42) );
  AND2X1 U229 ( .A(n372), .B(n439), .Y(n633) );
  INVX1 U230 ( .A(n633), .Y(n43) );
  AND2X1 U231 ( .A(n371), .B(n439), .Y(n632) );
  INVX1 U232 ( .A(n632), .Y(n44) );
  AND2X1 U233 ( .A(n370), .B(n439), .Y(n631) );
  INVX1 U234 ( .A(n631), .Y(n45) );
  AND2X1 U235 ( .A(n369), .B(n439), .Y(n630) );
  INVX1 U236 ( .A(n630), .Y(n46) );
  AND2X1 U237 ( .A(n412), .B(n439), .Y(n627) );
  INVX1 U238 ( .A(n627), .Y(n47) );
  AND2X1 U239 ( .A(n368), .B(n439), .Y(n620) );
  INVX1 U240 ( .A(n620), .Y(n48) );
  AND2X1 U241 ( .A(n367), .B(n439), .Y(n619) );
  INVX1 U242 ( .A(n619), .Y(n49) );
  AND2X1 U243 ( .A(n366), .B(n439), .Y(n618) );
  INVX1 U244 ( .A(n618), .Y(n50) );
  AND2X1 U245 ( .A(n365), .B(n439), .Y(n617) );
  INVX1 U246 ( .A(n617), .Y(n51) );
  AND2X1 U247 ( .A(n411), .B(n436), .Y(n616) );
  INVX1 U248 ( .A(n616), .Y(n52) );
  AND2X1 U249 ( .A(n364), .B(n436), .Y(n615) );
  INVX1 U250 ( .A(n615), .Y(n53) );
  AND2X1 U251 ( .A(n363), .B(n435), .Y(n614) );
  INVX1 U252 ( .A(n614), .Y(n54) );
  AND2X1 U253 ( .A(n362), .B(n434), .Y(n613) );
  INVX1 U254 ( .A(n613), .Y(n55) );
  AND2X1 U255 ( .A(n361), .B(n435), .Y(n612) );
  INVX1 U256 ( .A(n612), .Y(n56) );
  AND2X1 U257 ( .A(n410), .B(n434), .Y(n611) );
  INVX1 U258 ( .A(n611), .Y(n57) );
  AND2X1 U259 ( .A(n409), .B(n433), .Y(n610) );
  INVX1 U260 ( .A(n610), .Y(n58) );
  AND2X1 U261 ( .A(n408), .B(n436), .Y(n609) );
  INVX1 U262 ( .A(n609), .Y(n59) );
  AND2X1 U263 ( .A(n407), .B(n433), .Y(n608) );
  INVX1 U264 ( .A(n608), .Y(n60) );
  AND2X1 U265 ( .A(n424), .B(dataIn[55]), .Y(n587) );
  INVX1 U266 ( .A(n587), .Y(n61) );
  AND2X1 U267 ( .A(n596), .B(dataIn[51]), .Y(n583) );
  INVX1 U268 ( .A(n583), .Y(n62) );
  AND2X1 U269 ( .A(n596), .B(dataIn[49]), .Y(n581) );
  INVX1 U270 ( .A(n581), .Y(n63) );
  AND2X1 U271 ( .A(n596), .B(dataIn[26]), .Y(n558) );
  INVX1 U272 ( .A(n558), .Y(n64) );
  AND2X1 U273 ( .A(n596), .B(dataIn[14]), .Y(n546) );
  INVX1 U274 ( .A(n546), .Y(n65) );
  AND2X1 U275 ( .A(dataIn[63]), .B(n530), .Y(n529) );
  INVX1 U276 ( .A(n529), .Y(n66) );
  AND2X1 U277 ( .A(dataIn[62]), .B(n530), .Y(n528) );
  INVX1 U278 ( .A(n528), .Y(n67) );
  AND2X1 U279 ( .A(dataIn[51]), .B(n530), .Y(n517) );
  INVX1 U280 ( .A(n517), .Y(n68) );
  AND2X1 U283 ( .A(dataIn[50]), .B(n530), .Y(n516) );
  INVX1 U289 ( .A(n516), .Y(n69) );
  AND2X1 U291 ( .A(dataIn[38]), .B(n530), .Y(n504) );
  INVX1 U293 ( .A(n504), .Y(n70) );
  AND2X1 U295 ( .A(dataIn[37]), .B(n425), .Y(n503) );
  INVX1 U297 ( .A(n503), .Y(n71) );
  AND2X1 U299 ( .A(dataIn[36]), .B(n425), .Y(n502) );
  INVX1 U301 ( .A(n502), .Y(n72) );
  AND2X1 U303 ( .A(dataIn[26]), .B(n425), .Y(n492) );
  INVX1 U305 ( .A(n492), .Y(n73) );
  AND2X1 U307 ( .A(dataIn[24]), .B(n425), .Y(n490) );
  INVX1 U309 ( .A(n490), .Y(n74) );
  AND2X1 U311 ( .A(dataIn[14]), .B(n530), .Y(n480) );
  INVX1 U313 ( .A(n480), .Y(n75) );
  AND2X1 U315 ( .A(dataIn[11]), .B(n530), .Y(n477) );
  INVX1 U317 ( .A(n477), .Y(n76) );
  BUFX2 U319 ( .A(n464), .Y(n77) );
  OR2X1 U321 ( .A(outputBufferGrant[0]), .B(outputBufferGrant[1]), .Y(n597) );
  INVX1 U323 ( .A(n597), .Y(n78) );
  INVX1 U325 ( .A(n925), .Y(request[0]) );
  INVX1 U327 ( .A(n924), .Y(request[1]) );
  AND2X1 U329 ( .A(n424), .B(dataIn[54]), .Y(n586) );
  INVX1 U331 ( .A(n586), .Y(n81) );
  AND2X1 U333 ( .A(n596), .B(dataIn[50]), .Y(n582) );
  INVX1 U335 ( .A(n582), .Y(n82) );
  AND2X1 U337 ( .A(dataIn[61]), .B(n530), .Y(n527) );
  INVX1 U339 ( .A(n527), .Y(n83) );
  AND2X1 U341 ( .A(dataIn[47]), .B(n530), .Y(n513) );
  INVX1 U343 ( .A(n513), .Y(n84) );
  AND2X1 U345 ( .A(dataIn[35]), .B(n425), .Y(n501) );
  INVX1 U347 ( .A(n501), .Y(n85) );
  AND2X1 U349 ( .A(dataIn[23]), .B(n530), .Y(n489) );
  INVX1 U351 ( .A(n489), .Y(n86) );
  AND2X1 U353 ( .A(dataIn[10]), .B(n530), .Y(n476) );
  INVX1 U355 ( .A(n476), .Y(n87) );
  AND2X1 U357 ( .A(n596), .B(dataIn[38]), .Y(n570) );
  INVX1 U359 ( .A(n570), .Y(n88) );
  AND2X1 U361 ( .A(n596), .B(dataIn[25]), .Y(n557) );
  INVX1 U363 ( .A(n557), .Y(n89) );
  AND2X1 U365 ( .A(n596), .B(dataIn[12]), .Y(n544) );
  INVX1 U367 ( .A(n544), .Y(n90) );
  AND2X1 U369 ( .A(dataIn[60]), .B(n530), .Y(n526) );
  INVX1 U371 ( .A(n526), .Y(n91) );
  AND2X1 U373 ( .A(dataIn[46]), .B(n530), .Y(n512) );
  INVX1 U375 ( .A(n512), .Y(n92) );
  AND2X1 U377 ( .A(dataIn[34]), .B(n425), .Y(n500) );
  INVX1 U379 ( .A(n500), .Y(n93) );
  AND2X1 U381 ( .A(dataIn[22]), .B(n530), .Y(n488) );
  INVX1 U383 ( .A(n488), .Y(n94) );
  AND2X1 U385 ( .A(dataIn[9]), .B(n530), .Y(n475) );
  INVX1 U387 ( .A(n475), .Y(n95) );
  AND2X1 U389 ( .A(n424), .B(dataIn[52]), .Y(n584) );
  INVX1 U391 ( .A(n584), .Y(n96) );
  AND2X1 U393 ( .A(n596), .B(dataIn[37]), .Y(n569) );
  INVX1 U395 ( .A(n569), .Y(n97) );
  AND2X1 U397 ( .A(n596), .B(dataIn[24]), .Y(n556) );
  INVX1 U399 ( .A(n556), .Y(n98) );
  AND2X1 U401 ( .A(n596), .B(dataIn[11]), .Y(n543) );
  INVX1 U403 ( .A(n543), .Y(n99) );
  AND2X1 U405 ( .A(dataIn[59]), .B(n530), .Y(n525) );
  INVX1 U407 ( .A(n525), .Y(n100) );
  AND2X1 U409 ( .A(dataIn[45]), .B(n530), .Y(n511) );
  INVX1 U411 ( .A(n511), .Y(n101) );
  AND2X1 U413 ( .A(dataIn[33]), .B(n425), .Y(n499) );
  INVX1 U415 ( .A(n499), .Y(n102) );
  AND2X1 U417 ( .A(dataIn[21]), .B(n530), .Y(n487) );
  INVX1 U419 ( .A(n487), .Y(n103) );
  AND2X1 U421 ( .A(dataIn[8]), .B(n530), .Y(n474) );
  INVX1 U423 ( .A(n474), .Y(n104) );
  AND2X1 U425 ( .A(n424), .B(dataIn[63]), .Y(n595) );
  INVX1 U427 ( .A(n595), .Y(n105) );
  AND2X1 U429 ( .A(n596), .B(dataIn[48]), .Y(n580) );
  INVX1 U431 ( .A(n580), .Y(n106) );
  AND2X1 U433 ( .A(n596), .B(dataIn[36]), .Y(n568) );
  INVX1 U435 ( .A(n568), .Y(n107) );
  AND2X1 U437 ( .A(n596), .B(dataIn[23]), .Y(n555) );
  INVX1 U439 ( .A(n555), .Y(n108) );
  AND2X1 U441 ( .A(n596), .B(dataIn[10]), .Y(n542) );
  INVX1 U443 ( .A(n542), .Y(n109) );
  AND2X1 U445 ( .A(dataIn[58]), .B(n530), .Y(n524) );
  INVX1 U447 ( .A(n524), .Y(n110) );
  AND2X1 U449 ( .A(dataIn[44]), .B(n530), .Y(n510) );
  INVX1 U451 ( .A(n510), .Y(n111) );
  AND2X1 U453 ( .A(dataIn[32]), .B(n425), .Y(n498) );
  INVX1 U455 ( .A(n498), .Y(n112) );
  AND2X1 U457 ( .A(dataIn[20]), .B(n530), .Y(n486) );
  INVX1 U459 ( .A(n486), .Y(n113) );
  AND2X1 U461 ( .A(dataIn[7]), .B(n530), .Y(n473) );
  INVX1 U463 ( .A(n473), .Y(n114) );
  AND2X1 U465 ( .A(n424), .B(dataIn[62]), .Y(n594) );
  INVX1 U467 ( .A(n594), .Y(n115) );
  AND2X1 U469 ( .A(n596), .B(dataIn[47]), .Y(n579) );
  INVX1 U471 ( .A(n579), .Y(n116) );
  AND2X1 U473 ( .A(n596), .B(dataIn[35]), .Y(n567) );
  INVX1 U475 ( .A(n567), .Y(n117) );
  AND2X1 U477 ( .A(n596), .B(dataIn[22]), .Y(n554) );
  INVX1 U479 ( .A(n554), .Y(n118) );
  AND2X1 U481 ( .A(n596), .B(dataIn[9]), .Y(n541) );
  INVX1 U483 ( .A(n541), .Y(n119) );
  AND2X1 U485 ( .A(dataIn[57]), .B(n530), .Y(n523) );
  INVX1 U487 ( .A(n523), .Y(n120) );
  AND2X1 U489 ( .A(dataIn[43]), .B(n530), .Y(n509) );
  INVX1 U491 ( .A(n509), .Y(n121) );
  AND2X1 U493 ( .A(dataIn[31]), .B(n425), .Y(n497) );
  INVX1 U495 ( .A(n497), .Y(n122) );
  AND2X1 U497 ( .A(dataIn[19]), .B(n530), .Y(n485) );
  INVX1 U499 ( .A(n485), .Y(n123) );
  AND2X1 U501 ( .A(dataIn[6]), .B(n530), .Y(n472) );
  INVX1 U503 ( .A(n472), .Y(n124) );
  AND2X1 U505 ( .A(n424), .B(dataIn[61]), .Y(n593) );
  INVX1 U507 ( .A(n593), .Y(n125) );
  AND2X1 U509 ( .A(n596), .B(dataIn[46]), .Y(n578) );
  INVX1 U511 ( .A(n578), .Y(n126) );
  AND2X1 U513 ( .A(n596), .B(dataIn[34]), .Y(n566) );
  INVX1 U515 ( .A(n566), .Y(n127) );
  AND2X1 U517 ( .A(n596), .B(dataIn[21]), .Y(n553) );
  INVX1 U519 ( .A(n553), .Y(n128) );
  AND2X1 U521 ( .A(n596), .B(dataIn[8]), .Y(n540) );
  INVX1 U523 ( .A(n540), .Y(n129) );
  AND2X1 U525 ( .A(dataIn[55]), .B(n530), .Y(n521) );
  INVX1 U527 ( .A(n521), .Y(n130) );
  AND2X1 U529 ( .A(dataIn[42]), .B(n530), .Y(n508) );
  INVX1 U531 ( .A(n508), .Y(n131) );
  AND2X1 U533 ( .A(dataIn[30]), .B(n425), .Y(n496) );
  INVX1 U535 ( .A(n496), .Y(n132) );
  AND2X1 U537 ( .A(dataIn[18]), .B(n530), .Y(n484) );
  INVX1 U539 ( .A(n484), .Y(n133) );
  AND2X1 U541 ( .A(dataIn[5]), .B(n530), .Y(n471) );
  INVX1 U543 ( .A(n471), .Y(n134) );
  AND2X1 U545 ( .A(n424), .B(dataIn[60]), .Y(n592) );
  INVX1 U547 ( .A(n592), .Y(n135) );
  AND2X1 U549 ( .A(n596), .B(dataIn[45]), .Y(n577) );
  INVX1 U551 ( .A(n577), .Y(n136) );
  AND2X1 U552 ( .A(n596), .B(dataIn[33]), .Y(n565) );
  INVX1 U554 ( .A(n565), .Y(n137) );
  AND2X1 U556 ( .A(n596), .B(dataIn[20]), .Y(n552) );
  INVX1 U557 ( .A(n552), .Y(n138) );
  AND2X1 U559 ( .A(n596), .B(dataIn[7]), .Y(n539) );
  INVX1 U561 ( .A(n539), .Y(n139) );
  AND2X1 U563 ( .A(dataIn[54]), .B(n530), .Y(n520) );
  INVX1 U565 ( .A(n520), .Y(n148) );
  AND2X1 U567 ( .A(dataIn[41]), .B(n530), .Y(n507) );
  INVX1 U569 ( .A(n507), .Y(n149) );
  AND2X1 U571 ( .A(dataIn[29]), .B(n425), .Y(n495) );
  INVX1 U573 ( .A(n495), .Y(n150) );
  AND2X1 U575 ( .A(dataIn[17]), .B(n530), .Y(n483) );
  INVX1 U577 ( .A(n483), .Y(n151) );
  AND2X1 U579 ( .A(dataIn[4]), .B(n530), .Y(n470) );
  INVX1 U581 ( .A(n470), .Y(n160) );
  AND2X1 U583 ( .A(n424), .B(dataIn[59]), .Y(n591) );
  INVX1 U585 ( .A(n591), .Y(n161) );
  AND2X1 U587 ( .A(n596), .B(dataIn[44]), .Y(n576) );
  INVX1 U595 ( .A(n576), .Y(n162) );
  AND2X1 U599 ( .A(n596), .B(dataIn[32]), .Y(n564) );
  INVX1 U601 ( .A(n564), .Y(n163) );
  AND2X1 U603 ( .A(n596), .B(dataIn[19]), .Y(n551) );
  INVX1 U605 ( .A(n551), .Y(n164) );
  AND2X1 U607 ( .A(n596), .B(dataIn[6]), .Y(n538) );
  INVX1 U609 ( .A(n538), .Y(n165) );
  AND2X1 U611 ( .A(dataIn[56]), .B(n530), .Y(n522) );
  INVX1 U613 ( .A(n522), .Y(n166) );
  AND2X1 U615 ( .A(dataIn[40]), .B(n530), .Y(n506) );
  INVX1 U617 ( .A(n506), .Y(n167) );
  AND2X1 U619 ( .A(dataIn[28]), .B(n425), .Y(n494) );
  INVX1 U621 ( .A(n494), .Y(n168) );
  AND2X1 U623 ( .A(dataIn[16]), .B(n530), .Y(n482) );
  INVX1 U625 ( .A(n482), .Y(n170) );
  AND2X1 U627 ( .A(dataIn[3]), .B(n530), .Y(n469) );
  INVX1 U629 ( .A(n469), .Y(n171) );
  AND2X1 U631 ( .A(n424), .B(dataIn[58]), .Y(n590) );
  INVX1 U633 ( .A(n590), .Y(n172) );
  AND2X1 U635 ( .A(n596), .B(dataIn[43]), .Y(n575) );
  INVX1 U637 ( .A(n575), .Y(n173) );
  AND2X1 U639 ( .A(n596), .B(dataIn[31]), .Y(n563) );
  INVX1 U641 ( .A(n563), .Y(n174) );
  AND2X1 U643 ( .A(n596), .B(dataIn[18]), .Y(n550) );
  INVX1 U645 ( .A(n550), .Y(n175) );
  AND2X1 U647 ( .A(n596), .B(dataIn[5]), .Y(n537) );
  INVX1 U649 ( .A(n537), .Y(n176) );
  AND2X1 U651 ( .A(n808), .B(n807), .Y(n603) );
  INVX1 U653 ( .A(n603), .Y(n178) );
  AND2X1 U655 ( .A(n604), .B(n605), .Y(n169) );
  INVX1 U657 ( .A(n169), .Y(n179) );
  AND2X1 U659 ( .A(n868), .B(n867), .Y(n606) );
  INVX1 U661 ( .A(n606), .Y(n180) );
  AND2X1 U663 ( .A(dataIn[39]), .B(n530), .Y(n505) );
  INVX1 U665 ( .A(n505), .Y(n181) );
  AND2X1 U667 ( .A(dataIn[27]), .B(n425), .Y(n493) );
  INVX1 U669 ( .A(n493), .Y(n182) );
  AND2X1 U671 ( .A(dataIn[15]), .B(n530), .Y(n481) );
  INVX1 U673 ( .A(n481), .Y(n183) );
  AND2X1 U675 ( .A(dataIn[2]), .B(n530), .Y(n468) );
  INVX1 U677 ( .A(n468), .Y(n184) );
  AND2X1 U679 ( .A(n424), .B(dataIn[57]), .Y(n589) );
  INVX1 U681 ( .A(n589), .Y(n314) );
  AND2X1 U682 ( .A(n596), .B(dataIn[42]), .Y(n574) );
  INVX1 U683 ( .A(n574), .Y(n316) );
  AND2X1 U684 ( .A(n596), .B(dataIn[30]), .Y(n562) );
  INVX1 U685 ( .A(n562), .Y(n317) );
  AND2X1 U686 ( .A(n596), .B(dataIn[17]), .Y(n549) );
  INVX1 U687 ( .A(n549), .Y(n318) );
  AND2X1 U688 ( .A(n596), .B(dataIn[3]), .Y(n535) );
  INVX1 U689 ( .A(n535), .Y(n319) );
  AND2X1 U690 ( .A(dataIn[53]), .B(n530), .Y(n519) );
  INVX1 U691 ( .A(n519), .Y(n320) );
  AND2X1 U692 ( .A(n872), .B(n871), .Y(n607) );
  INVX1 U693 ( .A(n607), .Y(n321) );
  AND2X1 U694 ( .A(n600), .B(n601), .Y(n177) );
  INVX1 U695 ( .A(n177), .Y(n322) );
  AND2X1 U696 ( .A(n804), .B(n803), .Y(n602) );
  INVX1 U697 ( .A(n602), .Y(n323) );
  AND2X1 U698 ( .A(dataIn[13]), .B(n530), .Y(n479) );
  INVX1 U699 ( .A(n479), .Y(n324) );
  AND2X1 U700 ( .A(dataIn[1]), .B(n530), .Y(n467) );
  INVX1 U701 ( .A(n467), .Y(n325) );
  AND2X1 U702 ( .A(n424), .B(dataIn[53]), .Y(n585) );
  INVX1 U703 ( .A(n585), .Y(n326) );
  AND2X1 U704 ( .A(n596), .B(dataIn[41]), .Y(n573) );
  INVX1 U705 ( .A(n573), .Y(n327) );
  AND2X1 U706 ( .A(n596), .B(dataIn[29]), .Y(n561) );
  INVX1 U707 ( .A(n561), .Y(n328) );
  AND2X1 U708 ( .A(n596), .B(dataIn[15]), .Y(n547) );
  INVX1 U709 ( .A(n547), .Y(n329) );
  AND2X1 U710 ( .A(n424), .B(dataIn[2]), .Y(n534) );
  INVX1 U711 ( .A(n534), .Y(n330) );
  AND2X1 U712 ( .A(dataIn[52]), .B(n530), .Y(n518) );
  INVX1 U713 ( .A(n518), .Y(n331) );
  AND2X1 U714 ( .A(dataIn[49]), .B(n530), .Y(n515) );
  INVX1 U715 ( .A(n515), .Y(n332) );
  BUFX2 U716 ( .A(oddBuffer[49]), .Y(n333) );
  BUFX2 U717 ( .A(evenBuffer[53]), .Y(n334) );
  AND2X1 U718 ( .A(dataIn[25]), .B(n425), .Y(n491) );
  INVX1 U719 ( .A(n491), .Y(n335) );
  AND2X1 U720 ( .A(dataIn[12]), .B(n530), .Y(n478) );
  INVX1 U721 ( .A(n478), .Y(n336) );
  AND2X1 U722 ( .A(dataIn[0]), .B(n530), .Y(n466) );
  INVX1 U723 ( .A(n466), .Y(n337) );
  AND2X1 U724 ( .A(n424), .B(dataIn[56]), .Y(n588) );
  INVX1 U725 ( .A(n588), .Y(n338) );
  AND2X1 U726 ( .A(n596), .B(dataIn[39]), .Y(n571) );
  INVX1 U727 ( .A(n571), .Y(n339) );
  AND2X1 U728 ( .A(n596), .B(dataIn[27]), .Y(n559) );
  INVX1 U729 ( .A(n559), .Y(n340) );
  AND2X1 U730 ( .A(n596), .B(dataIn[13]), .Y(n545) );
  INVX1 U731 ( .A(n545), .Y(n341) );
  AND2X1 U732 ( .A(n596), .B(dataIn[1]), .Y(n533) );
  INVX1 U733 ( .A(n533), .Y(n342) );
  AND2X1 U734 ( .A(dataIn[48]), .B(n530), .Y(n514) );
  INVX1 U735 ( .A(n514), .Y(n343) );
  BUFX2 U736 ( .A(oddBuffer[53]), .Y(n344) );
  BUFX2 U737 ( .A(evenBuffer[49]), .Y(n345) );
  AND2X1 U738 ( .A(n596), .B(dataIn[40]), .Y(n572) );
  INVX1 U739 ( .A(n572), .Y(n346) );
  AND2X1 U740 ( .A(n596), .B(dataIn[28]), .Y(n560) );
  INVX1 U741 ( .A(n560), .Y(n347) );
  AND2X1 U742 ( .A(n596), .B(dataIn[16]), .Y(n548) );
  INVX1 U743 ( .A(n548), .Y(n348) );
  AND2X1 U744 ( .A(n596), .B(dataIn[4]), .Y(n536) );
  INVX1 U745 ( .A(n536), .Y(n349) );
  AND2X1 U746 ( .A(n596), .B(dataIn[0]), .Y(n532) );
  INVX1 U747 ( .A(n532), .Y(n350) );
  AND2X1 U748 ( .A(n437), .B(n465), .Y(n530) );
  INVX1 U749 ( .A(n530), .Y(n351) );
  BUFX2 U750 ( .A(oddBuffer[55]), .Y(n352) );
  BUFX2 U751 ( .A(oddBufferFull), .Y(n353) );
  BUFX2 U752 ( .A(oddBuffer[54]), .Y(n354) );
  BUFX2 U753 ( .A(oddBuffer[51]), .Y(n355) );
  BUFX2 U754 ( .A(oddBuffer[50]), .Y(n356) );
  BUFX2 U755 ( .A(oddBuffer[48]), .Y(n357) );
  BUFX2 U756 ( .A(evenBuffer[52]), .Y(n358) );
  AND2X1 U757 ( .A(sendIn), .B(n437), .Y(n598) );
  INVX1 U758 ( .A(n598), .Y(n359) );
  AND2X1 U759 ( .A(n531), .B(n442), .Y(n596) );
  INVX1 U760 ( .A(n596), .Y(n360) );
  BUFX2 U761 ( .A(oddBuffer[63]), .Y(n361) );
  BUFX2 U762 ( .A(oddBuffer[62]), .Y(n362) );
  BUFX2 U763 ( .A(oddBuffer[61]), .Y(n363) );
  BUFX2 U764 ( .A(oddBuffer[60]), .Y(n364) );
  BUFX2 U765 ( .A(oddBuffer[59]), .Y(n365) );
  BUFX2 U766 ( .A(oddBuffer[58]), .Y(n366) );
  BUFX2 U767 ( .A(oddBuffer[57]), .Y(n367) );
  BUFX2 U768 ( .A(oddBuffer[56]), .Y(n368) );
  BUFX2 U769 ( .A(oddBuffer[47]), .Y(n369) );
  BUFX2 U770 ( .A(oddBuffer[46]), .Y(n370) );
  BUFX2 U771 ( .A(oddBuffer[45]), .Y(n371) );
  BUFX2 U772 ( .A(oddBuffer[44]), .Y(n372) );
  BUFX2 U773 ( .A(oddBuffer[43]), .Y(n373) );
  BUFX2 U774 ( .A(oddBuffer[42]), .Y(n374) );
  BUFX2 U775 ( .A(oddBuffer[41]), .Y(n375) );
  BUFX2 U776 ( .A(oddBuffer[40]), .Y(n376) );
  BUFX2 U777 ( .A(oddBuffer[39]), .Y(n377) );
  BUFX2 U778 ( .A(oddBuffer[38]), .Y(n378) );
  BUFX2 U779 ( .A(oddBuffer[37]), .Y(n379) );
  BUFX2 U780 ( .A(oddBuffer[36]), .Y(n380) );
  BUFX2 U781 ( .A(oddBuffer[35]), .Y(n381) );
  BUFX2 U782 ( .A(oddBuffer[34]), .Y(n382) );
  BUFX2 U783 ( .A(oddBuffer[33]), .Y(n383) );
  BUFX2 U784 ( .A(oddBuffer[32]), .Y(n384) );
  BUFX2 U785 ( .A(oddBuffer[31]), .Y(n385) );
  BUFX2 U786 ( .A(oddBuffer[30]), .Y(n386) );
  BUFX2 U787 ( .A(oddBuffer[29]), .Y(n387) );
  BUFX2 U788 ( .A(oddBuffer[28]), .Y(n388) );
  BUFX2 U789 ( .A(oddBuffer[27]), .Y(n389) );
  BUFX2 U790 ( .A(oddBuffer[26]), .Y(n390) );
  BUFX2 U791 ( .A(oddBuffer[25]), .Y(n391) );
  BUFX2 U792 ( .A(oddBuffer[24]), .Y(n392) );
  BUFX2 U793 ( .A(oddBuffer[23]), .Y(n393) );
  BUFX2 U794 ( .A(oddBuffer[22]), .Y(n394) );
  BUFX2 U795 ( .A(oddBuffer[21]), .Y(n395) );
  BUFX2 U796 ( .A(oddBuffer[20]), .Y(n396) );
  BUFX2 U797 ( .A(oddBuffer[19]), .Y(n397) );
  BUFX2 U798 ( .A(oddBuffer[18]), .Y(n398) );
  BUFX2 U799 ( .A(oddBuffer[17]), .Y(n399) );
  BUFX2 U800 ( .A(oddBuffer[16]), .Y(n400) );
  BUFX2 U801 ( .A(oddBuffer[15]), .Y(n401) );
  BUFX2 U802 ( .A(oddBuffer[14]), .Y(n402) );
  BUFX2 U803 ( .A(oddBuffer[13]), .Y(n403) );
  BUFX2 U804 ( .A(oddBuffer[12]), .Y(n404) );
  BUFX2 U805 ( .A(oddBuffer[11]), .Y(n405) );
  BUFX2 U806 ( .A(oddBuffer[10]), .Y(n406) );
  BUFX2 U807 ( .A(oddBuffer[9]), .Y(n407) );
  BUFX2 U808 ( .A(oddBuffer[8]), .Y(n408) );
  BUFX2 U809 ( .A(oddBuffer[7]), .Y(n409) );
  BUFX2 U810 ( .A(oddBuffer[6]), .Y(n410) );
  BUFX2 U811 ( .A(oddBuffer[5]), .Y(n411) );
  BUFX2 U812 ( .A(oddBuffer[4]), .Y(n412) );
  BUFX2 U813 ( .A(oddBuffer[3]), .Y(n413) );
  BUFX2 U814 ( .A(oddBuffer[2]), .Y(n414) );
  BUFX2 U815 ( .A(oddBuffer[1]), .Y(n415) );
  BUFX2 U816 ( .A(oddBuffer[0]), .Y(n416) );
  BUFX2 U817 ( .A(evenBuffer[55]), .Y(n417) );
  BUFX2 U818 ( .A(evenBufferFull), .Y(n418) );
  BUFX2 U819 ( .A(evenBuffer[54]), .Y(n419) );
  BUFX2 U820 ( .A(evenBuffer[51]), .Y(n420) );
  BUFX2 U821 ( .A(evenBuffer[50]), .Y(n421) );
  BUFX2 U822 ( .A(oddBuffer[52]), .Y(n422) );
  BUFX2 U823 ( .A(evenBuffer[48]), .Y(n423) );
  INVX1 U824 ( .A(n441), .Y(n432) );
  INVX1 U825 ( .A(n440), .Y(n437) );
  INVX1 U826 ( .A(n442), .Y(n438) );
  INVX1 U827 ( .A(n442), .Y(n439) );
  INVX1 U828 ( .A(n440), .Y(n436) );
  INVX1 U829 ( .A(n440), .Y(n435) );
  INVX1 U830 ( .A(n441), .Y(n434) );
  INVX1 U831 ( .A(n441), .Y(n433) );
  INVX1 U832 ( .A(n351), .Y(n425) );
  INVX1 U833 ( .A(n360), .Y(n424) );
  INVX1 U834 ( .A(n429), .Y(n440) );
  INVX1 U835 ( .A(n429), .Y(n441) );
  INVX1 U836 ( .A(n431), .Y(n429) );
  INVX1 U837 ( .A(n430), .Y(n442) );
  INVX1 U838 ( .A(n431), .Y(n430) );
  INVX1 U839 ( .A(polarity), .Y(n431) );
  INVX1 U840 ( .A(reset), .Y(n428) );
  INVX1 U841 ( .A(reset), .Y(n426) );
  INVX1 U842 ( .A(reset), .Y(n427) );
  INVX1 U843 ( .A(n423), .Y(n874) );
  INVX1 U844 ( .A(n345), .Y(n873) );
  INVX1 U845 ( .A(n358), .Y(n870) );
  INVX1 U846 ( .A(n415), .Y(n857) );
  INVX1 U847 ( .A(n414), .Y(n856) );
  INVX1 U848 ( .A(n413), .Y(n855) );
  INVX1 U849 ( .A(n412), .Y(n854) );
  INVX1 U850 ( .A(n411), .Y(n853) );
  INVX1 U851 ( .A(n410), .Y(n852) );
  INVX1 U852 ( .A(n409), .Y(n851) );
  INVX1 U853 ( .A(n408), .Y(n850) );
  INVX1 U854 ( .A(n407), .Y(n849) );
  INVX1 U855 ( .A(n406), .Y(n848) );
  INVX1 U856 ( .A(n405), .Y(n847) );
  INVX1 U857 ( .A(n404), .Y(n846) );
  INVX1 U858 ( .A(n403), .Y(n845) );
  INVX1 U859 ( .A(n402), .Y(n844) );
  INVX1 U860 ( .A(n401), .Y(n843) );
  INVX1 U861 ( .A(n400), .Y(n842) );
  INVX1 U862 ( .A(n399), .Y(n841) );
  INVX1 U863 ( .A(n398), .Y(n840) );
  INVX1 U864 ( .A(n397), .Y(n839) );
  INVX1 U865 ( .A(n396), .Y(n838) );
  INVX1 U866 ( .A(n395), .Y(n837) );
  INVX1 U867 ( .A(n394), .Y(n836) );
  INVX1 U868 ( .A(n393), .Y(n835) );
  INVX1 U869 ( .A(n392), .Y(n834) );
  INVX1 U870 ( .A(n391), .Y(n833) );
  INVX1 U871 ( .A(n390), .Y(n832) );
  INVX1 U872 ( .A(n389), .Y(n831) );
  INVX1 U873 ( .A(n388), .Y(n830) );
  INVX1 U874 ( .A(n387), .Y(n829) );
  INVX1 U875 ( .A(n386), .Y(n828) );
  INVX1 U876 ( .A(n385), .Y(n827) );
  INVX1 U877 ( .A(n384), .Y(n826) );
  INVX1 U878 ( .A(n383), .Y(n825) );
  INVX1 U879 ( .A(n382), .Y(n824) );
  INVX1 U880 ( .A(n381), .Y(n823) );
  INVX1 U881 ( .A(n380), .Y(n822) );
  INVX1 U882 ( .A(n379), .Y(n821) );
  INVX1 U883 ( .A(n378), .Y(n820) );
  INVX1 U884 ( .A(n377), .Y(n819) );
  INVX1 U885 ( .A(n376), .Y(n818) );
  INVX1 U886 ( .A(n375), .Y(n817) );
  INVX1 U887 ( .A(n374), .Y(n816) );
  INVX1 U888 ( .A(n373), .Y(n815) );
  INVX1 U889 ( .A(n372), .Y(n814) );
  INVX1 U890 ( .A(n371), .Y(n813) );
  INVX1 U891 ( .A(n370), .Y(n812) );
  INVX1 U892 ( .A(n369), .Y(n811) );
  INVX1 U893 ( .A(n357), .Y(n810) );
  INVX1 U894 ( .A(n333), .Y(n809) );
  INVX1 U895 ( .A(n422), .Y(n806) );
  INVX1 U896 ( .A(n334), .Y(n869) );
  INVX1 U897 ( .A(n416), .Y(n858) );
  INVX1 U898 ( .A(n344), .Y(n805) );
  INVX1 U899 ( .A(n368), .Y(n802) );
  INVX1 U900 ( .A(n367), .Y(n459) );
  INVX1 U901 ( .A(n366), .Y(n458) );
  INVX1 U902 ( .A(n365), .Y(n457) );
  INVX1 U903 ( .A(n364), .Y(n456) );
  INVX1 U904 ( .A(n363), .Y(n455) );
  INVX1 U905 ( .A(n362), .Y(n454) );
  INVX1 U906 ( .A(n361), .Y(n453) );
  INVX1 U907 ( .A(n629), .Y(dataOut[48]) );
  INVX1 U908 ( .A(n628), .Y(dataOut[49]) );
  INVX1 U909 ( .A(n626), .Y(dataOut[50]) );
  INVX1 U910 ( .A(n625), .Y(dataOut[51]) );
  INVX1 U911 ( .A(n624), .Y(dataOut[52]) );
  INVX1 U912 ( .A(n623), .Y(dataOut[53]) );
  INVX1 U913 ( .A(n622), .Y(dataOut[54]) );
  INVX1 U914 ( .A(n621), .Y(dataOut[55]) );
  INVX1 U915 ( .A(n356), .Y(n808) );
  INVX1 U916 ( .A(n354), .Y(n804) );
  INVX1 U917 ( .A(n421), .Y(n872) );
  INVX1 U918 ( .A(n419), .Y(n868) );
  INVX1 U919 ( .A(n355), .Y(n807) );
  INVX1 U920 ( .A(n420), .Y(n871) );
  INVX1 U921 ( .A(n418), .Y(n452) );
  INVX1 U922 ( .A(n353), .Y(n451) );
  INVX1 U923 ( .A(n352), .Y(n803) );
  INVX1 U924 ( .A(n417), .Y(n867) );
  INVX1 U925 ( .A(sendIn), .Y(n923) );
  INVX1 U926 ( .A(evenBuffer[0]), .Y(n922) );
  INVX1 U927 ( .A(evenBuffer[1]), .Y(n921) );
  INVX1 U928 ( .A(evenBuffer[2]), .Y(n920) );
  INVX1 U929 ( .A(evenBuffer[3]), .Y(n919) );
  INVX1 U930 ( .A(evenBuffer[4]), .Y(n918) );
  INVX1 U931 ( .A(evenBuffer[5]), .Y(n917) );
  INVX1 U932 ( .A(evenBuffer[6]), .Y(n916) );
  INVX1 U933 ( .A(evenBuffer[7]), .Y(n915) );
  INVX1 U934 ( .A(evenBuffer[8]), .Y(n914) );
  INVX1 U935 ( .A(evenBuffer[9]), .Y(n913) );
  INVX1 U936 ( .A(evenBuffer[10]), .Y(n912) );
  INVX1 U937 ( .A(evenBuffer[11]), .Y(n911) );
  INVX1 U938 ( .A(evenBuffer[12]), .Y(n910) );
  INVX1 U939 ( .A(evenBuffer[13]), .Y(n909) );
  INVX1 U940 ( .A(evenBuffer[14]), .Y(n908) );
  INVX1 U941 ( .A(evenBuffer[15]), .Y(n907) );
  INVX1 U942 ( .A(evenBuffer[16]), .Y(n906) );
  INVX1 U943 ( .A(evenBuffer[17]), .Y(n905) );
  INVX1 U944 ( .A(evenBuffer[18]), .Y(n904) );
  INVX1 U945 ( .A(evenBuffer[19]), .Y(n903) );
  INVX1 U946 ( .A(evenBuffer[20]), .Y(n902) );
  INVX1 U947 ( .A(evenBuffer[21]), .Y(n901) );
  INVX1 U948 ( .A(evenBuffer[22]), .Y(n900) );
  INVX1 U949 ( .A(evenBuffer[23]), .Y(n899) );
  INVX1 U950 ( .A(evenBuffer[24]), .Y(n898) );
  INVX1 U951 ( .A(evenBuffer[25]), .Y(n897) );
  INVX1 U952 ( .A(evenBuffer[26]), .Y(n896) );
  INVX1 U953 ( .A(evenBuffer[27]), .Y(n895) );
  INVX1 U954 ( .A(evenBuffer[28]), .Y(n894) );
  INVX1 U955 ( .A(evenBuffer[29]), .Y(n893) );
  INVX1 U956 ( .A(evenBuffer[30]), .Y(n892) );
  INVX1 U957 ( .A(evenBuffer[31]), .Y(n891) );
  INVX1 U958 ( .A(evenBuffer[32]), .Y(n890) );
  INVX1 U959 ( .A(evenBuffer[33]), .Y(n889) );
  INVX1 U960 ( .A(evenBuffer[34]), .Y(n888) );
  INVX1 U961 ( .A(evenBuffer[35]), .Y(n887) );
  INVX1 U962 ( .A(evenBuffer[36]), .Y(n886) );
  INVX1 U963 ( .A(evenBuffer[37]), .Y(n885) );
  INVX1 U964 ( .A(evenBuffer[38]), .Y(n884) );
  INVX1 U965 ( .A(evenBuffer[39]), .Y(n883) );
  INVX1 U966 ( .A(evenBuffer[40]), .Y(n882) );
  INVX1 U967 ( .A(evenBuffer[41]), .Y(n881) );
  INVX1 U968 ( .A(evenBuffer[42]), .Y(n880) );
  INVX1 U969 ( .A(evenBuffer[43]), .Y(n879) );
  INVX1 U970 ( .A(evenBuffer[44]), .Y(n878) );
  INVX1 U971 ( .A(evenBuffer[45]), .Y(n877) );
  INVX1 U972 ( .A(evenBuffer[46]), .Y(n876) );
  INVX1 U973 ( .A(evenBuffer[47]), .Y(n875) );
  INVX1 U974 ( .A(evenBuffer[56]), .Y(n866) );
  INVX1 U975 ( .A(evenBuffer[57]), .Y(n865) );
  INVX1 U976 ( .A(evenBuffer[58]), .Y(n864) );
  INVX1 U977 ( .A(evenBuffer[59]), .Y(n863) );
  INVX1 U978 ( .A(evenBuffer[60]), .Y(n862) );
  INVX1 U979 ( .A(evenBuffer[61]), .Y(n861) );
  INVX1 U980 ( .A(evenBuffer[62]), .Y(n860) );
  INVX1 U981 ( .A(evenBuffer[63]), .Y(n859) );
  XNOR2X1 U982 ( .A(n352), .B(sub_131_aco_carry[7]), .Y(n159) );
  XNOR2X1 U983 ( .A(n354), .B(sub_131_aco_carry[6]), .Y(n158) );
  XNOR2X1 U984 ( .A(n344), .B(sub_131_aco_carry[5]), .Y(n157) );
  XNOR2X1 U985 ( .A(n422), .B(sub_131_aco_carry[4]), .Y(n156) );
  XNOR2X1 U986 ( .A(n355), .B(sub_131_aco_carry[3]), .Y(n155) );
  XNOR2X1 U987 ( .A(n356), .B(sub_131_aco_carry[2]), .Y(n154) );
  XNOR2X1 U988 ( .A(n333), .B(sub_131_aco_carry[1]), .Y(n153) );
  XNOR2X1 U989 ( .A(n357), .B(n177), .Y(n152) );
  XNOR2X1 U990 ( .A(n417), .B(sub_111_aco_carry[7]), .Y(n147) );
  XNOR2X1 U991 ( .A(n419), .B(sub_111_aco_carry[6]), .Y(n146) );
  XNOR2X1 U992 ( .A(n334), .B(sub_111_aco_carry[5]), .Y(n145) );
  XNOR2X1 U993 ( .A(n358), .B(sub_111_aco_carry[4]), .Y(n144) );
  XNOR2X1 U994 ( .A(n420), .B(sub_111_aco_carry[3]), .Y(n143) );
  XNOR2X1 U995 ( .A(n421), .B(sub_111_aco_carry[2]), .Y(n142) );
  XNOR2X1 U996 ( .A(n345), .B(sub_111_aco_carry[1]), .Y(n141) );
  XNOR2X1 U997 ( .A(n423), .B(n169), .Y(n140) );
endmodule


module inputBuffer_0 ( clk, reset, polarity, sendIn, readyIn, dataIn, dataOut, 
        request, outputBufferGrant );
  input [63:0] dataIn;
  output [63:0] dataOut;
  output [1:0] request;
  input [1:0] outputBufferGrant;
  input clk, reset, polarity, sendIn;
  output readyIn;
  wire   n1264, n1265, evenBufferFull, oddBufferFull, n140, n141, n142, n143,
         n144, n145, n146, n147, n152, n153, n154, n155, n156, n157, n158,
         n159, n169, n177, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263;
  wire   [63:0] evenBuffer;
  wire   [63:0] oddBuffer;
  wire   [7:1] sub_131_aco_carry;
  wire   [7:1] sub_111_aco_carry;

  NAND3X1 U281 ( .A(n169), .B(n437), .C(n418), .Y(n1262) );
  NAND3X1 U282 ( .A(n353), .B(n177), .C(n429), .Y(n1263) );
  NAND3X1 U284 ( .A(n309), .B(n438), .C(n418), .Y(n1260) );
  NAND3X1 U285 ( .A(n353), .B(n322), .C(n429), .Y(n1261) );
  NOR2X1 U286 ( .A(reset), .B(n77), .Y(readyIn) );
  AOI22X1 U287 ( .A(n429), .B(n449), .C(n448), .D(n439), .Y(n1259) );
  OAI21X1 U288 ( .A(n1258), .B(n919), .C(n337), .Y(n1051) );
  OAI21X1 U290 ( .A(n1258), .B(n918), .C(n325), .Y(n1050) );
  OAI21X1 U292 ( .A(n1258), .B(n917), .C(n314), .Y(n1049) );
  OAI21X1 U294 ( .A(n1258), .B(n916), .C(n302), .Y(n1048) );
  OAI21X1 U296 ( .A(n1258), .B(n915), .C(n292), .Y(n1047) );
  OAI21X1 U298 ( .A(n1258), .B(n914), .C(n282), .Y(n1046) );
  OAI21X1 U300 ( .A(n1258), .B(n913), .C(n272), .Y(n1045) );
  OAI21X1 U302 ( .A(n1258), .B(n912), .C(n262), .Y(n1044) );
  OAI21X1 U304 ( .A(n1258), .B(n911), .C(n252), .Y(n1043) );
  OAI21X1 U306 ( .A(n1258), .B(n910), .C(n243), .Y(n1042) );
  OAI21X1 U308 ( .A(n1258), .B(n909), .C(n235), .Y(n1041) );
  OAI21X1 U310 ( .A(n1258), .B(n908), .C(n76), .Y(n1040) );
  OAI21X1 U312 ( .A(n1258), .B(n907), .C(n336), .Y(n1039) );
  OAI21X1 U314 ( .A(n1258), .B(n906), .C(n324), .Y(n1038) );
  OAI21X1 U316 ( .A(n1258), .B(n905), .C(n75), .Y(n1037) );
  OAI21X1 U318 ( .A(n1258), .B(n904), .C(n313), .Y(n1036) );
  OAI21X1 U320 ( .A(n1258), .B(n903), .C(n301), .Y(n1035) );
  OAI21X1 U322 ( .A(n1258), .B(n902), .C(n291), .Y(n1034) );
  OAI21X1 U324 ( .A(n1258), .B(n901), .C(n281), .Y(n1033) );
  OAI21X1 U326 ( .A(n1258), .B(n900), .C(n271), .Y(n1032) );
  OAI21X1 U328 ( .A(n1258), .B(n899), .C(n261), .Y(n1031) );
  OAI21X1 U330 ( .A(n1258), .B(n898), .C(n251), .Y(n1030) );
  OAI21X1 U332 ( .A(n1258), .B(n897), .C(n242), .Y(n1029) );
  OAI21X1 U334 ( .A(n1258), .B(n896), .C(n234), .Y(n1028) );
  OAI21X1 U336 ( .A(n1258), .B(n895), .C(n74), .Y(n1027) );
  OAI21X1 U338 ( .A(n1258), .B(n894), .C(n335), .Y(n1026) );
  OAI21X1 U340 ( .A(n1258), .B(n893), .C(n73), .Y(n1025) );
  OAI21X1 U342 ( .A(n1258), .B(n892), .C(n312), .Y(n1024) );
  OAI21X1 U344 ( .A(n1258), .B(n891), .C(n300), .Y(n1023) );
  OAI21X1 U346 ( .A(n1258), .B(n890), .C(n290), .Y(n1022) );
  OAI21X1 U348 ( .A(n1258), .B(n889), .C(n280), .Y(n1021) );
  OAI21X1 U350 ( .A(n1258), .B(n888), .C(n270), .Y(n1020) );
  OAI21X1 U352 ( .A(n1258), .B(n887), .C(n260), .Y(n1019) );
  OAI21X1 U354 ( .A(n1258), .B(n886), .C(n250), .Y(n1018) );
  OAI21X1 U356 ( .A(n1258), .B(n885), .C(n241), .Y(n1017) );
  OAI21X1 U358 ( .A(n1258), .B(n884), .C(n233), .Y(n1016) );
  OAI21X1 U360 ( .A(n1258), .B(n883), .C(n72), .Y(n1015) );
  OAI21X1 U362 ( .A(n1258), .B(n882), .C(n71), .Y(n1014) );
  OAI21X1 U364 ( .A(n1258), .B(n881), .C(n70), .Y(n1013) );
  OAI21X1 U366 ( .A(n1258), .B(n880), .C(n311), .Y(n1012) );
  OAI21X1 U368 ( .A(n1258), .B(n879), .C(n299), .Y(n1011) );
  OAI21X1 U370 ( .A(n1258), .B(n878), .C(n289), .Y(n1010) );
  OAI21X1 U372 ( .A(n1258), .B(n877), .C(n279), .Y(n1009) );
  OAI21X1 U374 ( .A(n1258), .B(n876), .C(n269), .Y(n1008) );
  OAI21X1 U376 ( .A(n1258), .B(n875), .C(n259), .Y(n1007) );
  OAI21X1 U378 ( .A(n1258), .B(n874), .C(n249), .Y(n1006) );
  OAI21X1 U380 ( .A(n1258), .B(n873), .C(n240), .Y(n1005) );
  OAI21X1 U382 ( .A(n1258), .B(n872), .C(n232), .Y(n1004) );
  OAI21X1 U384 ( .A(n1258), .B(n871), .C(n343), .Y(n1003) );
  OAI21X1 U386 ( .A(n1258), .B(n870), .C(n332), .Y(n1002) );
  OAI21X1 U388 ( .A(n1258), .B(n869), .C(n69), .Y(n1001) );
  OAI21X1 U390 ( .A(n1258), .B(n868), .C(n68), .Y(n1000) );
  OAI21X1 U392 ( .A(n1258), .B(n867), .C(n331), .Y(n999) );
  OAI21X1 U394 ( .A(n1258), .B(n866), .C(n320), .Y(n998) );
  OAI21X1 U396 ( .A(n1258), .B(n865), .C(n288), .Y(n997) );
  OAI21X1 U398 ( .A(n1258), .B(n864), .C(n278), .Y(n996) );
  OAI21X1 U400 ( .A(n1258), .B(n863), .C(n298), .Y(n995) );
  OAI21X1 U402 ( .A(n1258), .B(n862), .C(n268), .Y(n994) );
  OAI21X1 U404 ( .A(n1258), .B(n861), .C(n258), .Y(n993) );
  OAI21X1 U406 ( .A(n1258), .B(n860), .C(n248), .Y(n992) );
  OAI21X1 U408 ( .A(n1258), .B(n859), .C(n239), .Y(n991) );
  OAI21X1 U410 ( .A(n1258), .B(n858), .C(n231), .Y(n990) );
  OAI21X1 U412 ( .A(n1258), .B(n857), .C(n67), .Y(n989) );
  OAI21X1 U414 ( .A(n1258), .B(n856), .C(n66), .Y(n988) );
  OAI21X1 U416 ( .A(n1192), .B(n855), .C(n350), .Y(n987) );
  OAI21X1 U418 ( .A(n1192), .B(n854), .C(n342), .Y(n986) );
  OAI21X1 U420 ( .A(n1192), .B(n853), .C(n330), .Y(n985) );
  OAI21X1 U422 ( .A(n1192), .B(n852), .C(n319), .Y(n984) );
  OAI21X1 U424 ( .A(n1192), .B(n851), .C(n349), .Y(n983) );
  OAI21X1 U426 ( .A(n1192), .B(n850), .C(n307), .Y(n982) );
  OAI21X1 U428 ( .A(n1192), .B(n849), .C(n297), .Y(n981) );
  OAI21X1 U430 ( .A(n1192), .B(n848), .C(n287), .Y(n980) );
  OAI21X1 U432 ( .A(n1192), .B(n847), .C(n277), .Y(n979) );
  OAI21X1 U434 ( .A(n1192), .B(n846), .C(n267), .Y(n978) );
  OAI21X1 U436 ( .A(n1192), .B(n845), .C(n257), .Y(n977) );
  OAI21X1 U438 ( .A(n1192), .B(n844), .C(n247), .Y(n976) );
  OAI21X1 U440 ( .A(n1192), .B(n843), .C(n238), .Y(n975) );
  OAI21X1 U442 ( .A(n1192), .B(n842), .C(n341), .Y(n974) );
  OAI21X1 U444 ( .A(n1192), .B(n841), .C(n65), .Y(n973) );
  OAI21X1 U446 ( .A(n1192), .B(n840), .C(n329), .Y(n972) );
  OAI21X1 U448 ( .A(n1192), .B(n839), .C(n348), .Y(n971) );
  OAI21X1 U450 ( .A(n1192), .B(n838), .C(n318), .Y(n970) );
  OAI21X1 U452 ( .A(n1192), .B(n837), .C(n306), .Y(n969) );
  OAI21X1 U454 ( .A(n1192), .B(n836), .C(n296), .Y(n968) );
  OAI21X1 U456 ( .A(n1192), .B(n835), .C(n286), .Y(n967) );
  OAI21X1 U458 ( .A(n1192), .B(n834), .C(n276), .Y(n966) );
  OAI21X1 U460 ( .A(n1192), .B(n833), .C(n266), .Y(n965) );
  OAI21X1 U462 ( .A(n1192), .B(n832), .C(n256), .Y(n964) );
  OAI21X1 U464 ( .A(n1192), .B(n831), .C(n246), .Y(n963) );
  OAI21X1 U466 ( .A(n1192), .B(n830), .C(n237), .Y(n962) );
  OAI21X1 U468 ( .A(n1192), .B(n829), .C(n64), .Y(n961) );
  OAI21X1 U470 ( .A(n1192), .B(n828), .C(n340), .Y(n960) );
  OAI21X1 U472 ( .A(n1192), .B(n827), .C(n347), .Y(n959) );
  OAI21X1 U474 ( .A(n1192), .B(n826), .C(n328), .Y(n958) );
  OAI21X1 U476 ( .A(n1192), .B(n825), .C(n317), .Y(n957) );
  OAI21X1 U478 ( .A(n1192), .B(n824), .C(n305), .Y(n956) );
  OAI21X1 U480 ( .A(n1192), .B(n823), .C(n295), .Y(n955) );
  OAI21X1 U482 ( .A(n1192), .B(n822), .C(n285), .Y(n954) );
  OAI21X1 U484 ( .A(n1192), .B(n821), .C(n275), .Y(n953) );
  OAI21X1 U486 ( .A(n1192), .B(n820), .C(n265), .Y(n952) );
  OAI21X1 U488 ( .A(n1192), .B(n819), .C(n255), .Y(n951) );
  OAI21X1 U490 ( .A(n1192), .B(n818), .C(n245), .Y(n950) );
  OAI21X1 U492 ( .A(n1192), .B(n817), .C(n236), .Y(n949) );
  OAI21X1 U494 ( .A(n1192), .B(n816), .C(n339), .Y(n948) );
  OAI21X1 U496 ( .A(n1192), .B(n815), .C(n346), .Y(n947) );
  OAI21X1 U498 ( .A(n1192), .B(n814), .C(n327), .Y(n946) );
  OAI21X1 U500 ( .A(n1192), .B(n813), .C(n316), .Y(n945) );
  OAI21X1 U502 ( .A(n1192), .B(n812), .C(n304), .Y(n944) );
  OAI21X1 U504 ( .A(n1192), .B(n811), .C(n294), .Y(n943) );
  OAI21X1 U506 ( .A(n1192), .B(n810), .C(n284), .Y(n942) );
  OAI21X1 U508 ( .A(n1192), .B(n809), .C(n274), .Y(n941) );
  OAI21X1 U510 ( .A(n1192), .B(n808), .C(n264), .Y(n940) );
  OAI21X1 U512 ( .A(n1192), .B(n807), .C(n254), .Y(n939) );
  OAI21X1 U514 ( .A(n1192), .B(n806), .C(n63), .Y(n938) );
  OAI21X1 U516 ( .A(n1192), .B(n805), .C(n230), .Y(n937) );
  OAI21X1 U518 ( .A(n1192), .B(n804), .C(n62), .Y(n936) );
  OAI21X1 U520 ( .A(n1192), .B(n803), .C(n244), .Y(n935) );
  OAI21X1 U522 ( .A(n1192), .B(n802), .C(n326), .Y(n934) );
  OAI21X1 U524 ( .A(n1192), .B(n459), .C(n229), .Y(n933) );
  OAI21X1 U526 ( .A(n1192), .B(n458), .C(n61), .Y(n932) );
  OAI21X1 U528 ( .A(n1192), .B(n457), .C(n338), .Y(n931) );
  OAI21X1 U530 ( .A(n1192), .B(n456), .C(n315), .Y(n930) );
  OAI21X1 U532 ( .A(n1192), .B(n455), .C(n303), .Y(n929) );
  OAI21X1 U534 ( .A(n1192), .B(n454), .C(n293), .Y(n928) );
  OAI21X1 U536 ( .A(n1192), .B(n453), .C(n283), .Y(n927) );
  OAI21X1 U538 ( .A(n1192), .B(n452), .C(n273), .Y(n926) );
  OAI21X1 U540 ( .A(n1192), .B(n451), .C(n263), .Y(n925) );
  OAI21X1 U542 ( .A(n1192), .B(n450), .C(n253), .Y(n924) );
  OAI21X1 U544 ( .A(n449), .B(n1258), .C(n351), .Y(n923) );
  OAI21X1 U546 ( .A(n429), .B(n78), .C(n359), .Y(n1258) );
  OAI21X1 U548 ( .A(n448), .B(n1192), .C(n360), .Y(n922) );
  OAI21X1 U550 ( .A(n429), .B(n921), .C(n1124), .Y(n1192) );
  NOR3X1 U553 ( .A(n323), .B(n344), .C(n422), .Y(n1122) );
  NOR3X1 U555 ( .A(n308), .B(n333), .C(n357), .Y(n1123) );
  NOR3X1 U558 ( .A(n310), .B(n334), .C(n358), .Y(n1118) );
  NOR3X1 U560 ( .A(n321), .B(n345), .C(n423), .Y(n1119) );
  OAI21X1 U562 ( .A(n430), .B(n910), .C(n60), .Y(dataOut[9]) );
  OAI21X1 U564 ( .A(n430), .B(n911), .C(n59), .Y(dataOut[8]) );
  OAI21X1 U566 ( .A(n430), .B(n912), .C(n58), .Y(dataOut[7]) );
  OAI21X1 U568 ( .A(n430), .B(n913), .C(n57), .Y(dataOut[6]) );
  OAI21X1 U570 ( .A(n430), .B(n856), .C(n56), .Y(dataOut[63]) );
  OAI21X1 U572 ( .A(n430), .B(n857), .C(n55), .Y(dataOut[62]) );
  OAI21X1 U574 ( .A(n430), .B(n858), .C(n54), .Y(dataOut[61]) );
  OAI21X1 U576 ( .A(n430), .B(n859), .C(n53), .Y(dataOut[60]) );
  OAI21X1 U578 ( .A(n430), .B(n914), .C(n52), .Y(dataOut[5]) );
  OAI21X1 U580 ( .A(n430), .B(n860), .C(n51), .Y(dataOut[59]) );
  OAI21X1 U582 ( .A(n431), .B(n861), .C(n50), .Y(dataOut[58]) );
  OAI21X1 U584 ( .A(n431), .B(n862), .C(n49), .Y(dataOut[57]) );
  OAI21X1 U586 ( .A(n431), .B(n863), .C(n48), .Y(dataOut[56]) );
  AOI22X1 U588 ( .A(n147), .B(n439), .C(n159), .D(n429), .Y(n1102) );
  AOI22X1 U589 ( .A(n146), .B(n439), .C(n158), .D(n429), .Y(n1101) );
  AOI22X1 U590 ( .A(n145), .B(n439), .C(n157), .D(n429), .Y(n1100) );
  AOI22X1 U591 ( .A(n144), .B(n439), .C(n156), .D(n429), .Y(n1099) );
  AOI22X1 U592 ( .A(n143), .B(n439), .C(n155), .D(n429), .Y(n1098) );
  AOI22X1 U593 ( .A(n142), .B(n439), .C(n154), .D(n429), .Y(n1097) );
  OAI21X1 U594 ( .A(n431), .B(n915), .C(n47), .Y(dataOut[4]) );
  AOI22X1 U596 ( .A(n141), .B(n439), .C(n153), .D(n429), .Y(n1095) );
  AOI22X1 U597 ( .A(n140), .B(n439), .C(n152), .D(n429), .Y(n1094) );
  OAI21X1 U598 ( .A(n431), .B(n872), .C(n46), .Y(dataOut[47]) );
  OAI21X1 U600 ( .A(n432), .B(n873), .C(n45), .Y(dataOut[46]) );
  OAI21X1 U602 ( .A(n432), .B(n874), .C(n44), .Y(dataOut[45]) );
  OAI21X1 U604 ( .A(n431), .B(n875), .C(n43), .Y(dataOut[44]) );
  OAI21X1 U606 ( .A(n432), .B(n876), .C(n42), .Y(dataOut[43]) );
  OAI21X1 U608 ( .A(n432), .B(n877), .C(n41), .Y(dataOut[42]) );
  OAI21X1 U610 ( .A(n432), .B(n878), .C(n40), .Y(dataOut[41]) );
  OAI21X1 U612 ( .A(n432), .B(n879), .C(n39), .Y(dataOut[40]) );
  OAI21X1 U614 ( .A(n432), .B(n916), .C(n38), .Y(dataOut[3]) );
  OAI21X1 U616 ( .A(n432), .B(n880), .C(n37), .Y(dataOut[39]) );
  OAI21X1 U618 ( .A(n433), .B(n881), .C(n36), .Y(dataOut[38]) );
  OAI21X1 U620 ( .A(n433), .B(n882), .C(n35), .Y(dataOut[37]) );
  OAI21X1 U622 ( .A(n432), .B(n883), .C(n34), .Y(dataOut[36]) );
  OAI21X1 U624 ( .A(n433), .B(n884), .C(n33), .Y(dataOut[35]) );
  OAI21X1 U626 ( .A(n433), .B(n885), .C(n32), .Y(dataOut[34]) );
  OAI21X1 U628 ( .A(n433), .B(n886), .C(n31), .Y(dataOut[33]) );
  OAI21X1 U630 ( .A(n433), .B(n887), .C(n30), .Y(dataOut[32]) );
  OAI21X1 U632 ( .A(n433), .B(n888), .C(n29), .Y(dataOut[31]) );
  OAI21X1 U634 ( .A(n433), .B(n889), .C(n28), .Y(dataOut[30]) );
  OAI21X1 U636 ( .A(n434), .B(n917), .C(n27), .Y(dataOut[2]) );
  OAI21X1 U638 ( .A(n434), .B(n890), .C(n26), .Y(dataOut[29]) );
  OAI21X1 U640 ( .A(n433), .B(n891), .C(n25), .Y(dataOut[28]) );
  OAI21X1 U642 ( .A(n434), .B(n892), .C(n24), .Y(dataOut[27]) );
  OAI21X1 U644 ( .A(n432), .B(n893), .C(n23), .Y(dataOut[26]) );
  OAI21X1 U646 ( .A(n434), .B(n894), .C(n22), .Y(dataOut[25]) );
  OAI21X1 U648 ( .A(n433), .B(n895), .C(n21), .Y(dataOut[24]) );
  OAI21X1 U650 ( .A(n433), .B(n896), .C(n20), .Y(dataOut[23]) );
  OAI21X1 U652 ( .A(n432), .B(n897), .C(n19), .Y(dataOut[22]) );
  OAI21X1 U654 ( .A(n433), .B(n898), .C(n18), .Y(dataOut[21]) );
  OAI21X1 U656 ( .A(n432), .B(n899), .C(n17), .Y(dataOut[20]) );
  OAI21X1 U658 ( .A(n433), .B(n918), .C(n16), .Y(dataOut[1]) );
  OAI21X1 U660 ( .A(n432), .B(n900), .C(n15), .Y(dataOut[19]) );
  OAI21X1 U662 ( .A(n431), .B(n901), .C(n14), .Y(dataOut[18]) );
  OAI21X1 U664 ( .A(n431), .B(n902), .C(n13), .Y(dataOut[17]) );
  OAI21X1 U666 ( .A(n431), .B(n903), .C(n12), .Y(dataOut[16]) );
  OAI21X1 U668 ( .A(n431), .B(n904), .C(n11), .Y(dataOut[15]) );
  OAI21X1 U670 ( .A(n431), .B(n905), .C(n10), .Y(dataOut[14]) );
  OAI21X1 U672 ( .A(n431), .B(n906), .C(n9), .Y(dataOut[13]) );
  OAI21X1 U674 ( .A(n430), .B(n907), .C(n8), .Y(dataOut[12]) );
  OAI21X1 U676 ( .A(n431), .B(n908), .C(n7), .Y(dataOut[11]) );
  OAI21X1 U678 ( .A(n430), .B(n909), .C(n6), .Y(dataOut[10]) );
  OAI21X1 U680 ( .A(n430), .B(n919), .C(n5), .Y(dataOut[0]) );
  DFFSR evenBufferFull_reg ( .D(n923), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBufferFull) );
  DFFSR oddBuffer_reg_3_ ( .D(n984), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[3]) );
  DFFSR oddBuffer_reg_2_ ( .D(n985), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[2]) );
  DFFSR oddBuffer_reg_1_ ( .D(n986), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[1]) );
  DFFSR oddBuffer_reg_0_ ( .D(n987), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[0]) );
  DFFSR oddBufferFull_reg ( .D(n922), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBufferFull) );
  DFFSR evenBuffer_reg_11_ ( .D(n1040), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[11]) );
  DFFSR evenBuffer_reg_63_ ( .D(n988), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[63]) );
  DFFSR evenBuffer_reg_62_ ( .D(n989), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[62]) );
  DFFSR evenBuffer_reg_51_ ( .D(n1000), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[51]) );
  DFFSR evenBuffer_reg_50_ ( .D(n1001), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[50]) );
  DFFSR evenBuffer_reg_38_ ( .D(n1013), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[38]) );
  DFFSR evenBuffer_reg_37_ ( .D(n1014), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[37]) );
  DFFSR evenBuffer_reg_36_ ( .D(n1015), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[36]) );
  DFFSR evenBuffer_reg_26_ ( .D(n1025), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[26]) );
  DFFSR evenBuffer_reg_24_ ( .D(n1027), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[24]) );
  DFFSR evenBuffer_reg_14_ ( .D(n1037), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[14]) );
  DFFSR oddBuffer_reg_51_ ( .D(n936), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[51]) );
  DFFSR oddBuffer_reg_49_ ( .D(n938), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[49]) );
  DFFSR oddBuffer_reg_55_ ( .D(n932), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[55]) );
  DFFSR oddBuffer_reg_26_ ( .D(n961), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[26]) );
  DFFSR oddBuffer_reg_14_ ( .D(n973), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[14]) );
  DFFSR evenBuffer_reg_61_ ( .D(n990), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[61]) );
  DFFSR evenBuffer_reg_60_ ( .D(n991), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[60]) );
  DFFSR evenBuffer_reg_59_ ( .D(n992), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[59]) );
  DFFSR evenBuffer_reg_58_ ( .D(n993), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[58]) );
  DFFSR evenBuffer_reg_57_ ( .D(n994), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[57]) );
  DFFSR evenBuffer_reg_56_ ( .D(n995), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[56]) );
  DFFSR evenBuffer_reg_55_ ( .D(n996), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[55]) );
  DFFSR evenBuffer_reg_54_ ( .D(n997), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[54]) );
  DFFSR evenBuffer_reg_53_ ( .D(n998), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[53]) );
  DFFSR evenBuffer_reg_52_ ( .D(n999), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[52]) );
  DFFSR evenBuffer_reg_0_ ( .D(n1051), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[0]) );
  DFFSR evenBuffer_reg_10_ ( .D(n1041), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[10]) );
  DFFSR evenBuffer_reg_9_ ( .D(n1042), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[9]) );
  DFFSR evenBuffer_reg_8_ ( .D(n1043), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[8]) );
  DFFSR evenBuffer_reg_7_ ( .D(n1044), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[7]) );
  DFFSR evenBuffer_reg_6_ ( .D(n1045), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[6]) );
  DFFSR evenBuffer_reg_5_ ( .D(n1046), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[5]) );
  DFFSR evenBuffer_reg_4_ ( .D(n1047), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[4]) );
  DFFSR evenBuffer_reg_3_ ( .D(n1048), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[3]) );
  DFFSR evenBuffer_reg_2_ ( .D(n1049), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[2]) );
  DFFSR evenBuffer_reg_1_ ( .D(n1050), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[1]) );
  DFFSR evenBuffer_reg_49_ ( .D(n1002), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[49]) );
  DFFSR evenBuffer_reg_48_ ( .D(n1003), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[48]) );
  DFFSR evenBuffer_reg_47_ ( .D(n1004), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[47]) );
  DFFSR evenBuffer_reg_46_ ( .D(n1005), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[46]) );
  DFFSR evenBuffer_reg_45_ ( .D(n1006), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[45]) );
  DFFSR evenBuffer_reg_44_ ( .D(n1007), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[44]) );
  DFFSR evenBuffer_reg_43_ ( .D(n1008), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[43]) );
  DFFSR evenBuffer_reg_42_ ( .D(n1009), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[42]) );
  DFFSR evenBuffer_reg_41_ ( .D(n1010), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[41]) );
  DFFSR evenBuffer_reg_40_ ( .D(n1011), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[40]) );
  DFFSR evenBuffer_reg_39_ ( .D(n1012), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[39]) );
  DFFSR evenBuffer_reg_35_ ( .D(n1016), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[35]) );
  DFFSR evenBuffer_reg_34_ ( .D(n1017), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[34]) );
  DFFSR evenBuffer_reg_33_ ( .D(n1018), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[33]) );
  DFFSR evenBuffer_reg_32_ ( .D(n1019), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[32]) );
  DFFSR evenBuffer_reg_31_ ( .D(n1020), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[31]) );
  DFFSR evenBuffer_reg_30_ ( .D(n1021), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[30]) );
  DFFSR evenBuffer_reg_29_ ( .D(n1022), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[29]) );
  DFFSR evenBuffer_reg_28_ ( .D(n1023), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[28]) );
  DFFSR evenBuffer_reg_27_ ( .D(n1024), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[27]) );
  DFFSR evenBuffer_reg_25_ ( .D(n1026), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[25]) );
  DFFSR evenBuffer_reg_23_ ( .D(n1028), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[23]) );
  DFFSR evenBuffer_reg_22_ ( .D(n1029), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[22]) );
  DFFSR evenBuffer_reg_21_ ( .D(n1030), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[21]) );
  DFFSR evenBuffer_reg_20_ ( .D(n1031), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[20]) );
  DFFSR evenBuffer_reg_19_ ( .D(n1032), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[19]) );
  DFFSR evenBuffer_reg_18_ ( .D(n1033), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[18]) );
  DFFSR evenBuffer_reg_17_ ( .D(n1034), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[17]) );
  DFFSR evenBuffer_reg_16_ ( .D(n1035), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[16]) );
  DFFSR evenBuffer_reg_15_ ( .D(n1036), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[15]) );
  DFFSR evenBuffer_reg_13_ ( .D(n1038), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[13]) );
  DFFSR evenBuffer_reg_12_ ( .D(n1039), .CLK(clk), .R(n920), .S(1'b1), .Q(
        evenBuffer[12]) );
  DFFSR oddBuffer_reg_50_ ( .D(n937), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[50]) );
  DFFSR oddBuffer_reg_48_ ( .D(n939), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[48]) );
  DFFSR oddBuffer_reg_47_ ( .D(n940), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[47]) );
  DFFSR oddBuffer_reg_46_ ( .D(n941), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[46]) );
  DFFSR oddBuffer_reg_45_ ( .D(n942), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[45]) );
  DFFSR oddBuffer_reg_44_ ( .D(n943), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[44]) );
  DFFSR oddBuffer_reg_43_ ( .D(n944), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[43]) );
  DFFSR oddBuffer_reg_42_ ( .D(n945), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[42]) );
  DFFSR oddBuffer_reg_41_ ( .D(n946), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[41]) );
  DFFSR oddBuffer_reg_40_ ( .D(n947), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[40]) );
  DFFSR oddBuffer_reg_63_ ( .D(n924), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[63]) );
  DFFSR oddBuffer_reg_62_ ( .D(n925), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[62]) );
  DFFSR oddBuffer_reg_61_ ( .D(n926), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[61]) );
  DFFSR oddBuffer_reg_60_ ( .D(n927), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[60]) );
  DFFSR oddBuffer_reg_59_ ( .D(n928), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[59]) );
  DFFSR oddBuffer_reg_58_ ( .D(n929), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[58]) );
  DFFSR oddBuffer_reg_57_ ( .D(n930), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[57]) );
  DFFSR oddBuffer_reg_56_ ( .D(n931), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[56]) );
  DFFSR oddBuffer_reg_54_ ( .D(n933), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[54]) );
  DFFSR oddBuffer_reg_53_ ( .D(n934), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[53]) );
  DFFSR oddBuffer_reg_52_ ( .D(n935), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[52]) );
  DFFSR oddBuffer_reg_27_ ( .D(n960), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[27]) );
  DFFSR oddBuffer_reg_25_ ( .D(n962), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[25]) );
  DFFSR oddBuffer_reg_24_ ( .D(n963), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[24]) );
  DFFSR oddBuffer_reg_23_ ( .D(n964), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[23]) );
  DFFSR oddBuffer_reg_22_ ( .D(n965), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[22]) );
  DFFSR oddBuffer_reg_21_ ( .D(n966), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[21]) );
  DFFSR oddBuffer_reg_20_ ( .D(n967), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[20]) );
  DFFSR oddBuffer_reg_19_ ( .D(n968), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[19]) );
  DFFSR oddBuffer_reg_18_ ( .D(n969), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[18]) );
  DFFSR oddBuffer_reg_17_ ( .D(n970), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[17]) );
  DFFSR oddBuffer_reg_16_ ( .D(n971), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[16]) );
  DFFSR oddBuffer_reg_15_ ( .D(n972), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[15]) );
  DFFSR oddBuffer_reg_13_ ( .D(n974), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[13]) );
  DFFSR oddBuffer_reg_12_ ( .D(n975), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[12]) );
  DFFSR oddBuffer_reg_11_ ( .D(n976), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[11]) );
  DFFSR oddBuffer_reg_10_ ( .D(n977), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[10]) );
  DFFSR oddBuffer_reg_9_ ( .D(n978), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[9]) );
  DFFSR oddBuffer_reg_8_ ( .D(n979), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[8]) );
  DFFSR oddBuffer_reg_7_ ( .D(n980), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[7]) );
  DFFSR oddBuffer_reg_6_ ( .D(n981), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[6]) );
  DFFSR oddBuffer_reg_5_ ( .D(n982), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[5]) );
  DFFSR oddBuffer_reg_4_ ( .D(n983), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[4]) );
  DFFSR oddBuffer_reg_39_ ( .D(n948), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[39]) );
  DFFSR oddBuffer_reg_38_ ( .D(n949), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[38]) );
  DFFSR oddBuffer_reg_37_ ( .D(n950), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[37]) );
  DFFSR oddBuffer_reg_36_ ( .D(n951), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[36]) );
  DFFSR oddBuffer_reg_35_ ( .D(n952), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[35]) );
  DFFSR oddBuffer_reg_34_ ( .D(n953), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[34]) );
  DFFSR oddBuffer_reg_33_ ( .D(n954), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[33]) );
  DFFSR oddBuffer_reg_32_ ( .D(n955), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[32]) );
  DFFSR oddBuffer_reg_31_ ( .D(n956), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[31]) );
  DFFSR oddBuffer_reg_30_ ( .D(n957), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[30]) );
  DFFSR oddBuffer_reg_29_ ( .D(n958), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[29]) );
  DFFSR oddBuffer_reg_28_ ( .D(n959), .CLK(clk), .R(n920), .S(1'b1), .Q(
        oddBuffer[28]) );
  AND2X1 U2 ( .A(n1), .B(n3), .Y(n1265) );
  OR2X1 U3 ( .A(n169), .B(n423), .Y(sub_111_aco_carry[1]) );
  OR2X1 U4 ( .A(n177), .B(n357), .Y(sub_131_aco_carry[1]) );
  OR2X1 U5 ( .A(sub_111_aco_carry[1]), .B(n345), .Y(sub_111_aco_carry[2]) );
  OR2X1 U6 ( .A(sub_131_aco_carry[1]), .B(n333), .Y(sub_131_aco_carry[2]) );
  OR2X1 U7 ( .A(sub_111_aco_carry[2]), .B(n421), .Y(sub_111_aco_carry[3]) );
  OR2X1 U8 ( .A(sub_131_aco_carry[2]), .B(n356), .Y(sub_131_aco_carry[3]) );
  OR2X1 U9 ( .A(sub_111_aco_carry[3]), .B(n420), .Y(sub_111_aco_carry[4]) );
  OR2X1 U10 ( .A(sub_131_aco_carry[3]), .B(n355), .Y(sub_131_aco_carry[4]) );
  OR2X1 U11 ( .A(sub_111_aco_carry[4]), .B(n358), .Y(sub_111_aco_carry[5]) );
  OR2X1 U12 ( .A(sub_131_aco_carry[4]), .B(n422), .Y(sub_131_aco_carry[5]) );
  OR2X1 U13 ( .A(sub_111_aco_carry[5]), .B(n334), .Y(sub_111_aco_carry[6]) );
  OR2X1 U14 ( .A(sub_131_aco_carry[5]), .B(n344), .Y(sub_131_aco_carry[6]) );
  OR2X1 U15 ( .A(sub_111_aco_carry[6]), .B(n419), .Y(sub_111_aco_carry[7]) );
  OR2X1 U16 ( .A(sub_131_aco_carry[6]), .B(n354), .Y(sub_131_aco_carry[7]) );
  AND2X1 U17 ( .A(n2), .B(n4), .Y(n1264) );
  OR2X1 U18 ( .A(n439), .B(n78), .Y(n1124) );
  BUFX2 U19 ( .A(n1261), .Y(n1) );
  BUFX2 U20 ( .A(n1263), .Y(n2) );
  BUFX2 U21 ( .A(n1260), .Y(n3) );
  BUFX2 U22 ( .A(n1262), .Y(n4) );
  AND2X1 U23 ( .A(n416), .B(n435), .Y(n1052) );
  INVX1 U24 ( .A(n1052), .Y(n5) );
  AND2X1 U25 ( .A(n406), .B(n434), .Y(n1053) );
  INVX1 U26 ( .A(n1053), .Y(n6) );
  AND2X1 U27 ( .A(n405), .B(n434), .Y(n1054) );
  INVX1 U28 ( .A(n1054), .Y(n7) );
  AND2X1 U29 ( .A(n404), .B(n434), .Y(n1055) );
  INVX1 U30 ( .A(n1055), .Y(n8) );
  AND2X1 U31 ( .A(n403), .B(n434), .Y(n1056) );
  INVX1 U32 ( .A(n1056), .Y(n9) );
  AND2X1 U33 ( .A(n402), .B(n434), .Y(n1057) );
  INVX1 U34 ( .A(n1057), .Y(n10) );
  AND2X1 U35 ( .A(n401), .B(n434), .Y(n1058) );
  INVX1 U36 ( .A(n1058), .Y(n11) );
  AND2X1 U37 ( .A(n400), .B(n435), .Y(n1059) );
  INVX1 U38 ( .A(n1059), .Y(n12) );
  AND2X1 U39 ( .A(n399), .B(n435), .Y(n1060) );
  INVX1 U40 ( .A(n1060), .Y(n13) );
  AND2X1 U41 ( .A(n398), .B(n434), .Y(n1061) );
  INVX1 U42 ( .A(n1061), .Y(n14) );
  AND2X1 U43 ( .A(n397), .B(n434), .Y(n1062) );
  INVX1 U44 ( .A(n1062), .Y(n15) );
  AND2X1 U45 ( .A(n415), .B(n435), .Y(n1063) );
  INVX1 U46 ( .A(n1063), .Y(n16) );
  AND2X1 U47 ( .A(n396), .B(n434), .Y(n1064) );
  INVX1 U48 ( .A(n1064), .Y(n17) );
  AND2X1 U49 ( .A(n395), .B(n434), .Y(n1065) );
  INVX1 U50 ( .A(n1065), .Y(n18) );
  AND2X1 U51 ( .A(n394), .B(n435), .Y(n1066) );
  INVX1 U52 ( .A(n1066), .Y(n19) );
  AND2X1 U53 ( .A(n393), .B(n434), .Y(n1067) );
  INVX1 U54 ( .A(n1067), .Y(n20) );
  AND2X1 U55 ( .A(n392), .B(n435), .Y(n1068) );
  INVX1 U56 ( .A(n1068), .Y(n21) );
  AND2X1 U57 ( .A(n391), .B(n435), .Y(n1069) );
  INVX1 U58 ( .A(n1069), .Y(n22) );
  AND2X1 U59 ( .A(n390), .B(n435), .Y(n1070) );
  INVX1 U60 ( .A(n1070), .Y(n23) );
  AND2X1 U61 ( .A(n389), .B(n435), .Y(n1071) );
  INVX1 U62 ( .A(n1071), .Y(n24) );
  AND2X1 U63 ( .A(n388), .B(n435), .Y(n1072) );
  INVX1 U64 ( .A(n1072), .Y(n25) );
  AND2X1 U65 ( .A(n387), .B(n435), .Y(n1073) );
  INVX1 U66 ( .A(n1073), .Y(n26) );
  AND2X1 U67 ( .A(n414), .B(n435), .Y(n1074) );
  INVX1 U68 ( .A(n1074), .Y(n27) );
  AND2X1 U69 ( .A(n386), .B(n435), .Y(n1075) );
  INVX1 U70 ( .A(n1075), .Y(n28) );
  AND2X1 U71 ( .A(n385), .B(n435), .Y(n1076) );
  INVX1 U72 ( .A(n1076), .Y(n29) );
  AND2X1 U73 ( .A(n384), .B(n435), .Y(n1077) );
  INVX1 U74 ( .A(n1077), .Y(n30) );
  AND2X1 U75 ( .A(n383), .B(n435), .Y(n1078) );
  INVX1 U76 ( .A(n1078), .Y(n31) );
  AND2X1 U77 ( .A(n382), .B(n435), .Y(n1079) );
  INVX1 U78 ( .A(n1079), .Y(n32) );
  AND2X1 U79 ( .A(n381), .B(n435), .Y(n1080) );
  INVX1 U80 ( .A(n1080), .Y(n33) );
  AND2X1 U81 ( .A(n380), .B(n436), .Y(n1081) );
  INVX1 U82 ( .A(n1081), .Y(n34) );
  AND2X1 U83 ( .A(n379), .B(n436), .Y(n1082) );
  INVX1 U84 ( .A(n1082), .Y(n35) );
  AND2X1 U85 ( .A(n378), .B(n436), .Y(n1083) );
  INVX1 U86 ( .A(n1083), .Y(n36) );
  AND2X1 U87 ( .A(n377), .B(n436), .Y(n1084) );
  INVX1 U88 ( .A(n1084), .Y(n37) );
  AND2X1 U89 ( .A(n413), .B(n436), .Y(n1085) );
  INVX1 U90 ( .A(n1085), .Y(n38) );
  AND2X1 U91 ( .A(n376), .B(n436), .Y(n1086) );
  INVX1 U92 ( .A(n1086), .Y(n39) );
  AND2X1 U93 ( .A(n375), .B(n436), .Y(n1087) );
  INVX1 U94 ( .A(n1087), .Y(n40) );
  AND2X1 U95 ( .A(n374), .B(n436), .Y(n1088) );
  INVX1 U96 ( .A(n1088), .Y(n41) );
  AND2X1 U97 ( .A(n373), .B(n436), .Y(n1089) );
  INVX1 U98 ( .A(n1089), .Y(n42) );
  AND2X1 U99 ( .A(n372), .B(n436), .Y(n1090) );
  INVX1 U100 ( .A(n1090), .Y(n43) );
  AND2X1 U101 ( .A(n371), .B(n436), .Y(n1091) );
  INVX1 U102 ( .A(n1091), .Y(n44) );
  AND2X1 U103 ( .A(n370), .B(n436), .Y(n1092) );
  INVX1 U104 ( .A(n1092), .Y(n45) );
  AND2X1 U105 ( .A(n369), .B(n436), .Y(n1093) );
  INVX1 U106 ( .A(n1093), .Y(n46) );
  AND2X1 U107 ( .A(n412), .B(n436), .Y(n1096) );
  INVX1 U108 ( .A(n1096), .Y(n47) );
  AND2X1 U109 ( .A(n368), .B(n436), .Y(n1103) );
  INVX1 U110 ( .A(n1103), .Y(n48) );
  AND2X1 U111 ( .A(n367), .B(n436), .Y(n1104) );
  INVX1 U112 ( .A(n1104), .Y(n49) );
  AND2X1 U113 ( .A(n366), .B(n436), .Y(n1105) );
  INVX1 U114 ( .A(n1105), .Y(n50) );
  AND2X1 U115 ( .A(n365), .B(n436), .Y(n1106) );
  INVX1 U116 ( .A(n1106), .Y(n51) );
  AND2X1 U117 ( .A(n411), .B(n431), .Y(n1107) );
  INVX1 U118 ( .A(n1107), .Y(n52) );
  AND2X1 U119 ( .A(n364), .B(n430), .Y(n1108) );
  INVX1 U120 ( .A(n1108), .Y(n53) );
  AND2X1 U121 ( .A(n363), .B(n433), .Y(n1109) );
  INVX1 U122 ( .A(n1109), .Y(n54) );
  AND2X1 U123 ( .A(n362), .B(n432), .Y(n1110) );
  INVX1 U124 ( .A(n1110), .Y(n55) );
  AND2X1 U125 ( .A(n361), .B(n431), .Y(n1111) );
  INVX1 U126 ( .A(n1111), .Y(n56) );
  AND2X1 U127 ( .A(n410), .B(n430), .Y(n1112) );
  INVX1 U128 ( .A(n1112), .Y(n57) );
  AND2X1 U129 ( .A(n409), .B(n433), .Y(n1113) );
  INVX1 U130 ( .A(n1113), .Y(n58) );
  AND2X1 U131 ( .A(n408), .B(n432), .Y(n1114) );
  INVX1 U132 ( .A(n1114), .Y(n59) );
  AND2X1 U133 ( .A(n407), .B(n431), .Y(n1115) );
  INVX1 U134 ( .A(n1115), .Y(n60) );
  AND2X1 U135 ( .A(n424), .B(dataIn[55]), .Y(n1136) );
  INVX1 U136 ( .A(n1136), .Y(n61) );
  AND2X1 U137 ( .A(n1127), .B(dataIn[51]), .Y(n1140) );
  INVX1 U138 ( .A(n1140), .Y(n62) );
  AND2X1 U139 ( .A(n1127), .B(dataIn[49]), .Y(n1142) );
  INVX1 U140 ( .A(n1142), .Y(n63) );
  AND2X1 U141 ( .A(n1127), .B(dataIn[26]), .Y(n1165) );
  INVX1 U142 ( .A(n1165), .Y(n64) );
  AND2X1 U143 ( .A(n1127), .B(dataIn[14]), .Y(n1177) );
  INVX1 U144 ( .A(n1177), .Y(n65) );
  AND2X1 U145 ( .A(dataIn[63]), .B(n1193), .Y(n1194) );
  INVX1 U146 ( .A(n1194), .Y(n66) );
  AND2X1 U147 ( .A(dataIn[62]), .B(n1193), .Y(n1195) );
  INVX1 U148 ( .A(n1195), .Y(n67) );
  AND2X1 U149 ( .A(dataIn[51]), .B(n1193), .Y(n1206) );
  INVX1 U150 ( .A(n1206), .Y(n68) );
  AND2X1 U151 ( .A(dataIn[50]), .B(n1193), .Y(n1207) );
  INVX1 U152 ( .A(n1207), .Y(n69) );
  AND2X1 U153 ( .A(dataIn[38]), .B(n1193), .Y(n1219) );
  INVX1 U154 ( .A(n1219), .Y(n70) );
  AND2X1 U155 ( .A(dataIn[37]), .B(n425), .Y(n1220) );
  INVX1 U156 ( .A(n1220), .Y(n71) );
  AND2X1 U157 ( .A(dataIn[36]), .B(n425), .Y(n1221) );
  INVX1 U158 ( .A(n1221), .Y(n72) );
  AND2X1 U159 ( .A(dataIn[26]), .B(n425), .Y(n1231) );
  INVX1 U160 ( .A(n1231), .Y(n73) );
  AND2X1 U161 ( .A(dataIn[24]), .B(n425), .Y(n1233) );
  INVX1 U162 ( .A(n1233), .Y(n74) );
  AND2X1 U163 ( .A(dataIn[14]), .B(n1193), .Y(n1243) );
  INVX1 U164 ( .A(n1243), .Y(n75) );
  AND2X1 U165 ( .A(dataIn[11]), .B(n1193), .Y(n1246) );
  INVX1 U166 ( .A(n1246), .Y(n76) );
  BUFX2 U167 ( .A(n1259), .Y(n77) );
  OR2X1 U168 ( .A(outputBufferGrant[0]), .B(outputBufferGrant[1]), .Y(n1126)
         );
  INVX1 U169 ( .A(n1126), .Y(n78) );
  INVX1 U170 ( .A(n1264), .Y(request[1]) );
  INVX1 U171 ( .A(n1265), .Y(request[0]) );
  INVX8 U172 ( .A(reset), .Y(n920) );
  AND2X1 U331 ( .A(n424), .B(dataIn[54]), .Y(n1137) );
  INVX1 U333 ( .A(n1137), .Y(n229) );
  AND2X1 U335 ( .A(n1127), .B(dataIn[50]), .Y(n1141) );
  INVX1 U337 ( .A(n1141), .Y(n230) );
  AND2X1 U339 ( .A(dataIn[61]), .B(n1193), .Y(n1196) );
  INVX1 U341 ( .A(n1196), .Y(n231) );
  AND2X1 U343 ( .A(dataIn[47]), .B(n1193), .Y(n1210) );
  INVX1 U345 ( .A(n1210), .Y(n232) );
  AND2X1 U347 ( .A(dataIn[35]), .B(n425), .Y(n1222) );
  INVX1 U349 ( .A(n1222), .Y(n233) );
  AND2X1 U351 ( .A(dataIn[23]), .B(n1193), .Y(n1234) );
  INVX1 U353 ( .A(n1234), .Y(n234) );
  AND2X1 U355 ( .A(dataIn[10]), .B(n1193), .Y(n1247) );
  INVX1 U357 ( .A(n1247), .Y(n235) );
  AND2X1 U359 ( .A(n1127), .B(dataIn[38]), .Y(n1153) );
  INVX1 U361 ( .A(n1153), .Y(n236) );
  AND2X1 U363 ( .A(n1127), .B(dataIn[25]), .Y(n1166) );
  INVX1 U365 ( .A(n1166), .Y(n237) );
  AND2X1 U367 ( .A(n1127), .B(dataIn[12]), .Y(n1179) );
  INVX1 U369 ( .A(n1179), .Y(n238) );
  AND2X1 U371 ( .A(dataIn[60]), .B(n1193), .Y(n1197) );
  INVX1 U373 ( .A(n1197), .Y(n239) );
  AND2X1 U375 ( .A(dataIn[46]), .B(n1193), .Y(n1211) );
  INVX1 U377 ( .A(n1211), .Y(n240) );
  AND2X1 U379 ( .A(dataIn[34]), .B(n425), .Y(n1223) );
  INVX1 U381 ( .A(n1223), .Y(n241) );
  AND2X1 U383 ( .A(dataIn[22]), .B(n1193), .Y(n1235) );
  INVX1 U385 ( .A(n1235), .Y(n242) );
  AND2X1 U387 ( .A(dataIn[9]), .B(n1193), .Y(n1248) );
  INVX1 U389 ( .A(n1248), .Y(n243) );
  AND2X1 U391 ( .A(n424), .B(dataIn[52]), .Y(n1139) );
  INVX1 U393 ( .A(n1139), .Y(n244) );
  AND2X1 U395 ( .A(n1127), .B(dataIn[37]), .Y(n1154) );
  INVX1 U397 ( .A(n1154), .Y(n245) );
  AND2X1 U399 ( .A(n1127), .B(dataIn[24]), .Y(n1167) );
  INVX1 U401 ( .A(n1167), .Y(n246) );
  AND2X1 U403 ( .A(n1127), .B(dataIn[11]), .Y(n1180) );
  INVX1 U405 ( .A(n1180), .Y(n247) );
  AND2X1 U407 ( .A(dataIn[59]), .B(n1193), .Y(n1198) );
  INVX1 U409 ( .A(n1198), .Y(n248) );
  AND2X1 U411 ( .A(dataIn[45]), .B(n1193), .Y(n1212) );
  INVX1 U413 ( .A(n1212), .Y(n249) );
  AND2X1 U415 ( .A(dataIn[33]), .B(n425), .Y(n1224) );
  INVX1 U417 ( .A(n1224), .Y(n250) );
  AND2X1 U419 ( .A(dataIn[21]), .B(n1193), .Y(n1236) );
  INVX1 U421 ( .A(n1236), .Y(n251) );
  AND2X1 U423 ( .A(dataIn[8]), .B(n1193), .Y(n1249) );
  INVX1 U425 ( .A(n1249), .Y(n252) );
  AND2X1 U427 ( .A(n424), .B(dataIn[63]), .Y(n1128) );
  INVX1 U429 ( .A(n1128), .Y(n253) );
  AND2X1 U431 ( .A(n1127), .B(dataIn[48]), .Y(n1143) );
  INVX1 U433 ( .A(n1143), .Y(n254) );
  AND2X1 U435 ( .A(n1127), .B(dataIn[36]), .Y(n1155) );
  INVX1 U437 ( .A(n1155), .Y(n255) );
  AND2X1 U439 ( .A(n1127), .B(dataIn[23]), .Y(n1168) );
  INVX1 U441 ( .A(n1168), .Y(n256) );
  AND2X1 U443 ( .A(n1127), .B(dataIn[10]), .Y(n1181) );
  INVX1 U445 ( .A(n1181), .Y(n257) );
  AND2X1 U447 ( .A(dataIn[58]), .B(n1193), .Y(n1199) );
  INVX1 U449 ( .A(n1199), .Y(n258) );
  AND2X1 U451 ( .A(dataIn[44]), .B(n1193), .Y(n1213) );
  INVX1 U453 ( .A(n1213), .Y(n259) );
  AND2X1 U455 ( .A(dataIn[32]), .B(n425), .Y(n1225) );
  INVX1 U457 ( .A(n1225), .Y(n260) );
  AND2X1 U459 ( .A(dataIn[20]), .B(n1193), .Y(n1237) );
  INVX1 U461 ( .A(n1237), .Y(n261) );
  AND2X1 U463 ( .A(dataIn[7]), .B(n1193), .Y(n1250) );
  INVX1 U465 ( .A(n1250), .Y(n262) );
  AND2X1 U467 ( .A(n424), .B(dataIn[62]), .Y(n1129) );
  INVX1 U469 ( .A(n1129), .Y(n263) );
  AND2X1 U471 ( .A(n1127), .B(dataIn[47]), .Y(n1144) );
  INVX1 U473 ( .A(n1144), .Y(n264) );
  AND2X1 U475 ( .A(n1127), .B(dataIn[35]), .Y(n1156) );
  INVX1 U477 ( .A(n1156), .Y(n265) );
  AND2X1 U479 ( .A(n1127), .B(dataIn[22]), .Y(n1169) );
  INVX1 U481 ( .A(n1169), .Y(n266) );
  AND2X1 U483 ( .A(n1127), .B(dataIn[9]), .Y(n1182) );
  INVX1 U485 ( .A(n1182), .Y(n267) );
  AND2X1 U487 ( .A(dataIn[57]), .B(n1193), .Y(n1200) );
  INVX1 U489 ( .A(n1200), .Y(n268) );
  AND2X1 U491 ( .A(dataIn[43]), .B(n1193), .Y(n1214) );
  INVX1 U493 ( .A(n1214), .Y(n269) );
  AND2X1 U495 ( .A(dataIn[31]), .B(n425), .Y(n1226) );
  INVX1 U497 ( .A(n1226), .Y(n270) );
  AND2X1 U499 ( .A(dataIn[19]), .B(n1193), .Y(n1238) );
  INVX1 U501 ( .A(n1238), .Y(n271) );
  AND2X1 U503 ( .A(dataIn[6]), .B(n1193), .Y(n1251) );
  INVX1 U505 ( .A(n1251), .Y(n272) );
  AND2X1 U507 ( .A(n424), .B(dataIn[61]), .Y(n1130) );
  INVX1 U509 ( .A(n1130), .Y(n273) );
  AND2X1 U511 ( .A(n1127), .B(dataIn[46]), .Y(n1145) );
  INVX1 U513 ( .A(n1145), .Y(n274) );
  AND2X1 U515 ( .A(n1127), .B(dataIn[34]), .Y(n1157) );
  INVX1 U517 ( .A(n1157), .Y(n275) );
  AND2X1 U519 ( .A(n1127), .B(dataIn[21]), .Y(n1170) );
  INVX1 U521 ( .A(n1170), .Y(n276) );
  AND2X1 U523 ( .A(n1127), .B(dataIn[8]), .Y(n1183) );
  INVX1 U525 ( .A(n1183), .Y(n277) );
  AND2X1 U527 ( .A(dataIn[55]), .B(n1193), .Y(n1202) );
  INVX1 U529 ( .A(n1202), .Y(n278) );
  AND2X1 U531 ( .A(dataIn[42]), .B(n1193), .Y(n1215) );
  INVX1 U533 ( .A(n1215), .Y(n279) );
  AND2X1 U535 ( .A(dataIn[30]), .B(n425), .Y(n1227) );
  INVX1 U537 ( .A(n1227), .Y(n280) );
  AND2X1 U539 ( .A(dataIn[18]), .B(n1193), .Y(n1239) );
  INVX1 U541 ( .A(n1239), .Y(n281) );
  AND2X1 U543 ( .A(dataIn[5]), .B(n1193), .Y(n1252) );
  INVX1 U545 ( .A(n1252), .Y(n282) );
  AND2X1 U547 ( .A(n424), .B(dataIn[60]), .Y(n1131) );
  INVX1 U549 ( .A(n1131), .Y(n283) );
  AND2X1 U551 ( .A(n1127), .B(dataIn[45]), .Y(n1146) );
  INVX1 U552 ( .A(n1146), .Y(n284) );
  AND2X1 U554 ( .A(n1127), .B(dataIn[33]), .Y(n1158) );
  INVX1 U556 ( .A(n1158), .Y(n285) );
  AND2X1 U557 ( .A(n1127), .B(dataIn[20]), .Y(n1171) );
  INVX1 U559 ( .A(n1171), .Y(n286) );
  AND2X1 U561 ( .A(n1127), .B(dataIn[7]), .Y(n1184) );
  INVX1 U563 ( .A(n1184), .Y(n287) );
  AND2X1 U565 ( .A(dataIn[54]), .B(n1193), .Y(n1203) );
  INVX1 U567 ( .A(n1203), .Y(n288) );
  AND2X1 U569 ( .A(dataIn[41]), .B(n1193), .Y(n1216) );
  INVX1 U571 ( .A(n1216), .Y(n289) );
  AND2X1 U573 ( .A(dataIn[29]), .B(n425), .Y(n1228) );
  INVX1 U575 ( .A(n1228), .Y(n290) );
  AND2X1 U577 ( .A(dataIn[17]), .B(n1193), .Y(n1240) );
  INVX1 U579 ( .A(n1240), .Y(n291) );
  AND2X1 U581 ( .A(dataIn[4]), .B(n1193), .Y(n1253) );
  INVX1 U583 ( .A(n1253), .Y(n292) );
  AND2X1 U585 ( .A(n424), .B(dataIn[59]), .Y(n1132) );
  INVX1 U587 ( .A(n1132), .Y(n293) );
  AND2X1 U595 ( .A(n1127), .B(dataIn[44]), .Y(n1147) );
  INVX1 U599 ( .A(n1147), .Y(n294) );
  AND2X1 U601 ( .A(n1127), .B(dataIn[32]), .Y(n1159) );
  INVX1 U603 ( .A(n1159), .Y(n295) );
  AND2X1 U605 ( .A(n1127), .B(dataIn[19]), .Y(n1172) );
  INVX1 U607 ( .A(n1172), .Y(n296) );
  AND2X1 U609 ( .A(n1127), .B(dataIn[6]), .Y(n1185) );
  INVX1 U611 ( .A(n1185), .Y(n297) );
  AND2X1 U613 ( .A(dataIn[56]), .B(n1193), .Y(n1201) );
  INVX1 U615 ( .A(n1201), .Y(n298) );
  AND2X1 U617 ( .A(dataIn[40]), .B(n1193), .Y(n1217) );
  INVX1 U619 ( .A(n1217), .Y(n299) );
  AND2X1 U621 ( .A(dataIn[28]), .B(n425), .Y(n1229) );
  INVX1 U623 ( .A(n1229), .Y(n300) );
  AND2X1 U625 ( .A(dataIn[16]), .B(n1193), .Y(n1241) );
  INVX1 U627 ( .A(n1241), .Y(n301) );
  AND2X1 U629 ( .A(dataIn[3]), .B(n1193), .Y(n1254) );
  INVX1 U631 ( .A(n1254), .Y(n302) );
  AND2X1 U633 ( .A(n424), .B(dataIn[58]), .Y(n1133) );
  INVX1 U635 ( .A(n1133), .Y(n303) );
  AND2X1 U637 ( .A(n1127), .B(dataIn[43]), .Y(n1148) );
  INVX1 U639 ( .A(n1148), .Y(n304) );
  AND2X1 U641 ( .A(n1127), .B(dataIn[31]), .Y(n1160) );
  INVX1 U643 ( .A(n1160), .Y(n305) );
  AND2X1 U645 ( .A(n1127), .B(dataIn[18]), .Y(n1173) );
  INVX1 U647 ( .A(n1173), .Y(n306) );
  AND2X1 U649 ( .A(n1127), .B(dataIn[5]), .Y(n1186) );
  INVX1 U651 ( .A(n1186), .Y(n307) );
  AND2X1 U653 ( .A(n805), .B(n804), .Y(n1120) );
  INVX1 U655 ( .A(n1120), .Y(n308) );
  AND2X1 U657 ( .A(n1119), .B(n1118), .Y(n169) );
  INVX1 U659 ( .A(n169), .Y(n309) );
  AND2X1 U661 ( .A(n865), .B(n864), .Y(n1117) );
  INVX1 U663 ( .A(n1117), .Y(n310) );
  AND2X1 U665 ( .A(dataIn[39]), .B(n1193), .Y(n1218) );
  INVX1 U667 ( .A(n1218), .Y(n311) );
  AND2X1 U669 ( .A(dataIn[27]), .B(n425), .Y(n1230) );
  INVX1 U671 ( .A(n1230), .Y(n312) );
  AND2X1 U673 ( .A(dataIn[15]), .B(n1193), .Y(n1242) );
  INVX1 U675 ( .A(n1242), .Y(n313) );
  AND2X1 U677 ( .A(dataIn[2]), .B(n1193), .Y(n1255) );
  INVX1 U679 ( .A(n1255), .Y(n314) );
  AND2X1 U681 ( .A(n424), .B(dataIn[57]), .Y(n1134) );
  INVX1 U682 ( .A(n1134), .Y(n315) );
  AND2X1 U683 ( .A(n1127), .B(dataIn[42]), .Y(n1149) );
  INVX1 U684 ( .A(n1149), .Y(n316) );
  AND2X1 U685 ( .A(n1127), .B(dataIn[30]), .Y(n1161) );
  INVX1 U686 ( .A(n1161), .Y(n317) );
  AND2X1 U687 ( .A(n1127), .B(dataIn[17]), .Y(n1174) );
  INVX1 U688 ( .A(n1174), .Y(n318) );
  AND2X1 U689 ( .A(n1127), .B(dataIn[3]), .Y(n1188) );
  INVX1 U690 ( .A(n1188), .Y(n319) );
  AND2X1 U691 ( .A(dataIn[53]), .B(n1193), .Y(n1204) );
  INVX1 U692 ( .A(n1204), .Y(n320) );
  AND2X1 U693 ( .A(n869), .B(n868), .Y(n1116) );
  INVX1 U694 ( .A(n1116), .Y(n321) );
  AND2X1 U695 ( .A(n1123), .B(n1122), .Y(n177) );
  INVX1 U696 ( .A(n177), .Y(n322) );
  AND2X1 U697 ( .A(n459), .B(n458), .Y(n1121) );
  INVX1 U698 ( .A(n1121), .Y(n323) );
  AND2X1 U699 ( .A(dataIn[13]), .B(n1193), .Y(n1244) );
  INVX1 U700 ( .A(n1244), .Y(n324) );
  AND2X1 U701 ( .A(dataIn[1]), .B(n1193), .Y(n1256) );
  INVX1 U702 ( .A(n1256), .Y(n325) );
  AND2X1 U703 ( .A(n424), .B(dataIn[53]), .Y(n1138) );
  INVX1 U704 ( .A(n1138), .Y(n326) );
  AND2X1 U705 ( .A(n1127), .B(dataIn[41]), .Y(n1150) );
  INVX1 U706 ( .A(n1150), .Y(n327) );
  AND2X1 U707 ( .A(n1127), .B(dataIn[29]), .Y(n1162) );
  INVX1 U708 ( .A(n1162), .Y(n328) );
  AND2X1 U709 ( .A(n1127), .B(dataIn[15]), .Y(n1176) );
  INVX1 U710 ( .A(n1176), .Y(n329) );
  AND2X1 U711 ( .A(n1127), .B(dataIn[2]), .Y(n1189) );
  INVX1 U712 ( .A(n1189), .Y(n330) );
  AND2X1 U713 ( .A(dataIn[52]), .B(n1193), .Y(n1205) );
  INVX1 U714 ( .A(n1205), .Y(n331) );
  AND2X1 U715 ( .A(dataIn[49]), .B(n1193), .Y(n1208) );
  INVX1 U716 ( .A(n1208), .Y(n332) );
  BUFX2 U717 ( .A(oddBuffer[49]), .Y(n333) );
  BUFX2 U718 ( .A(evenBuffer[53]), .Y(n334) );
  AND2X1 U719 ( .A(dataIn[25]), .B(n425), .Y(n1232) );
  INVX1 U720 ( .A(n1232), .Y(n335) );
  AND2X1 U721 ( .A(dataIn[12]), .B(n1193), .Y(n1245) );
  INVX1 U722 ( .A(n1245), .Y(n336) );
  AND2X1 U723 ( .A(dataIn[0]), .B(n1193), .Y(n1257) );
  INVX1 U724 ( .A(n1257), .Y(n337) );
  AND2X1 U725 ( .A(n424), .B(dataIn[56]), .Y(n1135) );
  INVX1 U726 ( .A(n1135), .Y(n338) );
  AND2X1 U727 ( .A(n1127), .B(dataIn[39]), .Y(n1152) );
  INVX1 U728 ( .A(n1152), .Y(n339) );
  AND2X1 U729 ( .A(n1127), .B(dataIn[27]), .Y(n1164) );
  INVX1 U730 ( .A(n1164), .Y(n340) );
  AND2X1 U731 ( .A(n1127), .B(dataIn[13]), .Y(n1178) );
  INVX1 U732 ( .A(n1178), .Y(n341) );
  AND2X1 U733 ( .A(n1127), .B(dataIn[1]), .Y(n1190) );
  INVX1 U734 ( .A(n1190), .Y(n342) );
  AND2X1 U735 ( .A(dataIn[48]), .B(n1193), .Y(n1209) );
  INVX1 U736 ( .A(n1209), .Y(n343) );
  BUFX2 U737 ( .A(oddBuffer[53]), .Y(n344) );
  BUFX2 U738 ( .A(evenBuffer[49]), .Y(n345) );
  AND2X1 U739 ( .A(n1127), .B(dataIn[40]), .Y(n1151) );
  INVX1 U740 ( .A(n1151), .Y(n346) );
  AND2X1 U741 ( .A(n1127), .B(dataIn[28]), .Y(n1163) );
  INVX1 U742 ( .A(n1163), .Y(n347) );
  AND2X1 U743 ( .A(n1127), .B(dataIn[16]), .Y(n1175) );
  INVX1 U744 ( .A(n1175), .Y(n348) );
  AND2X1 U745 ( .A(n1127), .B(dataIn[4]), .Y(n1187) );
  INVX1 U746 ( .A(n1187), .Y(n349) );
  AND2X1 U747 ( .A(n1127), .B(dataIn[0]), .Y(n1191) );
  INVX1 U748 ( .A(n1191), .Y(n350) );
  AND2X1 U749 ( .A(n434), .B(n1258), .Y(n1193) );
  INVX1 U750 ( .A(n1193), .Y(n351) );
  BUFX2 U751 ( .A(oddBuffer[55]), .Y(n352) );
  BUFX2 U752 ( .A(oddBufferFull), .Y(n353) );
  BUFX2 U753 ( .A(oddBuffer[54]), .Y(n354) );
  BUFX2 U754 ( .A(oddBuffer[51]), .Y(n355) );
  BUFX2 U755 ( .A(oddBuffer[50]), .Y(n356) );
  BUFX2 U756 ( .A(oddBuffer[48]), .Y(n357) );
  BUFX2 U757 ( .A(evenBuffer[52]), .Y(n358) );
  AND2X1 U758 ( .A(sendIn), .B(n434), .Y(n1125) );
  INVX1 U759 ( .A(n1125), .Y(n359) );
  AND2X1 U760 ( .A(n1192), .B(n439), .Y(n1127) );
  INVX1 U761 ( .A(n1127), .Y(n360) );
  BUFX2 U762 ( .A(oddBuffer[63]), .Y(n361) );
  BUFX2 U763 ( .A(oddBuffer[62]), .Y(n362) );
  BUFX2 U764 ( .A(oddBuffer[61]), .Y(n363) );
  BUFX2 U765 ( .A(oddBuffer[60]), .Y(n364) );
  BUFX2 U766 ( .A(oddBuffer[59]), .Y(n365) );
  BUFX2 U767 ( .A(oddBuffer[58]), .Y(n366) );
  BUFX2 U768 ( .A(oddBuffer[57]), .Y(n367) );
  BUFX2 U769 ( .A(oddBuffer[56]), .Y(n368) );
  BUFX2 U770 ( .A(oddBuffer[47]), .Y(n369) );
  BUFX2 U771 ( .A(oddBuffer[46]), .Y(n370) );
  BUFX2 U772 ( .A(oddBuffer[45]), .Y(n371) );
  BUFX2 U773 ( .A(oddBuffer[44]), .Y(n372) );
  BUFX2 U774 ( .A(oddBuffer[43]), .Y(n373) );
  BUFX2 U775 ( .A(oddBuffer[42]), .Y(n374) );
  BUFX2 U776 ( .A(oddBuffer[41]), .Y(n375) );
  BUFX2 U777 ( .A(oddBuffer[40]), .Y(n376) );
  BUFX2 U778 ( .A(oddBuffer[39]), .Y(n377) );
  BUFX2 U779 ( .A(oddBuffer[38]), .Y(n378) );
  BUFX2 U780 ( .A(oddBuffer[37]), .Y(n379) );
  BUFX2 U781 ( .A(oddBuffer[36]), .Y(n380) );
  BUFX2 U782 ( .A(oddBuffer[35]), .Y(n381) );
  BUFX2 U783 ( .A(oddBuffer[34]), .Y(n382) );
  BUFX2 U784 ( .A(oddBuffer[33]), .Y(n383) );
  BUFX2 U785 ( .A(oddBuffer[32]), .Y(n384) );
  BUFX2 U786 ( .A(oddBuffer[31]), .Y(n385) );
  BUFX2 U787 ( .A(oddBuffer[30]), .Y(n386) );
  BUFX2 U788 ( .A(oddBuffer[29]), .Y(n387) );
  BUFX2 U789 ( .A(oddBuffer[28]), .Y(n388) );
  BUFX2 U790 ( .A(oddBuffer[27]), .Y(n389) );
  BUFX2 U791 ( .A(oddBuffer[26]), .Y(n390) );
  BUFX2 U792 ( .A(oddBuffer[25]), .Y(n391) );
  BUFX2 U793 ( .A(oddBuffer[24]), .Y(n392) );
  BUFX2 U794 ( .A(oddBuffer[23]), .Y(n393) );
  BUFX2 U795 ( .A(oddBuffer[22]), .Y(n394) );
  BUFX2 U796 ( .A(oddBuffer[21]), .Y(n395) );
  BUFX2 U797 ( .A(oddBuffer[20]), .Y(n396) );
  BUFX2 U798 ( .A(oddBuffer[19]), .Y(n397) );
  BUFX2 U799 ( .A(oddBuffer[18]), .Y(n398) );
  BUFX2 U800 ( .A(oddBuffer[17]), .Y(n399) );
  BUFX2 U801 ( .A(oddBuffer[16]), .Y(n400) );
  BUFX2 U802 ( .A(oddBuffer[15]), .Y(n401) );
  BUFX2 U803 ( .A(oddBuffer[14]), .Y(n402) );
  BUFX2 U804 ( .A(oddBuffer[13]), .Y(n403) );
  BUFX2 U805 ( .A(oddBuffer[12]), .Y(n404) );
  BUFX2 U806 ( .A(oddBuffer[11]), .Y(n405) );
  BUFX2 U807 ( .A(oddBuffer[10]), .Y(n406) );
  BUFX2 U808 ( .A(oddBuffer[9]), .Y(n407) );
  BUFX2 U809 ( .A(oddBuffer[8]), .Y(n408) );
  BUFX2 U810 ( .A(oddBuffer[7]), .Y(n409) );
  BUFX2 U811 ( .A(oddBuffer[6]), .Y(n410) );
  BUFX2 U812 ( .A(oddBuffer[5]), .Y(n411) );
  BUFX2 U813 ( .A(oddBuffer[4]), .Y(n412) );
  BUFX2 U814 ( .A(oddBuffer[3]), .Y(n413) );
  BUFX2 U815 ( .A(oddBuffer[2]), .Y(n414) );
  BUFX2 U816 ( .A(oddBuffer[1]), .Y(n415) );
  BUFX2 U817 ( .A(oddBuffer[0]), .Y(n416) );
  BUFX2 U818 ( .A(evenBuffer[55]), .Y(n417) );
  BUFX2 U819 ( .A(evenBufferFull), .Y(n418) );
  BUFX2 U820 ( .A(evenBuffer[54]), .Y(n419) );
  BUFX2 U821 ( .A(evenBuffer[51]), .Y(n420) );
  BUFX2 U822 ( .A(evenBuffer[50]), .Y(n421) );
  BUFX2 U823 ( .A(oddBuffer[52]), .Y(n422) );
  BUFX2 U824 ( .A(evenBuffer[48]), .Y(n423) );
  INVX1 U825 ( .A(n438), .Y(n429) );
  INVX1 U826 ( .A(n437), .Y(n434) );
  INVX1 U827 ( .A(n439), .Y(n435) );
  INVX1 U828 ( .A(n439), .Y(n436) );
  INVX1 U829 ( .A(n437), .Y(n433) );
  INVX1 U830 ( .A(n437), .Y(n432) );
  INVX1 U831 ( .A(n438), .Y(n431) );
  INVX1 U832 ( .A(n438), .Y(n430) );
  INVX1 U833 ( .A(n351), .Y(n425) );
  INVX1 U834 ( .A(n360), .Y(n424) );
  INVX1 U835 ( .A(n426), .Y(n438) );
  INVX1 U836 ( .A(n426), .Y(n437) );
  INVX1 U837 ( .A(n428), .Y(n426) );
  INVX1 U838 ( .A(n427), .Y(n439) );
  INVX1 U839 ( .A(n428), .Y(n427) );
  INVX1 U840 ( .A(polarity), .Y(n428) );
  INVX1 U841 ( .A(n415), .Y(n854) );
  INVX1 U842 ( .A(n414), .Y(n853) );
  INVX1 U843 ( .A(n413), .Y(n852) );
  INVX1 U844 ( .A(n412), .Y(n851) );
  INVX1 U845 ( .A(n411), .Y(n850) );
  INVX1 U846 ( .A(n410), .Y(n849) );
  INVX1 U847 ( .A(n409), .Y(n848) );
  INVX1 U848 ( .A(n408), .Y(n847) );
  INVX1 U849 ( .A(n407), .Y(n846) );
  INVX1 U850 ( .A(n406), .Y(n845) );
  INVX1 U851 ( .A(n405), .Y(n844) );
  INVX1 U852 ( .A(n404), .Y(n843) );
  INVX1 U853 ( .A(n403), .Y(n842) );
  INVX1 U854 ( .A(n402), .Y(n841) );
  INVX1 U855 ( .A(n401), .Y(n840) );
  INVX1 U856 ( .A(n400), .Y(n839) );
  INVX1 U857 ( .A(n399), .Y(n838) );
  INVX1 U858 ( .A(n398), .Y(n837) );
  INVX1 U859 ( .A(n397), .Y(n836) );
  INVX1 U860 ( .A(n396), .Y(n835) );
  INVX1 U861 ( .A(n395), .Y(n834) );
  INVX1 U862 ( .A(n394), .Y(n833) );
  INVX1 U863 ( .A(n393), .Y(n832) );
  INVX1 U864 ( .A(n392), .Y(n831) );
  INVX1 U865 ( .A(n391), .Y(n830) );
  INVX1 U866 ( .A(n390), .Y(n829) );
  INVX1 U867 ( .A(n389), .Y(n828) );
  INVX1 U868 ( .A(n388), .Y(n827) );
  INVX1 U869 ( .A(n387), .Y(n826) );
  INVX1 U870 ( .A(n386), .Y(n825) );
  INVX1 U871 ( .A(n385), .Y(n824) );
  INVX1 U872 ( .A(n384), .Y(n823) );
  INVX1 U873 ( .A(n383), .Y(n822) );
  INVX1 U874 ( .A(n382), .Y(n821) );
  INVX1 U875 ( .A(n381), .Y(n820) );
  INVX1 U876 ( .A(n380), .Y(n819) );
  INVX1 U877 ( .A(n379), .Y(n818) );
  INVX1 U878 ( .A(n378), .Y(n817) );
  INVX1 U879 ( .A(n377), .Y(n816) );
  INVX1 U880 ( .A(n376), .Y(n815) );
  INVX1 U881 ( .A(n375), .Y(n814) );
  INVX1 U882 ( .A(n374), .Y(n813) );
  INVX1 U883 ( .A(n373), .Y(n812) );
  INVX1 U884 ( .A(n372), .Y(n811) );
  INVX1 U885 ( .A(n371), .Y(n810) );
  INVX1 U886 ( .A(n370), .Y(n809) );
  INVX1 U887 ( .A(n369), .Y(n808) );
  INVX1 U888 ( .A(n357), .Y(n807) );
  INVX1 U889 ( .A(n333), .Y(n806) );
  INVX1 U890 ( .A(n422), .Y(n803) );
  INVX1 U891 ( .A(n334), .Y(n866) );
  INVX1 U892 ( .A(n416), .Y(n855) );
  INVX1 U893 ( .A(n344), .Y(n802) );
  INVX1 U894 ( .A(n368), .Y(n457) );
  INVX1 U895 ( .A(n367), .Y(n456) );
  INVX1 U896 ( .A(n366), .Y(n455) );
  INVX1 U897 ( .A(n365), .Y(n454) );
  INVX1 U898 ( .A(n364), .Y(n453) );
  INVX1 U899 ( .A(n363), .Y(n452) );
  INVX1 U900 ( .A(n362), .Y(n451) );
  INVX1 U901 ( .A(n361), .Y(n450) );
  INVX1 U902 ( .A(n423), .Y(n871) );
  INVX1 U903 ( .A(n345), .Y(n870) );
  INVX1 U904 ( .A(n358), .Y(n867) );
  INVX1 U905 ( .A(n1094), .Y(dataOut[48]) );
  INVX1 U906 ( .A(n1095), .Y(dataOut[49]) );
  INVX1 U907 ( .A(n1097), .Y(dataOut[50]) );
  INVX1 U908 ( .A(n1098), .Y(dataOut[51]) );
  INVX1 U909 ( .A(n1099), .Y(dataOut[52]) );
  INVX1 U910 ( .A(n1100), .Y(dataOut[53]) );
  INVX1 U911 ( .A(n1101), .Y(dataOut[54]) );
  INVX1 U912 ( .A(n1102), .Y(dataOut[55]) );
  INVX1 U913 ( .A(n356), .Y(n805) );
  INVX1 U914 ( .A(n354), .Y(n459) );
  INVX1 U915 ( .A(n421), .Y(n869) );
  INVX1 U916 ( .A(n419), .Y(n865) );
  INVX1 U917 ( .A(n355), .Y(n804) );
  INVX1 U918 ( .A(n420), .Y(n868) );
  INVX1 U919 ( .A(n418), .Y(n449) );
  INVX1 U920 ( .A(n353), .Y(n448) );
  INVX1 U921 ( .A(n352), .Y(n458) );
  INVX1 U922 ( .A(n417), .Y(n864) );
  INVX1 U923 ( .A(sendIn), .Y(n921) );
  INVX1 U924 ( .A(evenBuffer[0]), .Y(n919) );
  INVX1 U925 ( .A(evenBuffer[1]), .Y(n918) );
  INVX1 U926 ( .A(evenBuffer[2]), .Y(n917) );
  INVX1 U927 ( .A(evenBuffer[3]), .Y(n916) );
  INVX1 U928 ( .A(evenBuffer[4]), .Y(n915) );
  INVX1 U929 ( .A(evenBuffer[5]), .Y(n914) );
  INVX1 U930 ( .A(evenBuffer[6]), .Y(n913) );
  INVX1 U931 ( .A(evenBuffer[7]), .Y(n912) );
  INVX1 U932 ( .A(evenBuffer[8]), .Y(n911) );
  INVX1 U933 ( .A(evenBuffer[9]), .Y(n910) );
  INVX1 U934 ( .A(evenBuffer[10]), .Y(n909) );
  INVX1 U935 ( .A(evenBuffer[11]), .Y(n908) );
  INVX1 U936 ( .A(evenBuffer[12]), .Y(n907) );
  INVX1 U937 ( .A(evenBuffer[13]), .Y(n906) );
  INVX1 U938 ( .A(evenBuffer[14]), .Y(n905) );
  INVX1 U939 ( .A(evenBuffer[15]), .Y(n904) );
  INVX1 U940 ( .A(evenBuffer[16]), .Y(n903) );
  INVX1 U941 ( .A(evenBuffer[17]), .Y(n902) );
  INVX1 U942 ( .A(evenBuffer[18]), .Y(n901) );
  INVX1 U943 ( .A(evenBuffer[19]), .Y(n900) );
  INVX1 U944 ( .A(evenBuffer[20]), .Y(n899) );
  INVX1 U945 ( .A(evenBuffer[21]), .Y(n898) );
  INVX1 U946 ( .A(evenBuffer[22]), .Y(n897) );
  INVX1 U947 ( .A(evenBuffer[23]), .Y(n896) );
  INVX1 U948 ( .A(evenBuffer[24]), .Y(n895) );
  INVX1 U949 ( .A(evenBuffer[25]), .Y(n894) );
  INVX1 U950 ( .A(evenBuffer[26]), .Y(n893) );
  INVX1 U951 ( .A(evenBuffer[27]), .Y(n892) );
  INVX1 U952 ( .A(evenBuffer[28]), .Y(n891) );
  INVX1 U953 ( .A(evenBuffer[29]), .Y(n890) );
  INVX1 U954 ( .A(evenBuffer[30]), .Y(n889) );
  INVX1 U955 ( .A(evenBuffer[31]), .Y(n888) );
  INVX1 U956 ( .A(evenBuffer[32]), .Y(n887) );
  INVX1 U957 ( .A(evenBuffer[33]), .Y(n886) );
  INVX1 U958 ( .A(evenBuffer[34]), .Y(n885) );
  INVX1 U959 ( .A(evenBuffer[35]), .Y(n884) );
  INVX1 U960 ( .A(evenBuffer[36]), .Y(n883) );
  INVX1 U961 ( .A(evenBuffer[37]), .Y(n882) );
  INVX1 U962 ( .A(evenBuffer[38]), .Y(n881) );
  INVX1 U963 ( .A(evenBuffer[39]), .Y(n880) );
  INVX1 U964 ( .A(evenBuffer[40]), .Y(n879) );
  INVX1 U965 ( .A(evenBuffer[41]), .Y(n878) );
  INVX1 U966 ( .A(evenBuffer[42]), .Y(n877) );
  INVX1 U967 ( .A(evenBuffer[43]), .Y(n876) );
  INVX1 U968 ( .A(evenBuffer[44]), .Y(n875) );
  INVX1 U969 ( .A(evenBuffer[45]), .Y(n874) );
  INVX1 U970 ( .A(evenBuffer[46]), .Y(n873) );
  INVX1 U971 ( .A(evenBuffer[47]), .Y(n872) );
  INVX1 U972 ( .A(evenBuffer[56]), .Y(n863) );
  INVX1 U973 ( .A(evenBuffer[57]), .Y(n862) );
  INVX1 U974 ( .A(evenBuffer[58]), .Y(n861) );
  INVX1 U975 ( .A(evenBuffer[59]), .Y(n860) );
  INVX1 U976 ( .A(evenBuffer[60]), .Y(n859) );
  INVX1 U977 ( .A(evenBuffer[61]), .Y(n858) );
  INVX1 U978 ( .A(evenBuffer[62]), .Y(n857) );
  INVX1 U979 ( .A(evenBuffer[63]), .Y(n856) );
  XNOR2X1 U980 ( .A(n352), .B(sub_131_aco_carry[7]), .Y(n159) );
  XNOR2X1 U981 ( .A(n354), .B(sub_131_aco_carry[6]), .Y(n158) );
  XNOR2X1 U982 ( .A(n344), .B(sub_131_aco_carry[5]), .Y(n157) );
  XNOR2X1 U983 ( .A(n422), .B(sub_131_aco_carry[4]), .Y(n156) );
  XNOR2X1 U984 ( .A(n355), .B(sub_131_aco_carry[3]), .Y(n155) );
  XNOR2X1 U985 ( .A(n356), .B(sub_131_aco_carry[2]), .Y(n154) );
  XNOR2X1 U986 ( .A(n333), .B(sub_131_aco_carry[1]), .Y(n153) );
  XNOR2X1 U987 ( .A(n357), .B(n177), .Y(n152) );
  XNOR2X1 U988 ( .A(n417), .B(sub_111_aco_carry[7]), .Y(n147) );
  XNOR2X1 U989 ( .A(n419), .B(sub_111_aco_carry[6]), .Y(n146) );
  XNOR2X1 U990 ( .A(n334), .B(sub_111_aco_carry[5]), .Y(n145) );
  XNOR2X1 U991 ( .A(n358), .B(sub_111_aco_carry[4]), .Y(n144) );
  XNOR2X1 U992 ( .A(n420), .B(sub_111_aco_carry[3]), .Y(n143) );
  XNOR2X1 U993 ( .A(n421), .B(sub_111_aco_carry[2]), .Y(n142) );
  XNOR2X1 U994 ( .A(n345), .B(sub_111_aco_carry[1]), .Y(n141) );
  XNOR2X1 U995 ( .A(n423), .B(n169), .Y(n140) );
endmodule


module inputBuffer_PE1 ( clk, reset, polarity, sendIn, readyIn, dataIn, 
        dataOut, request, outputBufferGrant );
  input [63:0] dataIn;
  output [63:0] dataOut;
  output [1:0] request;
  input [1:0] outputBufferGrant;
  input clk, reset, polarity, sendIn;
  output readyIn;
  wire   n927, n928, evenBufferFull, oddBufferFull, n139, n140, n141, n142,
         n143, n144, n145, n146, n150, n151, n152, n153, n154, n155, n156,
         n157, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n130, n132, n133,
         n134, n135, n136, n137, n138, n147, n148, n149, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926;
  wire   [63:0] evenBuffer;
  wire   [63:0] oddBuffer;

  DFFSR oddBufferFull_reg ( .D(n616), .CLK(clk), .R(n749), .S(1'b1), .Q(
        oddBufferFull) );
  DFFSR evenBufferFull_reg ( .D(n615), .CLK(clk), .R(n750), .S(1'b1), .Q(
        evenBufferFull) );
  DFFSR oddBuffer_reg_63_ ( .D(n614), .CLK(clk), .R(n750), .S(1'b1), .Q(
        oddBuffer[63]) );
  DFFSR oddBuffer_reg_62_ ( .D(n613), .CLK(clk), .R(n749), .S(1'b1), .Q(
        oddBuffer[62]) );
  DFFSR oddBuffer_reg_61_ ( .D(n612), .CLK(clk), .R(n750), .S(1'b1), .Q(
        oddBuffer[61]) );
  DFFSR oddBuffer_reg_60_ ( .D(n611), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[60]) );
  DFFSR oddBuffer_reg_59_ ( .D(n610), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[59]) );
  DFFSR oddBuffer_reg_58_ ( .D(n609), .CLK(clk), .R(n750), .S(1'b1), .Q(
        oddBuffer[58]) );
  DFFSR oddBuffer_reg_57_ ( .D(n608), .CLK(clk), .R(n750), .S(1'b1), .Q(
        oddBuffer[57]) );
  DFFSR oddBuffer_reg_56_ ( .D(n607), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[56]) );
  DFFSR oddBuffer_reg_55_ ( .D(n606), .CLK(clk), .R(n750), .S(1'b1), .Q(
        oddBuffer[55]) );
  DFFSR oddBuffer_reg_54_ ( .D(n605), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[54]) );
  DFFSR oddBuffer_reg_53_ ( .D(n604), .CLK(clk), .R(n749), .S(1'b1), .Q(
        oddBuffer[53]) );
  DFFSR oddBuffer_reg_52_ ( .D(n603), .CLK(clk), .R(n749), .S(1'b1), .Q(
        oddBuffer[52]) );
  DFFSR oddBuffer_reg_51_ ( .D(n602), .CLK(clk), .R(n749), .S(1'b1), .Q(
        oddBuffer[51]) );
  DFFSR oddBuffer_reg_50_ ( .D(n601), .CLK(clk), .R(n749), .S(1'b1), .Q(
        oddBuffer[50]) );
  DFFSR oddBuffer_reg_49_ ( .D(n600), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[49]) );
  DFFSR oddBuffer_reg_48_ ( .D(n599), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[48]) );
  DFFSR oddBuffer_reg_47_ ( .D(n598), .CLK(clk), .R(n750), .S(1'b1), .Q(
        oddBuffer[47]) );
  DFFSR oddBuffer_reg_46_ ( .D(n597), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[46]) );
  DFFSR oddBuffer_reg_45_ ( .D(n596), .CLK(clk), .R(n750), .S(1'b1), .Q(
        oddBuffer[45]) );
  DFFSR oddBuffer_reg_44_ ( .D(n595), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[44]) );
  DFFSR oddBuffer_reg_43_ ( .D(n594), .CLK(clk), .R(n750), .S(1'b1), .Q(
        oddBuffer[43]) );
  DFFSR oddBuffer_reg_42_ ( .D(n593), .CLK(clk), .R(n750), .S(1'b1), .Q(
        oddBuffer[42]) );
  DFFSR oddBuffer_reg_41_ ( .D(n592), .CLK(clk), .R(n750), .S(1'b1), .Q(
        oddBuffer[41]) );
  DFFSR oddBuffer_reg_40_ ( .D(n591), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[40]) );
  DFFSR oddBuffer_reg_39_ ( .D(n590), .CLK(clk), .R(n749), .S(1'b1), .Q(
        oddBuffer[39]) );
  DFFSR oddBuffer_reg_38_ ( .D(n589), .CLK(clk), .R(n750), .S(1'b1), .Q(
        oddBuffer[38]) );
  DFFSR oddBuffer_reg_37_ ( .D(n588), .CLK(clk), .R(n749), .S(1'b1), .Q(
        oddBuffer[37]) );
  DFFSR oddBuffer_reg_36_ ( .D(n587), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[36]) );
  DFFSR oddBuffer_reg_35_ ( .D(n586), .CLK(clk), .R(n750), .S(1'b1), .Q(
        oddBuffer[35]) );
  DFFSR oddBuffer_reg_34_ ( .D(n585), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[34]) );
  DFFSR oddBuffer_reg_33_ ( .D(n584), .CLK(clk), .R(n750), .S(1'b1), .Q(
        oddBuffer[33]) );
  DFFSR oddBuffer_reg_32_ ( .D(n583), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[32]) );
  DFFSR oddBuffer_reg_31_ ( .D(n582), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[31]) );
  DFFSR oddBuffer_reg_30_ ( .D(n581), .CLK(clk), .R(n750), .S(1'b1), .Q(
        oddBuffer[30]) );
  DFFSR oddBuffer_reg_29_ ( .D(n580), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[29]) );
  DFFSR oddBuffer_reg_28_ ( .D(n579), .CLK(clk), .R(n750), .S(1'b1), .Q(
        oddBuffer[28]) );
  DFFSR oddBuffer_reg_27_ ( .D(n578), .CLK(clk), .R(n749), .S(1'b1), .Q(
        oddBuffer[27]) );
  DFFSR oddBuffer_reg_26_ ( .D(n577), .CLK(clk), .R(n749), .S(1'b1), .Q(
        oddBuffer[26]) );
  DFFSR oddBuffer_reg_25_ ( .D(n576), .CLK(clk), .R(n749), .S(1'b1), .Q(
        oddBuffer[25]) );
  DFFSR oddBuffer_reg_24_ ( .D(n575), .CLK(clk), .R(n749), .S(1'b1), .Q(
        oddBuffer[24]) );
  DFFSR oddBuffer_reg_23_ ( .D(n574), .CLK(clk), .R(n750), .S(1'b1), .Q(
        oddBuffer[23]) );
  DFFSR oddBuffer_reg_22_ ( .D(n573), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[22]) );
  DFFSR oddBuffer_reg_21_ ( .D(n572), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[21]) );
  DFFSR oddBuffer_reg_20_ ( .D(n571), .CLK(clk), .R(n749), .S(1'b1), .Q(
        oddBuffer[20]) );
  DFFSR oddBuffer_reg_19_ ( .D(n570), .CLK(clk), .R(n749), .S(1'b1), .Q(
        oddBuffer[19]) );
  DFFSR oddBuffer_reg_18_ ( .D(n569), .CLK(clk), .R(n749), .S(1'b1), .Q(
        oddBuffer[18]) );
  DFFSR oddBuffer_reg_17_ ( .D(n568), .CLK(clk), .R(n750), .S(1'b1), .Q(
        oddBuffer[17]) );
  DFFSR oddBuffer_reg_16_ ( .D(n567), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[16]) );
  DFFSR oddBuffer_reg_15_ ( .D(n566), .CLK(clk), .R(n749), .S(1'b1), .Q(
        oddBuffer[15]) );
  DFFSR oddBuffer_reg_14_ ( .D(n565), .CLK(clk), .R(n750), .S(1'b1), .Q(
        oddBuffer[14]) );
  DFFSR oddBuffer_reg_13_ ( .D(n564), .CLK(clk), .R(n750), .S(1'b1), .Q(
        oddBuffer[13]) );
  DFFSR oddBuffer_reg_12_ ( .D(n563), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[12]) );
  DFFSR oddBuffer_reg_11_ ( .D(n562), .CLK(clk), .R(n749), .S(1'b1), .Q(
        oddBuffer[11]) );
  DFFSR oddBuffer_reg_10_ ( .D(n561), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[10]) );
  DFFSR oddBuffer_reg_9_ ( .D(n560), .CLK(clk), .R(n750), .S(1'b1), .Q(
        oddBuffer[9]) );
  DFFSR oddBuffer_reg_8_ ( .D(n559), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[8]) );
  DFFSR oddBuffer_reg_7_ ( .D(n558), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[7]) );
  DFFSR oddBuffer_reg_6_ ( .D(n557), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[6]) );
  DFFSR oddBuffer_reg_5_ ( .D(n556), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[5]) );
  DFFSR oddBuffer_reg_4_ ( .D(n555), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[4]) );
  DFFSR oddBuffer_reg_3_ ( .D(n554), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[3]) );
  DFFSR oddBuffer_reg_2_ ( .D(n553), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[2]) );
  DFFSR oddBuffer_reg_1_ ( .D(n552), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[1]) );
  DFFSR oddBuffer_reg_0_ ( .D(n551), .CLK(clk), .R(n751), .S(1'b1), .Q(
        oddBuffer[0]) );
  DFFSR evenBuffer_reg_63_ ( .D(n550), .CLK(clk), .R(n751), .S(1'b1), .Q(
        evenBuffer[63]) );
  DFFSR evenBuffer_reg_62_ ( .D(n549), .CLK(clk), .R(n751), .S(1'b1), .Q(
        evenBuffer[62]) );
  DFFSR evenBuffer_reg_61_ ( .D(n548), .CLK(clk), .R(n751), .S(1'b1), .Q(
        evenBuffer[61]) );
  DFFSR evenBuffer_reg_60_ ( .D(n547), .CLK(clk), .R(n751), .S(1'b1), .Q(
        evenBuffer[60]) );
  DFFSR evenBuffer_reg_59_ ( .D(n546), .CLK(clk), .R(n750), .S(1'b1), .Q(
        evenBuffer[59]) );
  DFFSR evenBuffer_reg_58_ ( .D(n545), .CLK(clk), .R(n749), .S(1'b1), .Q(
        evenBuffer[58]) );
  DFFSR evenBuffer_reg_57_ ( .D(n544), .CLK(clk), .R(n751), .S(1'b1), .Q(
        evenBuffer[57]) );
  DFFSR evenBuffer_reg_56_ ( .D(n543), .CLK(clk), .R(n750), .S(1'b1), .Q(
        evenBuffer[56]) );
  DFFSR evenBuffer_reg_55_ ( .D(n789), .CLK(clk), .R(n750), .S(1'b1), .Q(
        evenBuffer[55]) );
  DFFSR evenBuffer_reg_54_ ( .D(n790), .CLK(clk), .R(n749), .S(1'b1), .Q(
        evenBuffer[54]) );
  DFFSR evenBuffer_reg_53_ ( .D(n791), .CLK(clk), .R(n751), .S(1'b1), .Q(
        evenBuffer[53]) );
  DFFSR evenBuffer_reg_52_ ( .D(n792), .CLK(clk), .R(n751), .S(1'b1), .Q(
        evenBuffer[52]) );
  DFFSR evenBuffer_reg_51_ ( .D(n793), .CLK(clk), .R(n749), .S(1'b1), .Q(
        evenBuffer[51]) );
  DFFSR evenBuffer_reg_50_ ( .D(n794), .CLK(clk), .R(n750), .S(1'b1), .Q(
        evenBuffer[50]) );
  DFFSR evenBuffer_reg_49_ ( .D(n795), .CLK(clk), .R(n749), .S(1'b1), .Q(
        evenBuffer[49]) );
  DFFSR evenBuffer_reg_48_ ( .D(n796), .CLK(clk), .R(n751), .S(1'b1), .Q(
        evenBuffer[48]) );
  DFFSR evenBuffer_reg_47_ ( .D(n542), .CLK(clk), .R(n751), .S(1'b1), .Q(
        evenBuffer[47]) );
  DFFSR evenBuffer_reg_46_ ( .D(n541), .CLK(clk), .R(n750), .S(1'b1), .Q(
        evenBuffer[46]) );
  DFFSR evenBuffer_reg_45_ ( .D(n540), .CLK(clk), .R(n749), .S(1'b1), .Q(
        evenBuffer[45]) );
  DFFSR evenBuffer_reg_44_ ( .D(n539), .CLK(clk), .R(n749), .S(1'b1), .Q(
        evenBuffer[44]) );
  DFFSR evenBuffer_reg_43_ ( .D(n538), .CLK(clk), .R(n749), .S(1'b1), .Q(
        evenBuffer[43]) );
  DFFSR evenBuffer_reg_42_ ( .D(n537), .CLK(clk), .R(n751), .S(1'b1), .Q(
        evenBuffer[42]) );
  DFFSR evenBuffer_reg_41_ ( .D(n536), .CLK(clk), .R(n750), .S(1'b1), .Q(
        evenBuffer[41]) );
  DFFSR evenBuffer_reg_40_ ( .D(n535), .CLK(clk), .R(n751), .S(1'b1), .Q(
        evenBuffer[40]) );
  DFFSR evenBuffer_reg_39_ ( .D(n534), .CLK(clk), .R(n749), .S(1'b1), .Q(
        evenBuffer[39]) );
  DFFSR evenBuffer_reg_38_ ( .D(n533), .CLK(clk), .R(n750), .S(1'b1), .Q(
        evenBuffer[38]) );
  DFFSR evenBuffer_reg_37_ ( .D(n532), .CLK(clk), .R(n749), .S(1'b1), .Q(
        evenBuffer[37]) );
  DFFSR evenBuffer_reg_36_ ( .D(n531), .CLK(clk), .R(n749), .S(1'b1), .Q(
        evenBuffer[36]) );
  DFFSR evenBuffer_reg_35_ ( .D(n530), .CLK(clk), .R(n750), .S(1'b1), .Q(
        evenBuffer[35]) );
  DFFSR evenBuffer_reg_34_ ( .D(n529), .CLK(clk), .R(n749), .S(1'b1), .Q(
        evenBuffer[34]) );
  DFFSR evenBuffer_reg_33_ ( .D(n528), .CLK(clk), .R(n751), .S(1'b1), .Q(
        evenBuffer[33]) );
  DFFSR evenBuffer_reg_32_ ( .D(n527), .CLK(clk), .R(n750), .S(1'b1), .Q(
        evenBuffer[32]) );
  DFFSR evenBuffer_reg_31_ ( .D(n526), .CLK(clk), .R(n749), .S(1'b1), .Q(
        evenBuffer[31]) );
  DFFSR evenBuffer_reg_30_ ( .D(n525), .CLK(clk), .R(n751), .S(1'b1), .Q(
        evenBuffer[30]) );
  DFFSR evenBuffer_reg_29_ ( .D(n524), .CLK(clk), .R(n750), .S(1'b1), .Q(
        evenBuffer[29]) );
  DFFSR evenBuffer_reg_28_ ( .D(n523), .CLK(clk), .R(n749), .S(1'b1), .Q(
        evenBuffer[28]) );
  DFFSR evenBuffer_reg_27_ ( .D(n522), .CLK(clk), .R(n751), .S(1'b1), .Q(
        evenBuffer[27]) );
  DFFSR evenBuffer_reg_26_ ( .D(n521), .CLK(clk), .R(n750), .S(1'b1), .Q(
        evenBuffer[26]) );
  DFFSR evenBuffer_reg_25_ ( .D(n520), .CLK(clk), .R(n749), .S(1'b1), .Q(
        evenBuffer[25]) );
  DFFSR evenBuffer_reg_24_ ( .D(n519), .CLK(clk), .R(n751), .S(1'b1), .Q(
        evenBuffer[24]) );
  DFFSR evenBuffer_reg_23_ ( .D(n518), .CLK(clk), .R(n750), .S(1'b1), .Q(
        evenBuffer[23]) );
  DFFSR evenBuffer_reg_22_ ( .D(n517), .CLK(clk), .R(n750), .S(1'b1), .Q(
        evenBuffer[22]) );
  DFFSR evenBuffer_reg_21_ ( .D(n516), .CLK(clk), .R(n750), .S(1'b1), .Q(
        evenBuffer[21]) );
  DFFSR evenBuffer_reg_20_ ( .D(n515), .CLK(clk), .R(n750), .S(1'b1), .Q(
        evenBuffer[20]) );
  DFFSR evenBuffer_reg_19_ ( .D(n514), .CLK(clk), .R(n750), .S(1'b1), .Q(
        evenBuffer[19]) );
  DFFSR evenBuffer_reg_18_ ( .D(n513), .CLK(clk), .R(n750), .S(1'b1), .Q(
        evenBuffer[18]) );
  DFFSR evenBuffer_reg_17_ ( .D(n512), .CLK(clk), .R(n750), .S(1'b1), .Q(
        evenBuffer[17]) );
  DFFSR evenBuffer_reg_16_ ( .D(n511), .CLK(clk), .R(n750), .S(1'b1), .Q(
        evenBuffer[16]) );
  DFFSR evenBuffer_reg_15_ ( .D(n510), .CLK(clk), .R(n750), .S(1'b1), .Q(
        evenBuffer[15]) );
  DFFSR evenBuffer_reg_14_ ( .D(n509), .CLK(clk), .R(n750), .S(1'b1), .Q(
        evenBuffer[14]) );
  DFFSR evenBuffer_reg_13_ ( .D(n508), .CLK(clk), .R(n750), .S(1'b1), .Q(
        evenBuffer[13]) );
  DFFSR evenBuffer_reg_12_ ( .D(n507), .CLK(clk), .R(n750), .S(1'b1), .Q(
        evenBuffer[12]) );
  DFFSR evenBuffer_reg_11_ ( .D(n506), .CLK(clk), .R(n749), .S(1'b1), .Q(
        evenBuffer[11]) );
  DFFSR evenBuffer_reg_10_ ( .D(n505), .CLK(clk), .R(n749), .S(1'b1), .Q(
        evenBuffer[10]) );
  DFFSR evenBuffer_reg_9_ ( .D(n504), .CLK(clk), .R(n749), .S(1'b1), .Q(
        evenBuffer[9]) );
  DFFSR evenBuffer_reg_8_ ( .D(n503), .CLK(clk), .R(n749), .S(1'b1), .Q(
        evenBuffer[8]) );
  DFFSR evenBuffer_reg_7_ ( .D(n502), .CLK(clk), .R(n749), .S(1'b1), .Q(
        evenBuffer[7]) );
  DFFSR evenBuffer_reg_6_ ( .D(n501), .CLK(clk), .R(n749), .S(1'b1), .Q(
        evenBuffer[6]) );
  DFFSR evenBuffer_reg_5_ ( .D(n500), .CLK(clk), .R(n749), .S(1'b1), .Q(
        evenBuffer[5]) );
  DFFSR evenBuffer_reg_4_ ( .D(n499), .CLK(clk), .R(n749), .S(1'b1), .Q(
        evenBuffer[4]) );
  DFFSR evenBuffer_reg_3_ ( .D(n498), .CLK(clk), .R(n749), .S(1'b1), .Q(
        evenBuffer[3]) );
  DFFSR evenBuffer_reg_2_ ( .D(n497), .CLK(clk), .R(n749), .S(1'b1), .Q(
        evenBuffer[2]) );
  DFFSR evenBuffer_reg_1_ ( .D(n496), .CLK(clk), .R(n749), .S(1'b1), .Q(
        evenBuffer[1]) );
  DFFSR evenBuffer_reg_0_ ( .D(n495), .CLK(clk), .R(n749), .S(1'b1), .Q(
        evenBuffer[0]) );
  NAND3X1 U278 ( .A(n742), .B(n764), .C(n644), .Y(n292) );
  NAND3X1 U279 ( .A(n657), .B(n674), .C(n756), .Y(n291) );
  NAND3X1 U281 ( .A(n864), .B(n765), .C(n742), .Y(n294) );
  NAND3X1 U282 ( .A(n674), .B(n800), .C(n756), .Y(n293) );
  NOR2X1 U283 ( .A(reset), .B(n227), .Y(readyIn) );
  AOI22X1 U284 ( .A(n756), .B(n798), .C(n797), .D(n766), .Y(n295) );
  OAI21X1 U285 ( .A(n296), .B(n918), .C(n679), .Y(n495) );
  OAI21X1 U287 ( .A(n296), .B(n917), .C(n678), .Y(n496) );
  OAI21X1 U289 ( .A(n296), .B(n916), .C(n635), .Y(n497) );
  OAI21X1 U291 ( .A(n296), .B(n915), .C(n623), .Y(n498) );
  OAI21X1 U293 ( .A(n296), .B(n914), .C(n287), .Y(n499) );
  OAI21X1 U295 ( .A(n296), .B(n913), .C(n278), .Y(n500) );
  OAI21X1 U297 ( .A(n296), .B(n912), .C(n269), .Y(n501) );
  OAI21X1 U299 ( .A(n296), .B(n911), .C(n260), .Y(n502) );
  OAI21X1 U301 ( .A(n296), .B(n910), .C(n253), .Y(n503) );
  OAI21X1 U303 ( .A(n296), .B(n909), .C(n246), .Y(n504) );
  OAI21X1 U305 ( .A(n296), .B(n908), .C(n239), .Y(n505) );
  OAI21X1 U307 ( .A(n296), .B(n907), .C(n233), .Y(n506) );
  OAI21X1 U309 ( .A(n296), .B(n906), .C(n677), .Y(n507) );
  OAI21X1 U311 ( .A(n296), .B(n905), .C(n634), .Y(n508) );
  OAI21X1 U313 ( .A(n296), .B(n904), .C(n622), .Y(n509) );
  OAI21X1 U315 ( .A(n296), .B(n903), .C(n286), .Y(n510) );
  OAI21X1 U317 ( .A(n296), .B(n902), .C(n268), .Y(n511) );
  OAI21X1 U319 ( .A(n296), .B(n901), .C(n226), .Y(n512) );
  OAI21X1 U321 ( .A(n296), .B(n900), .C(n225), .Y(n513) );
  OAI21X1 U323 ( .A(n296), .B(n899), .C(n224), .Y(n514) );
  OAI21X1 U325 ( .A(n296), .B(n898), .C(n223), .Y(n515) );
  OAI21X1 U327 ( .A(n296), .B(n897), .C(n222), .Y(n516) );
  OAI21X1 U329 ( .A(n296), .B(n896), .C(n221), .Y(n517) );
  OAI21X1 U331 ( .A(n296), .B(n895), .C(n277), .Y(n518) );
  OAI21X1 U333 ( .A(n296), .B(n894), .C(n259), .Y(n519) );
  OAI21X1 U335 ( .A(n296), .B(n893), .C(n633), .Y(n520) );
  OAI21X1 U337 ( .A(n296), .B(n892), .C(n621), .Y(n521) );
  OAI21X1 U339 ( .A(n296), .B(n891), .C(n285), .Y(n522) );
  OAI21X1 U341 ( .A(n296), .B(n890), .C(n267), .Y(n523) );
  OAI21X1 U343 ( .A(n296), .B(n889), .C(n252), .Y(n524) );
  OAI21X1 U345 ( .A(n296), .B(n888), .C(n245), .Y(n525) );
  OAI21X1 U347 ( .A(n296), .B(n887), .C(n238), .Y(n526) );
  OAI21X1 U349 ( .A(n296), .B(n886), .C(n232), .Y(n527) );
  OAI21X1 U351 ( .A(n296), .B(n885), .C(n220), .Y(n528) );
  OAI21X1 U353 ( .A(n296), .B(n884), .C(n219), .Y(n529) );
  OAI21X1 U355 ( .A(n296), .B(n883), .C(n218), .Y(n530) );
  OAI21X1 U357 ( .A(n296), .B(n882), .C(n217), .Y(n531) );
  OAI21X1 U359 ( .A(n296), .B(n881), .C(n216), .Y(n532) );
  OAI21X1 U361 ( .A(n296), .B(n880), .C(n215), .Y(n533) );
  OAI21X1 U363 ( .A(n296), .B(n879), .C(n676), .Y(n534) );
  OAI21X1 U365 ( .A(n296), .B(n878), .C(n632), .Y(n535) );
  OAI21X1 U367 ( .A(n296), .B(n877), .C(n620), .Y(n536) );
  OAI21X1 U369 ( .A(n296), .B(n876), .C(n284), .Y(n537) );
  OAI21X1 U371 ( .A(n296), .B(n875), .C(n276), .Y(n538) );
  OAI21X1 U373 ( .A(n296), .B(n874), .C(n266), .Y(n539) );
  OAI21X1 U375 ( .A(n296), .B(n873), .C(n258), .Y(n540) );
  OAI21X1 U377 ( .A(n296), .B(n872), .C(n251), .Y(n541) );
  OAI21X1 U379 ( .A(n296), .B(n871), .C(n244), .Y(n542) );
  AOI22X1 U381 ( .A(dataIn[48]), .B(n361), .C(n740), .D(n752), .Y(n345) );
  AOI22X1 U382 ( .A(dataIn[49]), .B(n361), .C(n739), .D(n752), .Y(n346) );
  AOI22X1 U383 ( .A(dataIn[50]), .B(n361), .C(n738), .D(n752), .Y(n347) );
  AOI22X1 U384 ( .A(dataIn[51]), .B(n361), .C(n737), .D(n752), .Y(n348) );
  AOI22X1 U385 ( .A(dataIn[52]), .B(n361), .C(n736), .D(n752), .Y(n349) );
  AOI22X1 U386 ( .A(dataIn[53]), .B(n361), .C(n735), .D(n752), .Y(n350) );
  AOI22X1 U387 ( .A(dataIn[54]), .B(n361), .C(n743), .D(n752), .Y(n351) );
  AOI22X1 U388 ( .A(dataIn[55]), .B(n361), .C(n741), .D(n752), .Y(n352) );
  OAI21X1 U389 ( .A(n296), .B(n870), .C(n237), .Y(n543) );
  OAI21X1 U391 ( .A(n296), .B(n869), .C(n231), .Y(n544) );
  OAI21X1 U393 ( .A(n296), .B(n868), .C(n214), .Y(n545) );
  OAI21X1 U395 ( .A(n296), .B(n867), .C(n213), .Y(n546) );
  OAI21X1 U397 ( .A(n296), .B(n866), .C(n212), .Y(n547) );
  OAI21X1 U399 ( .A(n296), .B(n865), .C(n211), .Y(n548) );
  OAI21X1 U401 ( .A(n864), .B(n296), .C(n210), .Y(n549) );
  OAI21X1 U403 ( .A(n296), .B(n863), .C(n275), .Y(n550) );
  OAI21X1 U405 ( .A(n747), .B(n862), .C(n664), .Y(n551) );
  OAI21X1 U407 ( .A(n747), .B(n861), .C(n651), .Y(n552) );
  OAI21X1 U409 ( .A(n747), .B(n860), .C(n641), .Y(n553) );
  OAI21X1 U411 ( .A(n747), .B(n859), .C(n630), .Y(n554) );
  OAI21X1 U413 ( .A(n747), .B(n858), .C(n619), .Y(n555) );
  OAI21X1 U415 ( .A(n747), .B(n857), .C(n283), .Y(n556) );
  OAI21X1 U417 ( .A(n747), .B(n856), .C(n274), .Y(n557) );
  OAI21X1 U419 ( .A(n747), .B(n855), .C(n265), .Y(n558) );
  OAI21X1 U421 ( .A(n747), .B(n854), .C(n663), .Y(n559) );
  OAI21X1 U423 ( .A(n747), .B(n853), .C(n257), .Y(n560) );
  OAI21X1 U425 ( .A(n747), .B(n852), .C(n250), .Y(n561) );
  OAI21X1 U427 ( .A(n747), .B(n851), .C(n243), .Y(n562) );
  OAI21X1 U429 ( .A(n747), .B(n850), .C(n650), .Y(n563) );
  OAI21X1 U431 ( .A(n747), .B(n849), .C(n640), .Y(n564) );
  OAI21X1 U433 ( .A(n747), .B(n848), .C(n629), .Y(n565) );
  OAI21X1 U435 ( .A(n747), .B(n847), .C(n618), .Y(n566) );
  OAI21X1 U437 ( .A(n747), .B(n846), .C(n282), .Y(n567) );
  OAI21X1 U439 ( .A(n747), .B(n845), .C(n273), .Y(n568) );
  OAI21X1 U441 ( .A(n747), .B(n844), .C(n264), .Y(n569) );
  OAI21X1 U443 ( .A(n747), .B(n843), .C(n236), .Y(n570) );
  OAI21X1 U445 ( .A(n747), .B(n842), .C(n662), .Y(n571) );
  OAI21X1 U447 ( .A(n747), .B(n841), .C(n256), .Y(n572) );
  OAI21X1 U449 ( .A(n747), .B(n840), .C(n249), .Y(n573) );
  OAI21X1 U451 ( .A(n747), .B(n839), .C(n242), .Y(n574) );
  OAI21X1 U453 ( .A(n747), .B(n838), .C(n209), .Y(n575) );
  OAI21X1 U455 ( .A(n747), .B(n837), .C(n649), .Y(n576) );
  OAI21X1 U457 ( .A(n747), .B(n836), .C(n639), .Y(n577) );
  OAI21X1 U459 ( .A(n747), .B(n835), .C(n628), .Y(n578) );
  OAI21X1 U461 ( .A(n747), .B(n834), .C(n617), .Y(n579) );
  OAI21X1 U463 ( .A(n747), .B(n833), .C(n281), .Y(n580) );
  OAI21X1 U465 ( .A(n747), .B(n832), .C(n272), .Y(n581) );
  OAI21X1 U467 ( .A(n747), .B(n831), .C(n263), .Y(n582) );
  OAI21X1 U469 ( .A(n747), .B(n830), .C(n255), .Y(n583) );
  OAI21X1 U471 ( .A(n747), .B(n829), .C(n248), .Y(n584) );
  OAI21X1 U473 ( .A(n747), .B(n828), .C(n241), .Y(n585) );
  OAI21X1 U475 ( .A(n747), .B(n827), .C(n235), .Y(n586) );
  OAI21X1 U477 ( .A(n747), .B(n826), .C(n208), .Y(n587) );
  OAI21X1 U479 ( .A(n747), .B(n825), .C(n661), .Y(n588) );
  OAI21X1 U481 ( .A(n747), .B(n824), .C(n648), .Y(n589) );
  OAI21X1 U483 ( .A(n747), .B(n823), .C(n638), .Y(n590) );
  OAI21X1 U485 ( .A(n747), .B(n822), .C(n627), .Y(n591) );
  OAI21X1 U487 ( .A(n747), .B(n821), .C(n290), .Y(n592) );
  OAI21X1 U489 ( .A(n747), .B(n820), .C(n280), .Y(n593) );
  OAI21X1 U491 ( .A(n747), .B(n819), .C(n271), .Y(n594) );
  OAI21X1 U493 ( .A(n747), .B(n818), .C(n262), .Y(n595) );
  OAI21X1 U495 ( .A(n747), .B(n817), .C(n254), .Y(n596) );
  OAI21X1 U497 ( .A(n747), .B(n816), .C(n247), .Y(n597) );
  OAI21X1 U499 ( .A(n747), .B(n815), .C(n240), .Y(n598) );
  OAI21X1 U501 ( .A(n926), .B(n410), .C(n647), .Y(n599) );
  OAI21X1 U503 ( .A(n925), .B(n410), .C(n637), .Y(n600) );
  OAI21X1 U505 ( .A(n924), .B(n410), .C(n626), .Y(n601) );
  OAI21X1 U507 ( .A(n923), .B(n410), .C(n289), .Y(n602) );
  OAI21X1 U509 ( .A(n922), .B(n410), .C(n279), .Y(n603) );
  OAI21X1 U511 ( .A(n921), .B(n410), .C(n660), .Y(n604) );
  OAI21X1 U513 ( .A(n920), .B(n410), .C(n270), .Y(n605) );
  OAI21X1 U515 ( .A(n919), .B(n410), .C(n261), .Y(n606) );
  OAI21X1 U517 ( .A(n747), .B(n806), .C(n234), .Y(n607) );
  OAI21X1 U519 ( .A(n747), .B(n805), .C(n207), .Y(n608) );
  OAI21X1 U521 ( .A(n747), .B(n804), .C(n659), .Y(n609) );
  OAI21X1 U523 ( .A(n747), .B(n803), .C(n646), .Y(n610) );
  OAI21X1 U525 ( .A(n747), .B(n802), .C(n636), .Y(n611) );
  OAI21X1 U527 ( .A(n747), .B(n801), .C(n625), .Y(n612) );
  OAI21X1 U529 ( .A(n800), .B(n747), .C(n206), .Y(n613) );
  OAI21X1 U531 ( .A(n747), .B(n799), .C(n288), .Y(n614) );
  OAI21X1 U533 ( .A(n798), .B(n296), .C(n667), .Y(n615) );
  OAI21X1 U535 ( .A(n756), .B(n228), .C(n652), .Y(n296) );
  OAI21X1 U537 ( .A(n797), .B(n747), .C(n410), .Y(n616) );
  AOI21X1 U539 ( .A(n766), .B(sendIn), .C(n745), .Y(n412) );
  OAI21X1 U542 ( .A(n756), .B(n909), .C(n205), .Y(dataOut[9]) );
  OAI21X1 U544 ( .A(n758), .B(n910), .C(n204), .Y(dataOut[8]) );
  OAI21X1 U546 ( .A(n757), .B(n911), .C(n203), .Y(dataOut[7]) );
  OAI21X1 U548 ( .A(n757), .B(n912), .C(n202), .Y(dataOut[6]) );
  OAI21X1 U550 ( .A(n757), .B(n863), .C(n201), .Y(dataOut[63]) );
  OAI21X1 U552 ( .A(n758), .B(n864), .C(n624), .Y(dataOut[62]) );
  OAI21X1 U554 ( .A(n757), .B(n865), .C(n200), .Y(dataOut[61]) );
  OAI21X1 U556 ( .A(n757), .B(n866), .C(n199), .Y(dataOut[60]) );
  OAI21X1 U558 ( .A(n757), .B(n913), .C(n198), .Y(dataOut[5]) );
  OAI21X1 U560 ( .A(n758), .B(n867), .C(n197), .Y(dataOut[59]) );
  OAI21X1 U562 ( .A(n757), .B(n868), .C(n196), .Y(dataOut[58]) );
  OAI21X1 U564 ( .A(n757), .B(n869), .C(n195), .Y(dataOut[57]) );
  OAI21X1 U566 ( .A(n758), .B(n870), .C(n194), .Y(dataOut[56]) );
  AOI22X1 U568 ( .A(n146), .B(n766), .C(n157), .D(n756), .Y(n444) );
  AOI22X1 U569 ( .A(n145), .B(n766), .C(n156), .D(n756), .Y(n445) );
  AOI22X1 U570 ( .A(n144), .B(n766), .C(n155), .D(n756), .Y(n446) );
  AOI22X1 U571 ( .A(n143), .B(n766), .C(n154), .D(n756), .Y(n447) );
  AOI22X1 U572 ( .A(n142), .B(n766), .C(n153), .D(n756), .Y(n448) );
  AOI22X1 U573 ( .A(n141), .B(n766), .C(n152), .D(n756), .Y(n449) );
  OAI21X1 U574 ( .A(n758), .B(n914), .C(n193), .Y(dataOut[4]) );
  AOI22X1 U576 ( .A(n140), .B(n766), .C(n151), .D(n756), .Y(n451) );
  AOI22X1 U577 ( .A(n139), .B(n766), .C(n150), .D(n756), .Y(n452) );
  OAI21X1 U578 ( .A(n758), .B(n871), .C(n192), .Y(dataOut[47]) );
  OAI21X1 U580 ( .A(n758), .B(n872), .C(n191), .Y(dataOut[46]) );
  OAI21X1 U582 ( .A(n758), .B(n873), .C(n190), .Y(dataOut[45]) );
  OAI21X1 U584 ( .A(n759), .B(n874), .C(n189), .Y(dataOut[44]) );
  OAI21X1 U586 ( .A(n759), .B(n875), .C(n188), .Y(dataOut[43]) );
  OAI21X1 U588 ( .A(n758), .B(n876), .C(n187), .Y(dataOut[42]) );
  OAI21X1 U590 ( .A(n759), .B(n877), .C(n186), .Y(dataOut[41]) );
  OAI21X1 U592 ( .A(n759), .B(n878), .C(n185), .Y(dataOut[40]) );
  OAI21X1 U594 ( .A(n758), .B(n915), .C(n184), .Y(dataOut[3]) );
  OAI21X1 U596 ( .A(n759), .B(n879), .C(n183), .Y(dataOut[39]) );
  OAI21X1 U598 ( .A(n760), .B(n880), .C(n182), .Y(dataOut[38]) );
  OAI21X1 U600 ( .A(n759), .B(n881), .C(n181), .Y(dataOut[37]) );
  OAI21X1 U602 ( .A(n760), .B(n882), .C(n180), .Y(dataOut[36]) );
  OAI21X1 U604 ( .A(n760), .B(n883), .C(n179), .Y(dataOut[35]) );
  OAI21X1 U606 ( .A(n759), .B(n884), .C(n178), .Y(dataOut[34]) );
  OAI21X1 U608 ( .A(n760), .B(n885), .C(n177), .Y(dataOut[33]) );
  OAI21X1 U610 ( .A(n760), .B(n886), .C(n176), .Y(dataOut[32]) );
  OAI21X1 U612 ( .A(n759), .B(n887), .C(n175), .Y(dataOut[31]) );
  OAI21X1 U614 ( .A(n760), .B(n888), .C(n174), .Y(dataOut[30]) );
  OAI21X1 U616 ( .A(n760), .B(n916), .C(n173), .Y(dataOut[2]) );
  OAI21X1 U618 ( .A(n760), .B(n889), .C(n172), .Y(dataOut[29]) );
  OAI21X1 U620 ( .A(n761), .B(n890), .C(n171), .Y(dataOut[28]) );
  OAI21X1 U622 ( .A(n761), .B(n891), .C(n170), .Y(dataOut[27]) );
  OAI21X1 U624 ( .A(n760), .B(n892), .C(n169), .Y(dataOut[26]) );
  OAI21X1 U626 ( .A(n760), .B(n893), .C(n168), .Y(dataOut[25]) );
  OAI21X1 U628 ( .A(n761), .B(n894), .C(n167), .Y(dataOut[24]) );
  OAI21X1 U630 ( .A(n760), .B(n895), .C(n166), .Y(dataOut[23]) );
  OAI21X1 U632 ( .A(n759), .B(n896), .C(n165), .Y(dataOut[22]) );
  OAI21X1 U634 ( .A(n760), .B(n897), .C(n164), .Y(dataOut[21]) );
  OAI21X1 U636 ( .A(n760), .B(n898), .C(n163), .Y(dataOut[20]) );
  OAI21X1 U638 ( .A(n759), .B(n917), .C(n162), .Y(dataOut[1]) );
  OAI21X1 U640 ( .A(n759), .B(n899), .C(n161), .Y(dataOut[19]) );
  OAI21X1 U642 ( .A(n759), .B(n900), .C(n160), .Y(dataOut[18]) );
  OAI21X1 U644 ( .A(n758), .B(n901), .C(n159), .Y(dataOut[17]) );
  OAI21X1 U646 ( .A(n759), .B(n902), .C(n158), .Y(dataOut[16]) );
  OAI21X1 U648 ( .A(n758), .B(n903), .C(n149), .Y(dataOut[15]) );
  OAI21X1 U650 ( .A(n758), .B(n904), .C(n148), .Y(dataOut[14]) );
  OAI21X1 U652 ( .A(n757), .B(n905), .C(n147), .Y(dataOut[13]) );
  OAI21X1 U654 ( .A(n757), .B(n906), .C(n138), .Y(dataOut[12]) );
  OAI21X1 U656 ( .A(n757), .B(n907), .C(n137), .Y(dataOut[11]) );
  OAI21X1 U658 ( .A(n757), .B(n908), .C(n136), .Y(dataOut[10]) );
  OAI21X1 U660 ( .A(n757), .B(n918), .C(n135), .Y(dataOut[0]) );
  OR2X1 U132 ( .A(n766), .B(n228), .Y(n430) );
  AND2X1 U134 ( .A(n132), .B(n134), .Y(n927) );
  OR2X1 U135 ( .A(n658), .B(n743), .Y(n772) );
  OR2X1 U136 ( .A(n675), .B(n645), .Y(n783) );
  AND2X1 U137 ( .A(n130), .B(n133), .Y(n928) );
  AND2X1 U138 ( .A(n653), .B(n744), .Y(n417) );
  BUFX2 U139 ( .A(n293), .Y(n130) );
  BUFX2 U140 ( .A(n291), .Y(n132) );
  BUFX2 U141 ( .A(n294), .Y(n133) );
  BUFX2 U142 ( .A(n292), .Y(n134) );
  AND2X1 U143 ( .A(n734), .B(n762), .Y(n494) );
  INVX1 U144 ( .A(n494), .Y(n135) );
  AND2X1 U145 ( .A(n724), .B(n761), .Y(n493) );
  INVX1 U146 ( .A(n493), .Y(n136) );
  AND2X1 U147 ( .A(n723), .B(n761), .Y(n492) );
  INVX1 U148 ( .A(n492), .Y(n137) );
  AND2X1 U149 ( .A(n722), .B(n761), .Y(n491) );
  INVX1 U150 ( .A(n491), .Y(n138) );
  AND2X1 U151 ( .A(n721), .B(n761), .Y(n490) );
  INVX1 U152 ( .A(n490), .Y(n147) );
  AND2X1 U153 ( .A(n720), .B(n761), .Y(n489) );
  INVX1 U154 ( .A(n489), .Y(n148) );
  AND2X1 U155 ( .A(n719), .B(n762), .Y(n488) );
  INVX1 U156 ( .A(n488), .Y(n149) );
  AND2X1 U157 ( .A(n718), .B(n762), .Y(n487) );
  INVX1 U158 ( .A(n487), .Y(n158) );
  AND2X1 U159 ( .A(n717), .B(n761), .Y(n486) );
  INVX1 U160 ( .A(n486), .Y(n159) );
  AND2X1 U161 ( .A(n716), .B(n761), .Y(n485) );
  INVX1 U162 ( .A(n485), .Y(n160) );
  AND2X1 U163 ( .A(n715), .B(n762), .Y(n484) );
  INVX1 U164 ( .A(n484), .Y(n161) );
  AND2X1 U165 ( .A(n733), .B(n761), .Y(n483) );
  INVX1 U166 ( .A(n483), .Y(n162) );
  AND2X1 U167 ( .A(n714), .B(n761), .Y(n482) );
  INVX1 U168 ( .A(n482), .Y(n163) );
  AND2X1 U169 ( .A(n713), .B(n762), .Y(n481) );
  INVX1 U170 ( .A(n481), .Y(n164) );
  AND2X1 U171 ( .A(n712), .B(n761), .Y(n480) );
  INVX1 U172 ( .A(n480), .Y(n165) );
  AND2X1 U173 ( .A(n711), .B(n761), .Y(n479) );
  INVX1 U174 ( .A(n479), .Y(n166) );
  AND2X1 U175 ( .A(n710), .B(n762), .Y(n478) );
  INVX1 U176 ( .A(n478), .Y(n167) );
  AND2X1 U177 ( .A(n709), .B(n762), .Y(n477) );
  INVX1 U178 ( .A(n477), .Y(n168) );
  AND2X1 U179 ( .A(n708), .B(n762), .Y(n476) );
  INVX1 U180 ( .A(n476), .Y(n169) );
  AND2X1 U181 ( .A(n707), .B(n762), .Y(n475) );
  INVX1 U182 ( .A(n475), .Y(n170) );
  AND2X1 U183 ( .A(n706), .B(n762), .Y(n474) );
  INVX1 U184 ( .A(n474), .Y(n171) );
  AND2X1 U185 ( .A(n705), .B(n762), .Y(n473) );
  INVX1 U186 ( .A(n473), .Y(n172) );
  AND2X1 U187 ( .A(n732), .B(n762), .Y(n472) );
  INVX1 U188 ( .A(n472), .Y(n173) );
  AND2X1 U189 ( .A(n704), .B(n762), .Y(n471) );
  INVX1 U190 ( .A(n471), .Y(n174) );
  AND2X1 U191 ( .A(n703), .B(n762), .Y(n470) );
  INVX1 U192 ( .A(n470), .Y(n175) );
  AND2X1 U193 ( .A(n702), .B(n762), .Y(n469) );
  INVX1 U194 ( .A(n469), .Y(n176) );
  AND2X1 U195 ( .A(n701), .B(n762), .Y(n468) );
  INVX1 U196 ( .A(n468), .Y(n177) );
  AND2X1 U197 ( .A(n700), .B(n762), .Y(n467) );
  INVX1 U198 ( .A(n467), .Y(n178) );
  AND2X1 U199 ( .A(n699), .B(n762), .Y(n466) );
  INVX1 U200 ( .A(n466), .Y(n179) );
  AND2X1 U201 ( .A(n698), .B(n763), .Y(n465) );
  INVX1 U202 ( .A(n465), .Y(n180) );
  AND2X1 U203 ( .A(n697), .B(n763), .Y(n464) );
  INVX1 U204 ( .A(n464), .Y(n181) );
  AND2X1 U205 ( .A(n696), .B(n763), .Y(n463) );
  INVX1 U206 ( .A(n463), .Y(n182) );
  AND2X1 U207 ( .A(n695), .B(n763), .Y(n462) );
  INVX1 U208 ( .A(n462), .Y(n183) );
  AND2X1 U209 ( .A(n731), .B(n763), .Y(n461) );
  INVX1 U210 ( .A(n461), .Y(n184) );
  AND2X1 U211 ( .A(n694), .B(n763), .Y(n460) );
  INVX1 U212 ( .A(n460), .Y(n185) );
  AND2X1 U213 ( .A(n693), .B(n763), .Y(n459) );
  INVX1 U214 ( .A(n459), .Y(n186) );
  AND2X1 U215 ( .A(n692), .B(n763), .Y(n458) );
  INVX1 U216 ( .A(n458), .Y(n187) );
  AND2X1 U217 ( .A(n691), .B(n763), .Y(n457) );
  INVX1 U218 ( .A(n457), .Y(n188) );
  AND2X1 U219 ( .A(n690), .B(n763), .Y(n456) );
  INVX1 U220 ( .A(n456), .Y(n189) );
  AND2X1 U221 ( .A(n689), .B(n763), .Y(n455) );
  INVX1 U222 ( .A(n455), .Y(n190) );
  AND2X1 U223 ( .A(n688), .B(n763), .Y(n454) );
  INVX1 U224 ( .A(n454), .Y(n191) );
  AND2X1 U225 ( .A(n687), .B(n763), .Y(n453) );
  INVX1 U226 ( .A(n453), .Y(n192) );
  AND2X1 U227 ( .A(n730), .B(n763), .Y(n450) );
  INVX1 U228 ( .A(n450), .Y(n193) );
  AND2X1 U229 ( .A(n686), .B(n763), .Y(n443) );
  INVX1 U230 ( .A(n443), .Y(n194) );
  AND2X1 U231 ( .A(n685), .B(n763), .Y(n442) );
  INVX1 U232 ( .A(n442), .Y(n195) );
  AND2X1 U233 ( .A(n684), .B(n763), .Y(n441) );
  INVX1 U234 ( .A(n441), .Y(n196) );
  AND2X1 U235 ( .A(n683), .B(n763), .Y(n440) );
  INVX1 U236 ( .A(n440), .Y(n197) );
  AND2X1 U237 ( .A(n729), .B(n758), .Y(n439) );
  INVX1 U238 ( .A(n439), .Y(n198) );
  AND2X1 U239 ( .A(n682), .B(n760), .Y(n438) );
  INVX1 U240 ( .A(n438), .Y(n199) );
  AND2X1 U241 ( .A(n681), .B(n759), .Y(n437) );
  INVX1 U242 ( .A(n437), .Y(n200) );
  AND2X1 U243 ( .A(n680), .B(n757), .Y(n435) );
  INVX1 U244 ( .A(n435), .Y(n201) );
  AND2X1 U245 ( .A(n728), .B(n758), .Y(n434) );
  INVX1 U246 ( .A(n434), .Y(n202) );
  AND2X1 U247 ( .A(n727), .B(n757), .Y(n433) );
  INVX1 U248 ( .A(n433), .Y(n203) );
  AND2X1 U249 ( .A(n726), .B(n760), .Y(n432) );
  INVX1 U250 ( .A(n432), .Y(n204) );
  AND2X1 U251 ( .A(n725), .B(n759), .Y(n431) );
  INVX1 U252 ( .A(n431), .Y(n205) );
  AND2X1 U253 ( .A(n746), .B(dataIn[62]), .Y(n426) );
  INVX1 U254 ( .A(n426), .Y(n206) );
  AND2X1 U255 ( .A(n746), .B(dataIn[57]), .Y(n421) );
  INVX1 U256 ( .A(n421), .Y(n207) );
  AND2X1 U257 ( .A(n746), .B(dataIn[36]), .Y(n398) );
  INVX1 U258 ( .A(n398), .Y(n208) );
  AND2X1 U259 ( .A(n746), .B(dataIn[24]), .Y(n386) );
  INVX1 U260 ( .A(n386), .Y(n209) );
  AND2X1 U261 ( .A(dataIn[62]), .B(n361), .Y(n359) );
  INVX1 U262 ( .A(n359), .Y(n210) );
  AND2X1 U263 ( .A(dataIn[61]), .B(n361), .Y(n358) );
  INVX1 U264 ( .A(n358), .Y(n211) );
  AND2X1 U265 ( .A(dataIn[60]), .B(n361), .Y(n357) );
  INVX1 U266 ( .A(n357), .Y(n212) );
  AND2X1 U267 ( .A(dataIn[59]), .B(n361), .Y(n356) );
  INVX1 U268 ( .A(n356), .Y(n213) );
  AND2X1 U269 ( .A(dataIn[58]), .B(n361), .Y(n355) );
  INVX1 U270 ( .A(n355), .Y(n214) );
  AND2X1 U271 ( .A(dataIn[38]), .B(n361), .Y(n335) );
  INVX1 U272 ( .A(n335), .Y(n215) );
  AND2X1 U273 ( .A(dataIn[37]), .B(n361), .Y(n334) );
  INVX1 U274 ( .A(n334), .Y(n216) );
  AND2X1 U275 ( .A(dataIn[36]), .B(n361), .Y(n333) );
  INVX1 U276 ( .A(n333), .Y(n217) );
  AND2X1 U277 ( .A(dataIn[35]), .B(n361), .Y(n332) );
  INVX1 U280 ( .A(n332), .Y(n218) );
  AND2X1 U286 ( .A(dataIn[34]), .B(n361), .Y(n331) );
  INVX1 U288 ( .A(n331), .Y(n219) );
  AND2X1 U290 ( .A(dataIn[33]), .B(n361), .Y(n330) );
  INVX1 U292 ( .A(n330), .Y(n220) );
  AND2X1 U294 ( .A(dataIn[22]), .B(n748), .Y(n319) );
  INVX1 U296 ( .A(n319), .Y(n221) );
  AND2X1 U298 ( .A(dataIn[21]), .B(n748), .Y(n318) );
  INVX1 U300 ( .A(n318), .Y(n222) );
  AND2X1 U302 ( .A(dataIn[20]), .B(n748), .Y(n317) );
  INVX1 U304 ( .A(n317), .Y(n223) );
  AND2X1 U306 ( .A(dataIn[19]), .B(n748), .Y(n316) );
  INVX1 U308 ( .A(n316), .Y(n224) );
  AND2X1 U310 ( .A(dataIn[18]), .B(n748), .Y(n315) );
  INVX1 U312 ( .A(n315), .Y(n225) );
  AND2X1 U314 ( .A(dataIn[17]), .B(n748), .Y(n314) );
  INVX1 U316 ( .A(n314), .Y(n226) );
  BUFX2 U318 ( .A(n295), .Y(n227) );
  OR2X1 U320 ( .A(outputBufferGrant[0]), .B(outputBufferGrant[1]), .Y(n428) );
  INVX1 U322 ( .A(n428), .Y(n228) );
  INVX1 U324 ( .A(n928), .Y(request[0]) );
  INVX1 U326 ( .A(n927), .Y(request[1]) );
  AND2X1 U328 ( .A(dataIn[57]), .B(n361), .Y(n354) );
  INVX1 U330 ( .A(n354), .Y(n231) );
  AND2X1 U332 ( .A(dataIn[32]), .B(n361), .Y(n329) );
  INVX1 U334 ( .A(n329), .Y(n232) );
  AND2X1 U336 ( .A(dataIn[11]), .B(n748), .Y(n308) );
  INVX1 U338 ( .A(n308), .Y(n233) );
  AND2X1 U340 ( .A(n746), .B(dataIn[56]), .Y(n420) );
  INVX1 U342 ( .A(n420), .Y(n234) );
  AND2X1 U344 ( .A(n746), .B(dataIn[35]), .Y(n397) );
  INVX1 U346 ( .A(n397), .Y(n235) );
  AND2X1 U348 ( .A(n746), .B(dataIn[19]), .Y(n381) );
  INVX1 U350 ( .A(n381), .Y(n236) );
  AND2X1 U352 ( .A(dataIn[56]), .B(n361), .Y(n353) );
  INVX1 U354 ( .A(n353), .Y(n237) );
  AND2X1 U356 ( .A(dataIn[31]), .B(n361), .Y(n328) );
  INVX1 U358 ( .A(n328), .Y(n238) );
  AND2X1 U360 ( .A(dataIn[10]), .B(n748), .Y(n307) );
  INVX1 U362 ( .A(n307), .Y(n239) );
  AND2X1 U364 ( .A(n746), .B(dataIn[47]), .Y(n409) );
  INVX1 U366 ( .A(n409), .Y(n240) );
  AND2X1 U368 ( .A(n746), .B(dataIn[34]), .Y(n396) );
  INVX1 U370 ( .A(n396), .Y(n241) );
  AND2X1 U372 ( .A(n746), .B(dataIn[23]), .Y(n385) );
  INVX1 U374 ( .A(n385), .Y(n242) );
  AND2X1 U376 ( .A(n746), .B(dataIn[11]), .Y(n373) );
  INVX1 U378 ( .A(n373), .Y(n243) );
  AND2X1 U380 ( .A(dataIn[47]), .B(n361), .Y(n344) );
  INVX1 U390 ( .A(n344), .Y(n244) );
  AND2X1 U392 ( .A(dataIn[30]), .B(n361), .Y(n327) );
  INVX1 U394 ( .A(n327), .Y(n245) );
  AND2X1 U396 ( .A(dataIn[9]), .B(n748), .Y(n306) );
  INVX1 U398 ( .A(n306), .Y(n246) );
  AND2X1 U400 ( .A(n746), .B(dataIn[46]), .Y(n408) );
  INVX1 U402 ( .A(n408), .Y(n247) );
  AND2X1 U404 ( .A(n746), .B(dataIn[33]), .Y(n395) );
  INVX1 U406 ( .A(n395), .Y(n248) );
  AND2X1 U408 ( .A(n746), .B(dataIn[22]), .Y(n384) );
  INVX1 U410 ( .A(n384), .Y(n249) );
  AND2X1 U412 ( .A(n746), .B(dataIn[10]), .Y(n372) );
  INVX1 U414 ( .A(n372), .Y(n250) );
  AND2X1 U416 ( .A(dataIn[46]), .B(n361), .Y(n343) );
  INVX1 U418 ( .A(n343), .Y(n251) );
  AND2X1 U420 ( .A(dataIn[29]), .B(n361), .Y(n326) );
  INVX1 U422 ( .A(n326), .Y(n252) );
  AND2X1 U424 ( .A(dataIn[8]), .B(n748), .Y(n305) );
  INVX1 U426 ( .A(n305), .Y(n253) );
  AND2X1 U428 ( .A(n746), .B(dataIn[45]), .Y(n407) );
  INVX1 U430 ( .A(n407), .Y(n254) );
  AND2X1 U432 ( .A(n746), .B(dataIn[32]), .Y(n394) );
  INVX1 U434 ( .A(n394), .Y(n255) );
  AND2X1 U436 ( .A(n746), .B(dataIn[21]), .Y(n383) );
  INVX1 U438 ( .A(n383), .Y(n256) );
  AND2X1 U440 ( .A(n746), .B(dataIn[9]), .Y(n371) );
  INVX1 U442 ( .A(n371), .Y(n257) );
  AND2X1 U444 ( .A(dataIn[45]), .B(n361), .Y(n342) );
  INVX1 U446 ( .A(n342), .Y(n258) );
  AND2X1 U448 ( .A(dataIn[24]), .B(n361), .Y(n321) );
  INVX1 U450 ( .A(n321), .Y(n259) );
  AND2X1 U452 ( .A(dataIn[7]), .B(n748), .Y(n304) );
  INVX1 U454 ( .A(n304), .Y(n260) );
  AND2X1 U456 ( .A(n673), .B(n744), .Y(n419) );
  INVX1 U458 ( .A(n419), .Y(n261) );
  AND2X1 U460 ( .A(n746), .B(dataIn[44]), .Y(n406) );
  INVX1 U462 ( .A(n406), .Y(n262) );
  AND2X1 U464 ( .A(n746), .B(dataIn[31]), .Y(n393) );
  INVX1 U466 ( .A(n393), .Y(n263) );
  AND2X1 U468 ( .A(n746), .B(dataIn[18]), .Y(n380) );
  INVX1 U470 ( .A(n380), .Y(n264) );
  AND2X1 U472 ( .A(n746), .B(dataIn[7]), .Y(n369) );
  INVX1 U474 ( .A(n369), .Y(n265) );
  AND2X1 U476 ( .A(dataIn[44]), .B(n361), .Y(n341) );
  INVX1 U478 ( .A(n341), .Y(n266) );
  AND2X1 U480 ( .A(dataIn[28]), .B(n361), .Y(n325) );
  INVX1 U482 ( .A(n325), .Y(n267) );
  AND2X1 U484 ( .A(dataIn[16]), .B(n748), .Y(n313) );
  INVX1 U486 ( .A(n313), .Y(n268) );
  AND2X1 U488 ( .A(dataIn[6]), .B(n361), .Y(n303) );
  INVX1 U490 ( .A(n303), .Y(n269) );
  AND2X1 U492 ( .A(n645), .B(n744), .Y(n418) );
  INVX1 U494 ( .A(n418), .Y(n270) );
  AND2X1 U496 ( .A(n746), .B(dataIn[43]), .Y(n405) );
  INVX1 U498 ( .A(n405), .Y(n271) );
  AND2X1 U500 ( .A(n746), .B(dataIn[30]), .Y(n392) );
  INVX1 U502 ( .A(n392), .Y(n272) );
  AND2X1 U504 ( .A(n746), .B(dataIn[17]), .Y(n379) );
  INVX1 U506 ( .A(n379), .Y(n273) );
  AND2X1 U508 ( .A(n746), .B(dataIn[6]), .Y(n368) );
  INVX1 U510 ( .A(n368), .Y(n274) );
  AND2X1 U512 ( .A(dataIn[63]), .B(n361), .Y(n360) );
  INVX1 U514 ( .A(n360), .Y(n275) );
  AND2X1 U516 ( .A(dataIn[43]), .B(n361), .Y(n340) );
  INVX1 U518 ( .A(n340), .Y(n276) );
  AND2X1 U520 ( .A(dataIn[23]), .B(n361), .Y(n320) );
  INVX1 U522 ( .A(n320), .Y(n277) );
  AND2X1 U524 ( .A(dataIn[5]), .B(n748), .Y(n302) );
  INVX1 U526 ( .A(n302), .Y(n278) );
  AND2X1 U528 ( .A(n668), .B(n744), .Y(n416) );
  INVX1 U530 ( .A(n416), .Y(n279) );
  AND2X1 U532 ( .A(n746), .B(dataIn[42]), .Y(n404) );
  INVX1 U534 ( .A(n404), .Y(n280) );
  AND2X1 U536 ( .A(n746), .B(dataIn[29]), .Y(n391) );
  INVX1 U538 ( .A(n391), .Y(n281) );
  AND2X1 U540 ( .A(n746), .B(dataIn[16]), .Y(n378) );
  INVX1 U541 ( .A(n378), .Y(n282) );
  AND2X1 U543 ( .A(n746), .B(dataIn[5]), .Y(n367) );
  INVX1 U545 ( .A(n367), .Y(n283) );
  AND2X1 U547 ( .A(dataIn[42]), .B(n361), .Y(n339) );
  INVX1 U549 ( .A(n339), .Y(n284) );
  AND2X1 U551 ( .A(dataIn[27]), .B(n361), .Y(n324) );
  INVX1 U553 ( .A(n324), .Y(n285) );
  AND2X1 U555 ( .A(dataIn[15]), .B(n748), .Y(n312) );
  INVX1 U557 ( .A(n312), .Y(n286) );
  AND2X1 U559 ( .A(dataIn[4]), .B(n361), .Y(n301) );
  INVX1 U561 ( .A(n301), .Y(n287) );
  AND2X1 U563 ( .A(n746), .B(dataIn[63]), .Y(n427) );
  INVX1 U565 ( .A(n427), .Y(n288) );
  AND2X1 U567 ( .A(n669), .B(n744), .Y(n415) );
  INVX1 U575 ( .A(n415), .Y(n289) );
  AND2X1 U579 ( .A(n746), .B(dataIn[41]), .Y(n403) );
  INVX1 U581 ( .A(n403), .Y(n290) );
  AND2X1 U583 ( .A(n746), .B(dataIn[28]), .Y(n390) );
  INVX1 U585 ( .A(n390), .Y(n617) );
  AND2X1 U587 ( .A(n746), .B(dataIn[15]), .Y(n377) );
  INVX1 U589 ( .A(n377), .Y(n618) );
  AND2X1 U591 ( .A(n746), .B(dataIn[4]), .Y(n366) );
  INVX1 U593 ( .A(n366), .Y(n619) );
  AND2X1 U595 ( .A(dataIn[41]), .B(n361), .Y(n338) );
  INVX1 U597 ( .A(n338), .Y(n620) );
  AND2X1 U599 ( .A(dataIn[26]), .B(n361), .Y(n323) );
  INVX1 U601 ( .A(n323), .Y(n621) );
  AND2X1 U603 ( .A(dataIn[14]), .B(n748), .Y(n311) );
  INVX1 U605 ( .A(n311), .Y(n622) );
  AND2X1 U607 ( .A(dataIn[3]), .B(n361), .Y(n300) );
  INVX1 U609 ( .A(n300), .Y(n623) );
  AND2X1 U611 ( .A(n761), .B(n657), .Y(n436) );
  INVX1 U613 ( .A(n436), .Y(n624) );
  AND2X1 U615 ( .A(n746), .B(dataIn[61]), .Y(n425) );
  INVX1 U617 ( .A(n425), .Y(n625) );
  AND2X1 U619 ( .A(n670), .B(n744), .Y(n414) );
  INVX1 U621 ( .A(n414), .Y(n626) );
  AND2X1 U623 ( .A(n746), .B(dataIn[40]), .Y(n402) );
  INVX1 U625 ( .A(n402), .Y(n627) );
  AND2X1 U627 ( .A(n746), .B(dataIn[27]), .Y(n389) );
  INVX1 U629 ( .A(n389), .Y(n628) );
  AND2X1 U631 ( .A(n746), .B(dataIn[14]), .Y(n376) );
  INVX1 U633 ( .A(n376), .Y(n629) );
  AND2X1 U635 ( .A(n746), .B(dataIn[3]), .Y(n365) );
  INVX1 U637 ( .A(n365), .Y(n630) );
  AND2X1 U639 ( .A(n780), .B(n787), .Y(n781) );
  INVX1 U641 ( .A(n781), .Y(n631) );
  AND2X1 U643 ( .A(dataIn[40]), .B(n361), .Y(n337) );
  INVX1 U645 ( .A(n337), .Y(n632) );
  AND2X1 U647 ( .A(dataIn[25]), .B(n361), .Y(n322) );
  INVX1 U649 ( .A(n322), .Y(n633) );
  AND2X1 U651 ( .A(dataIn[13]), .B(n748), .Y(n310) );
  INVX1 U653 ( .A(n310), .Y(n634) );
  AND2X1 U655 ( .A(dataIn[2]), .B(n361), .Y(n299) );
  INVX1 U657 ( .A(n299), .Y(n635) );
  AND2X1 U659 ( .A(n746), .B(dataIn[60]), .Y(n424) );
  INVX1 U661 ( .A(n424), .Y(n636) );
  AND2X1 U662 ( .A(n671), .B(n744), .Y(n413) );
  INVX1 U663 ( .A(n413), .Y(n637) );
  AND2X1 U664 ( .A(n746), .B(dataIn[39]), .Y(n401) );
  INVX1 U665 ( .A(n401), .Y(n638) );
  AND2X1 U666 ( .A(n746), .B(dataIn[26]), .Y(n388) );
  INVX1 U667 ( .A(n388), .Y(n639) );
  AND2X1 U668 ( .A(n746), .B(dataIn[13]), .Y(n375) );
  INVX1 U669 ( .A(n375), .Y(n640) );
  AND2X1 U670 ( .A(n746), .B(dataIn[2]), .Y(n364) );
  INVX1 U671 ( .A(n364), .Y(n641) );
  AND2X1 U672 ( .A(n769), .B(n776), .Y(n770) );
  INVX1 U673 ( .A(n770), .Y(n642) );
  AND2X1 U674 ( .A(n778), .B(n785), .Y(n779) );
  INVX1 U675 ( .A(n779), .Y(n643) );
  BUFX2 U676 ( .A(evenBuffer[62]), .Y(n644) );
  BUFX2 U677 ( .A(oddBuffer[54]), .Y(n645) );
  AND2X1 U678 ( .A(n746), .B(dataIn[59]), .Y(n423) );
  INVX1 U679 ( .A(n423), .Y(n646) );
  AND2X1 U680 ( .A(n672), .B(n744), .Y(n411) );
  INVX1 U681 ( .A(n411), .Y(n647) );
  AND2X1 U682 ( .A(n746), .B(dataIn[38]), .Y(n400) );
  INVX1 U683 ( .A(n400), .Y(n648) );
  AND2X1 U684 ( .A(n746), .B(dataIn[25]), .Y(n387) );
  INVX1 U685 ( .A(n387), .Y(n649) );
  AND2X1 U686 ( .A(n746), .B(dataIn[12]), .Y(n374) );
  INVX1 U687 ( .A(n374), .Y(n650) );
  AND2X1 U688 ( .A(n746), .B(dataIn[1]), .Y(n363) );
  INVX1 U689 ( .A(n363), .Y(n651) );
  AND2X1 U690 ( .A(sendIn), .B(n761), .Y(n429) );
  INVX1 U691 ( .A(n429), .Y(n652) );
  BUFX2 U692 ( .A(oddBuffer[53]), .Y(n653) );
  AND2X1 U693 ( .A(n779), .B(n786), .Y(n780) );
  INVX1 U694 ( .A(n780), .Y(n654) );
  AND2X1 U695 ( .A(n767), .B(n774), .Y(n768) );
  INVX1 U696 ( .A(n768), .Y(n655) );
  AND2X1 U697 ( .A(n784), .B(n150), .Y(n778) );
  INVX1 U698 ( .A(n778), .Y(n656) );
  BUFX2 U699 ( .A(oddBuffer[62]), .Y(n657) );
  AND2X1 U700 ( .A(n770), .B(n777), .Y(n771) );
  INVX1 U701 ( .A(n771), .Y(n658) );
  AND2X1 U702 ( .A(n746), .B(dataIn[58]), .Y(n422) );
  INVX1 U703 ( .A(n422), .Y(n659) );
  INVX1 U704 ( .A(n417), .Y(n660) );
  AND2X1 U705 ( .A(n746), .B(dataIn[37]), .Y(n399) );
  INVX1 U706 ( .A(n399), .Y(n661) );
  AND2X1 U707 ( .A(n746), .B(dataIn[20]), .Y(n382) );
  INVX1 U708 ( .A(n382), .Y(n662) );
  AND2X1 U709 ( .A(n746), .B(dataIn[8]), .Y(n370) );
  INVX1 U710 ( .A(n370), .Y(n663) );
  AND2X1 U711 ( .A(n746), .B(dataIn[0]), .Y(n362) );
  INVX1 U712 ( .A(n362), .Y(n664) );
  AND2X1 U713 ( .A(n768), .B(n775), .Y(n769) );
  INVX1 U714 ( .A(n769), .Y(n665) );
  AND2X1 U715 ( .A(n773), .B(n139), .Y(n767) );
  INVX1 U716 ( .A(n767), .Y(n666) );
  AND2X1 U717 ( .A(n761), .B(n296), .Y(n361) );
  INVX1 U718 ( .A(n361), .Y(n667) );
  BUFX2 U719 ( .A(oddBuffer[52]), .Y(n668) );
  BUFX2 U720 ( .A(oddBuffer[51]), .Y(n669) );
  BUFX2 U721 ( .A(oddBuffer[50]), .Y(n670) );
  BUFX2 U722 ( .A(oddBuffer[49]), .Y(n671) );
  BUFX2 U723 ( .A(oddBuffer[48]), .Y(n672) );
  BUFX2 U724 ( .A(oddBuffer[55]), .Y(n673) );
  BUFX2 U725 ( .A(oddBufferFull), .Y(n674) );
  AND2X1 U726 ( .A(n781), .B(n788), .Y(n782) );
  INVX1 U727 ( .A(n782), .Y(n675) );
  AND2X1 U728 ( .A(dataIn[39]), .B(n361), .Y(n336) );
  INVX1 U729 ( .A(n336), .Y(n676) );
  AND2X1 U730 ( .A(dataIn[12]), .B(n748), .Y(n309) );
  INVX1 U731 ( .A(n309), .Y(n677) );
  AND2X1 U732 ( .A(dataIn[1]), .B(n361), .Y(n298) );
  INVX1 U733 ( .A(n298), .Y(n678) );
  AND2X1 U734 ( .A(dataIn[0]), .B(n361), .Y(n297) );
  INVX1 U735 ( .A(n297), .Y(n679) );
  BUFX2 U736 ( .A(oddBuffer[63]), .Y(n680) );
  BUFX2 U737 ( .A(oddBuffer[61]), .Y(n681) );
  BUFX2 U738 ( .A(oddBuffer[60]), .Y(n682) );
  BUFX2 U739 ( .A(oddBuffer[59]), .Y(n683) );
  BUFX2 U740 ( .A(oddBuffer[58]), .Y(n684) );
  BUFX2 U741 ( .A(oddBuffer[57]), .Y(n685) );
  BUFX2 U742 ( .A(oddBuffer[56]), .Y(n686) );
  BUFX2 U743 ( .A(oddBuffer[47]), .Y(n687) );
  BUFX2 U744 ( .A(oddBuffer[46]), .Y(n688) );
  BUFX2 U745 ( .A(oddBuffer[45]), .Y(n689) );
  BUFX2 U746 ( .A(oddBuffer[44]), .Y(n690) );
  BUFX2 U747 ( .A(oddBuffer[43]), .Y(n691) );
  BUFX2 U748 ( .A(oddBuffer[42]), .Y(n692) );
  BUFX2 U749 ( .A(oddBuffer[41]), .Y(n693) );
  BUFX2 U750 ( .A(oddBuffer[40]), .Y(n694) );
  BUFX2 U751 ( .A(oddBuffer[39]), .Y(n695) );
  BUFX2 U752 ( .A(oddBuffer[38]), .Y(n696) );
  BUFX2 U753 ( .A(oddBuffer[37]), .Y(n697) );
  BUFX2 U754 ( .A(oddBuffer[36]), .Y(n698) );
  BUFX2 U755 ( .A(oddBuffer[35]), .Y(n699) );
  BUFX2 U756 ( .A(oddBuffer[34]), .Y(n700) );
  BUFX2 U757 ( .A(oddBuffer[33]), .Y(n701) );
  BUFX2 U758 ( .A(oddBuffer[32]), .Y(n702) );
  BUFX2 U759 ( .A(oddBuffer[31]), .Y(n703) );
  BUFX2 U760 ( .A(oddBuffer[30]), .Y(n704) );
  BUFX2 U761 ( .A(oddBuffer[29]), .Y(n705) );
  BUFX2 U762 ( .A(oddBuffer[28]), .Y(n706) );
  BUFX2 U763 ( .A(oddBuffer[27]), .Y(n707) );
  BUFX2 U764 ( .A(oddBuffer[26]), .Y(n708) );
  BUFX2 U765 ( .A(oddBuffer[25]), .Y(n709) );
  BUFX2 U766 ( .A(oddBuffer[24]), .Y(n710) );
  BUFX2 U767 ( .A(oddBuffer[23]), .Y(n711) );
  BUFX2 U768 ( .A(oddBuffer[22]), .Y(n712) );
  BUFX2 U769 ( .A(oddBuffer[21]), .Y(n713) );
  BUFX2 U770 ( .A(oddBuffer[20]), .Y(n714) );
  BUFX2 U771 ( .A(oddBuffer[19]), .Y(n715) );
  BUFX2 U772 ( .A(oddBuffer[18]), .Y(n716) );
  BUFX2 U773 ( .A(oddBuffer[17]), .Y(n717) );
  BUFX2 U774 ( .A(oddBuffer[16]), .Y(n718) );
  BUFX2 U775 ( .A(oddBuffer[15]), .Y(n719) );
  BUFX2 U776 ( .A(oddBuffer[14]), .Y(n720) );
  BUFX2 U777 ( .A(oddBuffer[13]), .Y(n721) );
  BUFX2 U778 ( .A(oddBuffer[12]), .Y(n722) );
  BUFX2 U779 ( .A(oddBuffer[11]), .Y(n723) );
  BUFX2 U780 ( .A(oddBuffer[10]), .Y(n724) );
  BUFX2 U781 ( .A(oddBuffer[9]), .Y(n725) );
  BUFX2 U782 ( .A(oddBuffer[8]), .Y(n726) );
  BUFX2 U783 ( .A(oddBuffer[7]), .Y(n727) );
  BUFX2 U784 ( .A(oddBuffer[6]), .Y(n728) );
  BUFX2 U785 ( .A(oddBuffer[5]), .Y(n729) );
  BUFX2 U786 ( .A(oddBuffer[4]), .Y(n730) );
  BUFX2 U787 ( .A(oddBuffer[3]), .Y(n731) );
  BUFX2 U788 ( .A(oddBuffer[2]), .Y(n732) );
  BUFX2 U789 ( .A(oddBuffer[1]), .Y(n733) );
  BUFX2 U790 ( .A(oddBuffer[0]), .Y(n734) );
  BUFX2 U791 ( .A(evenBuffer[53]), .Y(n735) );
  BUFX2 U792 ( .A(evenBuffer[52]), .Y(n736) );
  BUFX2 U793 ( .A(evenBuffer[51]), .Y(n737) );
  BUFX2 U794 ( .A(evenBuffer[50]), .Y(n738) );
  BUFX2 U795 ( .A(evenBuffer[49]), .Y(n739) );
  BUFX2 U796 ( .A(evenBuffer[48]), .Y(n740) );
  BUFX2 U797 ( .A(evenBuffer[55]), .Y(n741) );
  BUFX2 U798 ( .A(evenBufferFull), .Y(n742) );
  BUFX2 U799 ( .A(evenBuffer[54]), .Y(n743) );
  BUFX2 U800 ( .A(n412), .Y(n744) );
  INVX1 U801 ( .A(n430), .Y(n745) );
  INVX1 U802 ( .A(n667), .Y(n748) );
  INVX1 U803 ( .A(n765), .Y(n756) );
  INVX1 U804 ( .A(n764), .Y(n761) );
  INVX1 U805 ( .A(n766), .Y(n762) );
  INVX1 U806 ( .A(n766), .Y(n763) );
  INVX1 U807 ( .A(n764), .Y(n760) );
  INVX1 U808 ( .A(n764), .Y(n759) );
  INVX1 U809 ( .A(n765), .Y(n758) );
  INVX1 U810 ( .A(n765), .Y(n757) );
  AND2X1 U811 ( .A(n747), .B(n766), .Y(n746) );
  INVX1 U812 ( .A(n746), .Y(n410) );
  INVX1 U813 ( .A(n753), .Y(n764) );
  INVX1 U814 ( .A(n753), .Y(n765) );
  INVX1 U815 ( .A(n744), .Y(n747) );
  INVX1 U816 ( .A(n755), .Y(n753) );
  INVX1 U817 ( .A(n754), .Y(n766) );
  INVX1 U818 ( .A(n755), .Y(n754) );
  INVX1 U819 ( .A(polarity), .Y(n755) );
  INVX1 U820 ( .A(reset), .Y(n751) );
  INVX1 U821 ( .A(reset), .Y(n749) );
  INVX1 U822 ( .A(reset), .Y(n750) );
  INVX1 U823 ( .A(n452), .Y(dataOut[48]) );
  INVX1 U824 ( .A(n451), .Y(dataOut[49]) );
  INVX1 U825 ( .A(n449), .Y(dataOut[50]) );
  INVX1 U826 ( .A(n448), .Y(dataOut[51]) );
  INVX1 U827 ( .A(n447), .Y(dataOut[52]) );
  INVX1 U828 ( .A(n446), .Y(dataOut[53]) );
  INVX1 U829 ( .A(n296), .Y(n752) );
  INVX1 U830 ( .A(dataIn[48]), .Y(n926) );
  INVX1 U831 ( .A(dataIn[49]), .Y(n925) );
  INVX1 U832 ( .A(dataIn[50]), .Y(n924) );
  INVX1 U833 ( .A(dataIn[51]), .Y(n923) );
  INVX1 U834 ( .A(dataIn[52]), .Y(n922) );
  INVX1 U835 ( .A(dataIn[53]), .Y(n921) );
  INVX1 U836 ( .A(dataIn[54]), .Y(n920) );
  INVX1 U837 ( .A(dataIn[55]), .Y(n919) );
  INVX1 U838 ( .A(n684), .Y(n804) );
  INVX1 U839 ( .A(n683), .Y(n803) );
  INVX1 U840 ( .A(n682), .Y(n802) );
  INVX1 U841 ( .A(n681), .Y(n801) );
  INVX1 U842 ( .A(n680), .Y(n799) );
  INVX1 U843 ( .A(n722), .Y(n850) );
  INVX1 U844 ( .A(n721), .Y(n849) );
  INVX1 U845 ( .A(n720), .Y(n848) );
  INVX1 U846 ( .A(n719), .Y(n847) );
  INVX1 U847 ( .A(n718), .Y(n846) );
  INVX1 U848 ( .A(n717), .Y(n845) );
  INVX1 U849 ( .A(n716), .Y(n844) );
  INVX1 U850 ( .A(n715), .Y(n843) );
  INVX1 U851 ( .A(n714), .Y(n842) );
  INVX1 U852 ( .A(n713), .Y(n841) );
  INVX1 U853 ( .A(n712), .Y(n840) );
  INVX1 U854 ( .A(n711), .Y(n839) );
  INVX1 U855 ( .A(n710), .Y(n838) );
  INVX1 U856 ( .A(n733), .Y(n861) );
  INVX1 U857 ( .A(n732), .Y(n860) );
  INVX1 U858 ( .A(n731), .Y(n859) );
  INVX1 U859 ( .A(n730), .Y(n858) );
  INVX1 U860 ( .A(n729), .Y(n857) );
  INVX1 U861 ( .A(n728), .Y(n856) );
  INVX1 U862 ( .A(n727), .Y(n855) );
  INVX1 U863 ( .A(n726), .Y(n854) );
  INVX1 U864 ( .A(n725), .Y(n853) );
  INVX1 U865 ( .A(n724), .Y(n852) );
  INVX1 U866 ( .A(n723), .Y(n851) );
  INVX1 U867 ( .A(n445), .Y(dataOut[54]) );
  INVX1 U868 ( .A(n734), .Y(n862) );
  INVX1 U869 ( .A(n709), .Y(n837) );
  INVX1 U870 ( .A(n708), .Y(n836) );
  INVX1 U871 ( .A(n707), .Y(n835) );
  INVX1 U872 ( .A(n706), .Y(n834) );
  INVX1 U873 ( .A(n705), .Y(n833) );
  INVX1 U874 ( .A(n704), .Y(n832) );
  INVX1 U875 ( .A(n703), .Y(n831) );
  INVX1 U876 ( .A(n702), .Y(n830) );
  INVX1 U877 ( .A(n701), .Y(n829) );
  INVX1 U878 ( .A(n700), .Y(n828) );
  INVX1 U879 ( .A(n699), .Y(n827) );
  INVX1 U880 ( .A(n698), .Y(n826) );
  INVX1 U881 ( .A(n697), .Y(n825) );
  INVX1 U882 ( .A(n696), .Y(n824) );
  INVX1 U883 ( .A(n695), .Y(n823) );
  INVX1 U884 ( .A(n694), .Y(n822) );
  INVX1 U885 ( .A(n693), .Y(n821) );
  INVX1 U886 ( .A(n692), .Y(n820) );
  INVX1 U887 ( .A(n691), .Y(n819) );
  INVX1 U888 ( .A(n690), .Y(n818) );
  INVX1 U889 ( .A(n689), .Y(n817) );
  INVX1 U890 ( .A(n688), .Y(n816) );
  INVX1 U891 ( .A(n687), .Y(n815) );
  INVX1 U892 ( .A(n686), .Y(n806) );
  INVX1 U893 ( .A(n685), .Y(n805) );
  INVX1 U894 ( .A(n444), .Y(dataOut[55]) );
  INVX1 U895 ( .A(n742), .Y(n798) );
  INVX1 U896 ( .A(n674), .Y(n797) );
  INVX1 U897 ( .A(n345), .Y(n796) );
  INVX1 U898 ( .A(n346), .Y(n795) );
  INVX1 U899 ( .A(n347), .Y(n794) );
  INVX1 U900 ( .A(n348), .Y(n793) );
  INVX1 U901 ( .A(n349), .Y(n792) );
  INVX1 U902 ( .A(n350), .Y(n791) );
  INVX1 U903 ( .A(n351), .Y(n790) );
  INVX1 U904 ( .A(n352), .Y(n789) );
  INVX1 U905 ( .A(n657), .Y(n800) );
  INVX1 U906 ( .A(n644), .Y(n864) );
  INVX1 U907 ( .A(n740), .Y(n139) );
  INVX1 U908 ( .A(n672), .Y(n150) );
  INVX1 U909 ( .A(n739), .Y(n773) );
  INVX1 U910 ( .A(n738), .Y(n774) );
  INVX1 U911 ( .A(n737), .Y(n775) );
  INVX1 U912 ( .A(n736), .Y(n776) );
  INVX1 U913 ( .A(n735), .Y(n777) );
  INVX1 U914 ( .A(n671), .Y(n784) );
  INVX1 U915 ( .A(n670), .Y(n785) );
  INVX1 U916 ( .A(n669), .Y(n786) );
  INVX1 U917 ( .A(n668), .Y(n787) );
  INVX1 U918 ( .A(n653), .Y(n788) );
  INVX1 U919 ( .A(evenBuffer[0]), .Y(n918) );
  INVX1 U920 ( .A(evenBuffer[1]), .Y(n917) );
  INVX1 U921 ( .A(evenBuffer[2]), .Y(n916) );
  INVX1 U922 ( .A(evenBuffer[3]), .Y(n915) );
  INVX1 U923 ( .A(evenBuffer[4]), .Y(n914) );
  INVX1 U924 ( .A(evenBuffer[5]), .Y(n913) );
  INVX1 U925 ( .A(evenBuffer[6]), .Y(n912) );
  INVX1 U926 ( .A(evenBuffer[7]), .Y(n911) );
  INVX1 U927 ( .A(evenBuffer[8]), .Y(n910) );
  INVX1 U928 ( .A(evenBuffer[9]), .Y(n909) );
  INVX1 U929 ( .A(evenBuffer[10]), .Y(n908) );
  INVX1 U930 ( .A(evenBuffer[11]), .Y(n907) );
  INVX1 U931 ( .A(evenBuffer[12]), .Y(n906) );
  INVX1 U932 ( .A(evenBuffer[13]), .Y(n905) );
  INVX1 U933 ( .A(evenBuffer[14]), .Y(n904) );
  INVX1 U934 ( .A(evenBuffer[15]), .Y(n903) );
  INVX1 U935 ( .A(evenBuffer[16]), .Y(n902) );
  INVX1 U936 ( .A(evenBuffer[17]), .Y(n901) );
  INVX1 U937 ( .A(evenBuffer[18]), .Y(n900) );
  INVX1 U938 ( .A(evenBuffer[19]), .Y(n899) );
  INVX1 U939 ( .A(evenBuffer[20]), .Y(n898) );
  INVX1 U940 ( .A(evenBuffer[21]), .Y(n897) );
  INVX1 U941 ( .A(evenBuffer[22]), .Y(n896) );
  INVX1 U942 ( .A(evenBuffer[23]), .Y(n895) );
  INVX1 U943 ( .A(evenBuffer[24]), .Y(n894) );
  INVX1 U944 ( .A(evenBuffer[25]), .Y(n893) );
  INVX1 U945 ( .A(evenBuffer[26]), .Y(n892) );
  INVX1 U946 ( .A(evenBuffer[27]), .Y(n891) );
  INVX1 U947 ( .A(evenBuffer[28]), .Y(n890) );
  INVX1 U948 ( .A(evenBuffer[29]), .Y(n889) );
  INVX1 U949 ( .A(evenBuffer[30]), .Y(n888) );
  INVX1 U950 ( .A(evenBuffer[31]), .Y(n887) );
  INVX1 U951 ( .A(evenBuffer[32]), .Y(n886) );
  INVX1 U952 ( .A(evenBuffer[33]), .Y(n885) );
  INVX1 U953 ( .A(evenBuffer[34]), .Y(n884) );
  INVX1 U954 ( .A(evenBuffer[35]), .Y(n883) );
  INVX1 U955 ( .A(evenBuffer[36]), .Y(n882) );
  INVX1 U956 ( .A(evenBuffer[37]), .Y(n881) );
  INVX1 U957 ( .A(evenBuffer[38]), .Y(n880) );
  INVX1 U958 ( .A(evenBuffer[39]), .Y(n879) );
  INVX1 U959 ( .A(evenBuffer[40]), .Y(n878) );
  INVX1 U960 ( .A(evenBuffer[41]), .Y(n877) );
  INVX1 U961 ( .A(evenBuffer[42]), .Y(n876) );
  INVX1 U962 ( .A(evenBuffer[43]), .Y(n875) );
  INVX1 U963 ( .A(evenBuffer[44]), .Y(n874) );
  INVX1 U964 ( .A(evenBuffer[45]), .Y(n873) );
  INVX1 U965 ( .A(evenBuffer[46]), .Y(n872) );
  INVX1 U966 ( .A(evenBuffer[47]), .Y(n871) );
  INVX1 U967 ( .A(evenBuffer[56]), .Y(n870) );
  INVX1 U968 ( .A(evenBuffer[57]), .Y(n869) );
  INVX1 U969 ( .A(evenBuffer[58]), .Y(n868) );
  INVX1 U970 ( .A(evenBuffer[59]), .Y(n867) );
  INVX1 U971 ( .A(evenBuffer[60]), .Y(n866) );
  INVX1 U972 ( .A(evenBuffer[61]), .Y(n865) );
  INVX1 U973 ( .A(evenBuffer[63]), .Y(n863) );
  OAI21X1 U974 ( .A(n139), .B(n773), .C(n666), .Y(n140) );
  OAI21X1 U975 ( .A(n767), .B(n774), .C(n655), .Y(n141) );
  OAI21X1 U976 ( .A(n768), .B(n775), .C(n665), .Y(n142) );
  OAI21X1 U977 ( .A(n769), .B(n776), .C(n642), .Y(n143) );
  OAI21X1 U978 ( .A(n770), .B(n777), .C(n658), .Y(n144) );
  XNOR2X1 U979 ( .A(n743), .B(n658), .Y(n145) );
  XNOR2X1 U980 ( .A(n741), .B(n772), .Y(n146) );
  OAI21X1 U981 ( .A(n150), .B(n784), .C(n656), .Y(n151) );
  OAI21X1 U982 ( .A(n778), .B(n785), .C(n643), .Y(n152) );
  OAI21X1 U983 ( .A(n779), .B(n786), .C(n654), .Y(n153) );
  OAI21X1 U984 ( .A(n780), .B(n787), .C(n631), .Y(n154) );
  OAI21X1 U985 ( .A(n781), .B(n788), .C(n675), .Y(n155) );
  XNOR2X1 U986 ( .A(n645), .B(n675), .Y(n156) );
  XNOR2X1 U987 ( .A(n673), .B(n783), .Y(n157) );
endmodule


module outputBuffer_2 ( clk, reset, polarity, inputBufferRequest, dataIn0, 
        dataIn1, sendOut, readyOut, dataOut, InputBufferGrant );
  input [1:0] inputBufferRequest;
  input [63:0] dataIn0;
  input [63:0] dataIn1;
  output [63:0] dataOut;
  output [1:0] InputBufferGrant;
  input clk, reset, polarity, readyOut;
  output sendOut;
  wire   evenBufferFull, oddBufferFull, priorityRegEven, priorityRegOdd, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n340, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n132, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908;
  wire   [63:0] evenBuffer;
  wire   [63:0] oddBuffer;

  DFFSR evenBufferFull_reg ( .D(n621), .CLK(clk), .R(n758), .S(1'b1), .Q(
        evenBufferFull) );
  DFFSR priorityRegEven_reg ( .D(n619), .CLK(clk), .R(n758), .S(1'b1), .Q(
        priorityRegEven) );
  DFFSR priorityRegOdd_reg ( .D(n618), .CLK(clk), .R(n758), .S(1'b1), .Q(
        priorityRegOdd) );
  DFFSR oddBufferFull_reg ( .D(n620), .CLK(clk), .R(n757), .S(1'b1), .Q(
        oddBufferFull) );
  DFFSR oddBuffer_reg_63_ ( .D(n554), .CLK(clk), .R(n758), .S(1'b1), .Q(
        oddBuffer[63]) );
  DFFSR oddBuffer_reg_62_ ( .D(n555), .CLK(clk), .R(n758), .S(1'b1), .Q(
        oddBuffer[62]) );
  DFFSR oddBuffer_reg_61_ ( .D(n556), .CLK(clk), .R(n757), .S(1'b1), .Q(
        oddBuffer[61]) );
  DFFSR oddBuffer_reg_60_ ( .D(n557), .CLK(clk), .R(n756), .S(1'b1), .Q(
        oddBuffer[60]) );
  DFFSR oddBuffer_reg_59_ ( .D(n558), .CLK(clk), .R(n758), .S(1'b1), .Q(
        oddBuffer[59]) );
  DFFSR oddBuffer_reg_58_ ( .D(n559), .CLK(clk), .R(n756), .S(1'b1), .Q(
        oddBuffer[58]) );
  DFFSR oddBuffer_reg_57_ ( .D(n560), .CLK(clk), .R(n757), .S(1'b1), .Q(
        oddBuffer[57]) );
  DFFSR oddBuffer_reg_56_ ( .D(n561), .CLK(clk), .R(n756), .S(1'b1), .Q(
        oddBuffer[56]) );
  DFFSR oddBuffer_reg_55_ ( .D(n562), .CLK(clk), .R(n757), .S(1'b1), .Q(
        oddBuffer[55]) );
  DFFSR oddBuffer_reg_54_ ( .D(n563), .CLK(clk), .R(n757), .S(1'b1), .Q(
        oddBuffer[54]) );
  DFFSR oddBuffer_reg_53_ ( .D(n564), .CLK(clk), .R(n757), .S(1'b1), .Q(
        oddBuffer[53]) );
  DFFSR oddBuffer_reg_52_ ( .D(n565), .CLK(clk), .R(n758), .S(1'b1), .Q(
        oddBuffer[52]) );
  DFFSR oddBuffer_reg_51_ ( .D(n566), .CLK(clk), .R(n756), .S(1'b1), .Q(
        oddBuffer[51]) );
  DFFSR oddBuffer_reg_50_ ( .D(n567), .CLK(clk), .R(n757), .S(1'b1), .Q(
        oddBuffer[50]) );
  DFFSR oddBuffer_reg_49_ ( .D(n568), .CLK(clk), .R(n758), .S(1'b1), .Q(
        oddBuffer[49]) );
  DFFSR oddBuffer_reg_48_ ( .D(n569), .CLK(clk), .R(n757), .S(1'b1), .Q(
        oddBuffer[48]) );
  DFFSR oddBuffer_reg_47_ ( .D(n570), .CLK(clk), .R(n756), .S(1'b1), .Q(
        oddBuffer[47]) );
  DFFSR oddBuffer_reg_46_ ( .D(n571), .CLK(clk), .R(n757), .S(1'b1), .Q(
        oddBuffer[46]) );
  DFFSR oddBuffer_reg_45_ ( .D(n572), .CLK(clk), .R(n758), .S(1'b1), .Q(
        oddBuffer[45]) );
  DFFSR oddBuffer_reg_44_ ( .D(n573), .CLK(clk), .R(n756), .S(1'b1), .Q(
        oddBuffer[44]) );
  DFFSR oddBuffer_reg_43_ ( .D(n574), .CLK(clk), .R(n756), .S(1'b1), .Q(
        oddBuffer[43]) );
  DFFSR oddBuffer_reg_42_ ( .D(n575), .CLK(clk), .R(n757), .S(1'b1), .Q(
        oddBuffer[42]) );
  DFFSR oddBuffer_reg_41_ ( .D(n576), .CLK(clk), .R(n756), .S(1'b1), .Q(
        oddBuffer[41]) );
  DFFSR oddBuffer_reg_40_ ( .D(n577), .CLK(clk), .R(n756), .S(1'b1), .Q(
        oddBuffer[40]) );
  DFFSR oddBuffer_reg_39_ ( .D(n578), .CLK(clk), .R(n757), .S(1'b1), .Q(
        oddBuffer[39]) );
  DFFSR oddBuffer_reg_38_ ( .D(n579), .CLK(clk), .R(n758), .S(1'b1), .Q(
        oddBuffer[38]) );
  DFFSR oddBuffer_reg_37_ ( .D(n580), .CLK(clk), .R(n758), .S(1'b1), .Q(
        oddBuffer[37]) );
  DFFSR oddBuffer_reg_36_ ( .D(n581), .CLK(clk), .R(n756), .S(1'b1), .Q(
        oddBuffer[36]) );
  DFFSR oddBuffer_reg_35_ ( .D(n582), .CLK(clk), .R(n758), .S(1'b1), .Q(
        oddBuffer[35]) );
  DFFSR oddBuffer_reg_34_ ( .D(n583), .CLK(clk), .R(n756), .S(1'b1), .Q(
        oddBuffer[34]) );
  DFFSR oddBuffer_reg_33_ ( .D(n584), .CLK(clk), .R(n758), .S(1'b1), .Q(
        oddBuffer[33]) );
  DFFSR oddBuffer_reg_32_ ( .D(n585), .CLK(clk), .R(n758), .S(1'b1), .Q(
        oddBuffer[32]) );
  DFFSR oddBuffer_reg_31_ ( .D(n586), .CLK(clk), .R(n757), .S(1'b1), .Q(
        oddBuffer[31]) );
  DFFSR oddBuffer_reg_30_ ( .D(n587), .CLK(clk), .R(n758), .S(1'b1), .Q(
        oddBuffer[30]) );
  DFFSR oddBuffer_reg_29_ ( .D(n588), .CLK(clk), .R(n757), .S(1'b1), .Q(
        oddBuffer[29]) );
  DFFSR oddBuffer_reg_28_ ( .D(n589), .CLK(clk), .R(n758), .S(1'b1), .Q(
        oddBuffer[28]) );
  DFFSR oddBuffer_reg_27_ ( .D(n590), .CLK(clk), .R(n756), .S(1'b1), .Q(
        oddBuffer[27]) );
  DFFSR oddBuffer_reg_26_ ( .D(n591), .CLK(clk), .R(n756), .S(1'b1), .Q(
        oddBuffer[26]) );
  DFFSR oddBuffer_reg_25_ ( .D(n592), .CLK(clk), .R(n758), .S(1'b1), .Q(
        oddBuffer[25]) );
  DFFSR oddBuffer_reg_24_ ( .D(n593), .CLK(clk), .R(n757), .S(1'b1), .Q(
        oddBuffer[24]) );
  DFFSR oddBuffer_reg_23_ ( .D(n594), .CLK(clk), .R(n758), .S(1'b1), .Q(
        oddBuffer[23]) );
  DFFSR oddBuffer_reg_22_ ( .D(n595), .CLK(clk), .R(n756), .S(1'b1), .Q(
        oddBuffer[22]) );
  DFFSR oddBuffer_reg_21_ ( .D(n596), .CLK(clk), .R(n756), .S(1'b1), .Q(
        oddBuffer[21]) );
  DFFSR oddBuffer_reg_20_ ( .D(n597), .CLK(clk), .R(n757), .S(1'b1), .Q(
        oddBuffer[20]) );
  DFFSR oddBuffer_reg_19_ ( .D(n598), .CLK(clk), .R(n758), .S(1'b1), .Q(
        oddBuffer[19]) );
  DFFSR oddBuffer_reg_18_ ( .D(n599), .CLK(clk), .R(n756), .S(1'b1), .Q(
        oddBuffer[18]) );
  DFFSR oddBuffer_reg_17_ ( .D(n600), .CLK(clk), .R(n756), .S(1'b1), .Q(
        oddBuffer[17]) );
  DFFSR oddBuffer_reg_16_ ( .D(n601), .CLK(clk), .R(n757), .S(1'b1), .Q(
        oddBuffer[16]) );
  DFFSR oddBuffer_reg_15_ ( .D(n602), .CLK(clk), .R(n758), .S(1'b1), .Q(
        oddBuffer[15]) );
  DFFSR oddBuffer_reg_14_ ( .D(n603), .CLK(clk), .R(n756), .S(1'b1), .Q(
        oddBuffer[14]) );
  DFFSR oddBuffer_reg_13_ ( .D(n604), .CLK(clk), .R(n757), .S(1'b1), .Q(
        oddBuffer[13]) );
  DFFSR oddBuffer_reg_12_ ( .D(n605), .CLK(clk), .R(n757), .S(1'b1), .Q(
        oddBuffer[12]) );
  DFFSR oddBuffer_reg_11_ ( .D(n606), .CLK(clk), .R(n758), .S(1'b1), .Q(
        oddBuffer[11]) );
  DFFSR oddBuffer_reg_10_ ( .D(n607), .CLK(clk), .R(n756), .S(1'b1), .Q(
        oddBuffer[10]) );
  DFFSR oddBuffer_reg_9_ ( .D(n608), .CLK(clk), .R(n758), .S(1'b1), .Q(
        oddBuffer[9]) );
  DFFSR oddBuffer_reg_8_ ( .D(n609), .CLK(clk), .R(n757), .S(1'b1), .Q(
        oddBuffer[8]) );
  DFFSR oddBuffer_reg_7_ ( .D(n610), .CLK(clk), .R(n758), .S(1'b1), .Q(
        oddBuffer[7]) );
  DFFSR oddBuffer_reg_6_ ( .D(n611), .CLK(clk), .R(n756), .S(1'b1), .Q(
        oddBuffer[6]) );
  DFFSR oddBuffer_reg_5_ ( .D(n612), .CLK(clk), .R(n757), .S(1'b1), .Q(
        oddBuffer[5]) );
  DFFSR oddBuffer_reg_4_ ( .D(n613), .CLK(clk), .R(n758), .S(1'b1), .Q(
        oddBuffer[4]) );
  DFFSR oddBuffer_reg_3_ ( .D(n614), .CLK(clk), .R(n756), .S(1'b1), .Q(
        oddBuffer[3]) );
  DFFSR oddBuffer_reg_2_ ( .D(n615), .CLK(clk), .R(n757), .S(1'b1), .Q(
        oddBuffer[2]) );
  DFFSR oddBuffer_reg_1_ ( .D(n616), .CLK(clk), .R(n758), .S(1'b1), .Q(
        oddBuffer[1]) );
  DFFSR oddBuffer_reg_0_ ( .D(n617), .CLK(clk), .R(n756), .S(1'b1), .Q(
        oddBuffer[0]) );
  DFFSR evenBuffer_reg_63_ ( .D(n490), .CLK(clk), .R(n757), .S(1'b1), .Q(
        evenBuffer[63]) );
  DFFSR evenBuffer_reg_62_ ( .D(n491), .CLK(clk), .R(n758), .S(1'b1), .Q(
        evenBuffer[62]) );
  DFFSR evenBuffer_reg_61_ ( .D(n492), .CLK(clk), .R(n756), .S(1'b1), .Q(
        evenBuffer[61]) );
  DFFSR evenBuffer_reg_60_ ( .D(n493), .CLK(clk), .R(n757), .S(1'b1), .Q(
        evenBuffer[60]) );
  DFFSR evenBuffer_reg_59_ ( .D(n494), .CLK(clk), .R(n757), .S(1'b1), .Q(
        evenBuffer[59]) );
  DFFSR evenBuffer_reg_58_ ( .D(n495), .CLK(clk), .R(n758), .S(1'b1), .Q(
        evenBuffer[58]) );
  DFFSR evenBuffer_reg_57_ ( .D(n496), .CLK(clk), .R(n757), .S(1'b1), .Q(
        evenBuffer[57]) );
  DFFSR evenBuffer_reg_56_ ( .D(n497), .CLK(clk), .R(n756), .S(1'b1), .Q(
        evenBuffer[56]) );
  DFFSR evenBuffer_reg_55_ ( .D(n498), .CLK(clk), .R(n756), .S(1'b1), .Q(
        evenBuffer[55]) );
  DFFSR evenBuffer_reg_54_ ( .D(n499), .CLK(clk), .R(n758), .S(1'b1), .Q(
        evenBuffer[54]) );
  DFFSR evenBuffer_reg_53_ ( .D(n500), .CLK(clk), .R(n756), .S(1'b1), .Q(
        evenBuffer[53]) );
  DFFSR evenBuffer_reg_52_ ( .D(n501), .CLK(clk), .R(n756), .S(1'b1), .Q(
        evenBuffer[52]) );
  DFFSR evenBuffer_reg_51_ ( .D(n502), .CLK(clk), .R(n758), .S(1'b1), .Q(
        evenBuffer[51]) );
  DFFSR evenBuffer_reg_50_ ( .D(n503), .CLK(clk), .R(n756), .S(1'b1), .Q(
        evenBuffer[50]) );
  DFFSR evenBuffer_reg_49_ ( .D(n504), .CLK(clk), .R(n757), .S(1'b1), .Q(
        evenBuffer[49]) );
  DFFSR evenBuffer_reg_48_ ( .D(n505), .CLK(clk), .R(n757), .S(1'b1), .Q(
        evenBuffer[48]) );
  DFFSR evenBuffer_reg_47_ ( .D(n506), .CLK(clk), .R(n758), .S(1'b1), .Q(
        evenBuffer[47]) );
  DFFSR evenBuffer_reg_46_ ( .D(n507), .CLK(clk), .R(n756), .S(1'b1), .Q(
        evenBuffer[46]) );
  DFFSR evenBuffer_reg_45_ ( .D(n508), .CLK(clk), .R(n757), .S(1'b1), .Q(
        evenBuffer[45]) );
  DFFSR evenBuffer_reg_44_ ( .D(n509), .CLK(clk), .R(n756), .S(1'b1), .Q(
        evenBuffer[44]) );
  DFFSR evenBuffer_reg_43_ ( .D(n510), .CLK(clk), .R(n757), .S(1'b1), .Q(
        evenBuffer[43]) );
  DFFSR evenBuffer_reg_42_ ( .D(n511), .CLK(clk), .R(n756), .S(1'b1), .Q(
        evenBuffer[42]) );
  DFFSR evenBuffer_reg_41_ ( .D(n512), .CLK(clk), .R(n758), .S(1'b1), .Q(
        evenBuffer[41]) );
  DFFSR evenBuffer_reg_40_ ( .D(n513), .CLK(clk), .R(n756), .S(1'b1), .Q(
        evenBuffer[40]) );
  DFFSR evenBuffer_reg_39_ ( .D(n514), .CLK(clk), .R(n758), .S(1'b1), .Q(
        evenBuffer[39]) );
  DFFSR evenBuffer_reg_38_ ( .D(n515), .CLK(clk), .R(n757), .S(1'b1), .Q(
        evenBuffer[38]) );
  DFFSR evenBuffer_reg_37_ ( .D(n516), .CLK(clk), .R(n757), .S(1'b1), .Q(
        evenBuffer[37]) );
  DFFSR evenBuffer_reg_36_ ( .D(n517), .CLK(clk), .R(n757), .S(1'b1), .Q(
        evenBuffer[36]) );
  DFFSR evenBuffer_reg_35_ ( .D(n518), .CLK(clk), .R(n758), .S(1'b1), .Q(
        evenBuffer[35]) );
  DFFSR evenBuffer_reg_34_ ( .D(n519), .CLK(clk), .R(n758), .S(1'b1), .Q(
        evenBuffer[34]) );
  DFFSR evenBuffer_reg_33_ ( .D(n520), .CLK(clk), .R(n758), .S(1'b1), .Q(
        evenBuffer[33]) );
  DFFSR evenBuffer_reg_32_ ( .D(n521), .CLK(clk), .R(n758), .S(1'b1), .Q(
        evenBuffer[32]) );
  DFFSR evenBuffer_reg_31_ ( .D(n522), .CLK(clk), .R(n758), .S(1'b1), .Q(
        evenBuffer[31]) );
  DFFSR evenBuffer_reg_30_ ( .D(n523), .CLK(clk), .R(n758), .S(1'b1), .Q(
        evenBuffer[30]) );
  DFFSR evenBuffer_reg_29_ ( .D(n524), .CLK(clk), .R(n758), .S(1'b1), .Q(
        evenBuffer[29]) );
  DFFSR evenBuffer_reg_28_ ( .D(n525), .CLK(clk), .R(n758), .S(1'b1), .Q(
        evenBuffer[28]) );
  DFFSR evenBuffer_reg_27_ ( .D(n526), .CLK(clk), .R(n758), .S(1'b1), .Q(
        evenBuffer[27]) );
  DFFSR evenBuffer_reg_26_ ( .D(n527), .CLK(clk), .R(n758), .S(1'b1), .Q(
        evenBuffer[26]) );
  DFFSR evenBuffer_reg_25_ ( .D(n528), .CLK(clk), .R(n758), .S(1'b1), .Q(
        evenBuffer[25]) );
  DFFSR evenBuffer_reg_24_ ( .D(n529), .CLK(clk), .R(n758), .S(1'b1), .Q(
        evenBuffer[24]) );
  DFFSR evenBuffer_reg_23_ ( .D(n530), .CLK(clk), .R(n757), .S(1'b1), .Q(
        evenBuffer[23]) );
  DFFSR evenBuffer_reg_22_ ( .D(n531), .CLK(clk), .R(n757), .S(1'b1), .Q(
        evenBuffer[22]) );
  DFFSR evenBuffer_reg_21_ ( .D(n532), .CLK(clk), .R(n757), .S(1'b1), .Q(
        evenBuffer[21]) );
  DFFSR evenBuffer_reg_20_ ( .D(n533), .CLK(clk), .R(n757), .S(1'b1), .Q(
        evenBuffer[20]) );
  DFFSR evenBuffer_reg_19_ ( .D(n534), .CLK(clk), .R(n757), .S(1'b1), .Q(
        evenBuffer[19]) );
  DFFSR evenBuffer_reg_18_ ( .D(n535), .CLK(clk), .R(n757), .S(1'b1), .Q(
        evenBuffer[18]) );
  DFFSR evenBuffer_reg_17_ ( .D(n536), .CLK(clk), .R(n757), .S(1'b1), .Q(
        evenBuffer[17]) );
  DFFSR evenBuffer_reg_16_ ( .D(n537), .CLK(clk), .R(n757), .S(1'b1), .Q(
        evenBuffer[16]) );
  DFFSR evenBuffer_reg_15_ ( .D(n538), .CLK(clk), .R(n757), .S(1'b1), .Q(
        evenBuffer[15]) );
  DFFSR evenBuffer_reg_14_ ( .D(n539), .CLK(clk), .R(n757), .S(1'b1), .Q(
        evenBuffer[14]) );
  DFFSR evenBuffer_reg_13_ ( .D(n540), .CLK(clk), .R(n757), .S(1'b1), .Q(
        evenBuffer[13]) );
  DFFSR evenBuffer_reg_12_ ( .D(n541), .CLK(clk), .R(n757), .S(1'b1), .Q(
        evenBuffer[12]) );
  DFFSR evenBuffer_reg_11_ ( .D(n542), .CLK(clk), .R(n756), .S(1'b1), .Q(
        evenBuffer[11]) );
  DFFSR evenBuffer_reg_10_ ( .D(n543), .CLK(clk), .R(n756), .S(1'b1), .Q(
        evenBuffer[10]) );
  DFFSR evenBuffer_reg_9_ ( .D(n544), .CLK(clk), .R(n756), .S(1'b1), .Q(
        evenBuffer[9]) );
  DFFSR evenBuffer_reg_8_ ( .D(n545), .CLK(clk), .R(n756), .S(1'b1), .Q(
        evenBuffer[8]) );
  DFFSR evenBuffer_reg_7_ ( .D(n546), .CLK(clk), .R(n756), .S(1'b1), .Q(
        evenBuffer[7]) );
  DFFSR evenBuffer_reg_6_ ( .D(n547), .CLK(clk), .R(n756), .S(1'b1), .Q(
        evenBuffer[6]) );
  DFFSR evenBuffer_reg_5_ ( .D(n548), .CLK(clk), .R(n756), .S(1'b1), .Q(
        evenBuffer[5]) );
  DFFSR evenBuffer_reg_4_ ( .D(n549), .CLK(clk), .R(n756), .S(1'b1), .Q(
        evenBuffer[4]) );
  DFFSR evenBuffer_reg_3_ ( .D(n550), .CLK(clk), .R(n756), .S(1'b1), .Q(
        evenBuffer[3]) );
  DFFSR evenBuffer_reg_2_ ( .D(n551), .CLK(clk), .R(n756), .S(1'b1), .Q(
        evenBuffer[2]) );
  DFFSR evenBuffer_reg_1_ ( .D(n552), .CLK(clk), .R(n756), .S(1'b1), .Q(
        evenBuffer[1]) );
  DFFSR evenBuffer_reg_0_ ( .D(n553), .CLK(clk), .R(n756), .S(1'b1), .Q(
        evenBuffer[0]) );
  OAI21X1 U275 ( .A(n272), .B(n845), .C(n262), .Y(n490) );
  AOI22X1 U276 ( .A(dataIn1[63]), .B(n762), .C(dataIn0[63]), .D(n761), .Y(n273) );
  OAI21X1 U277 ( .A(n272), .B(n846), .C(n261), .Y(n491) );
  AOI22X1 U278 ( .A(dataIn1[62]), .B(n762), .C(dataIn0[62]), .D(n761), .Y(n276) );
  OAI21X1 U279 ( .A(n272), .B(n847), .C(n260), .Y(n492) );
  AOI22X1 U280 ( .A(dataIn1[61]), .B(n762), .C(dataIn0[61]), .D(n761), .Y(n277) );
  OAI21X1 U281 ( .A(n272), .B(n848), .C(n259), .Y(n493) );
  AOI22X1 U282 ( .A(dataIn1[60]), .B(n762), .C(dataIn0[60]), .D(n761), .Y(n278) );
  OAI21X1 U283 ( .A(n272), .B(n849), .C(n258), .Y(n494) );
  AOI22X1 U284 ( .A(dataIn1[59]), .B(n762), .C(dataIn0[59]), .D(n761), .Y(n279) );
  OAI21X1 U285 ( .A(n272), .B(n850), .C(n257), .Y(n495) );
  AOI22X1 U286 ( .A(dataIn1[58]), .B(n762), .C(dataIn0[58]), .D(n761), .Y(n280) );
  OAI21X1 U287 ( .A(n272), .B(n851), .C(n256), .Y(n496) );
  AOI22X1 U288 ( .A(dataIn1[57]), .B(n762), .C(dataIn0[57]), .D(n761), .Y(n281) );
  OAI21X1 U289 ( .A(n272), .B(n852), .C(n255), .Y(n497) );
  AOI22X1 U290 ( .A(dataIn1[56]), .B(n762), .C(dataIn0[56]), .D(n761), .Y(n282) );
  OAI21X1 U291 ( .A(n272), .B(n853), .C(n254), .Y(n498) );
  AOI22X1 U292 ( .A(dataIn1[55]), .B(n762), .C(dataIn0[55]), .D(n761), .Y(n283) );
  OAI21X1 U293 ( .A(n272), .B(n854), .C(n253), .Y(n499) );
  AOI22X1 U294 ( .A(dataIn1[54]), .B(n762), .C(dataIn0[54]), .D(n761), .Y(n284) );
  OAI21X1 U295 ( .A(n272), .B(n855), .C(n252), .Y(n500) );
  AOI22X1 U296 ( .A(dataIn1[53]), .B(n762), .C(dataIn0[53]), .D(n761), .Y(n285) );
  OAI21X1 U297 ( .A(n272), .B(n856), .C(n251), .Y(n501) );
  AOI22X1 U298 ( .A(dataIn1[52]), .B(n762), .C(dataIn0[52]), .D(n761), .Y(n286) );
  OAI21X1 U299 ( .A(n272), .B(n857), .C(n250), .Y(n502) );
  AOI22X1 U300 ( .A(dataIn1[51]), .B(n762), .C(dataIn0[51]), .D(n761), .Y(n287) );
  OAI21X1 U301 ( .A(n272), .B(n858), .C(n249), .Y(n503) );
  AOI22X1 U302 ( .A(dataIn1[50]), .B(n762), .C(dataIn0[50]), .D(n761), .Y(n288) );
  OAI21X1 U303 ( .A(n272), .B(n859), .C(n248), .Y(n504) );
  AOI22X1 U304 ( .A(dataIn1[49]), .B(n762), .C(dataIn0[49]), .D(n761), .Y(n289) );
  OAI21X1 U305 ( .A(n272), .B(n860), .C(n247), .Y(n505) );
  AOI22X1 U306 ( .A(dataIn1[48]), .B(n762), .C(dataIn0[48]), .D(n761), .Y(n290) );
  OAI21X1 U307 ( .A(n272), .B(n861), .C(n246), .Y(n506) );
  AOI22X1 U308 ( .A(dataIn1[47]), .B(n762), .C(dataIn0[47]), .D(n761), .Y(n291) );
  OAI21X1 U309 ( .A(n272), .B(n862), .C(n245), .Y(n507) );
  AOI22X1 U310 ( .A(dataIn1[46]), .B(n762), .C(dataIn0[46]), .D(n761), .Y(n292) );
  OAI21X1 U311 ( .A(n272), .B(n863), .C(n244), .Y(n508) );
  AOI22X1 U312 ( .A(dataIn1[45]), .B(n762), .C(dataIn0[45]), .D(n761), .Y(n293) );
  OAI21X1 U313 ( .A(n272), .B(n864), .C(n243), .Y(n509) );
  AOI22X1 U314 ( .A(dataIn1[44]), .B(n762), .C(dataIn0[44]), .D(n761), .Y(n294) );
  OAI21X1 U315 ( .A(n272), .B(n865), .C(n242), .Y(n510) );
  AOI22X1 U316 ( .A(dataIn1[43]), .B(n762), .C(dataIn0[43]), .D(n761), .Y(n295) );
  OAI21X1 U317 ( .A(n272), .B(n866), .C(n241), .Y(n511) );
  AOI22X1 U318 ( .A(dataIn1[42]), .B(n762), .C(dataIn0[42]), .D(n761), .Y(n296) );
  OAI21X1 U319 ( .A(n272), .B(n867), .C(n240), .Y(n512) );
  AOI22X1 U320 ( .A(dataIn1[41]), .B(n762), .C(dataIn0[41]), .D(n761), .Y(n297) );
  OAI21X1 U321 ( .A(n272), .B(n868), .C(n239), .Y(n513) );
  AOI22X1 U322 ( .A(dataIn1[40]), .B(n762), .C(dataIn0[40]), .D(n761), .Y(n298) );
  OAI21X1 U323 ( .A(n272), .B(n869), .C(n238), .Y(n514) );
  AOI22X1 U324 ( .A(dataIn1[39]), .B(n762), .C(dataIn0[39]), .D(n761), .Y(n299) );
  OAI21X1 U325 ( .A(n272), .B(n870), .C(n237), .Y(n515) );
  AOI22X1 U326 ( .A(dataIn1[38]), .B(n762), .C(dataIn0[38]), .D(n761), .Y(n300) );
  OAI21X1 U327 ( .A(n272), .B(n871), .C(n236), .Y(n516) );
  AOI22X1 U328 ( .A(dataIn1[37]), .B(n762), .C(dataIn0[37]), .D(n761), .Y(n301) );
  OAI21X1 U329 ( .A(n272), .B(n872), .C(n235), .Y(n517) );
  AOI22X1 U330 ( .A(dataIn1[36]), .B(n762), .C(dataIn0[36]), .D(n761), .Y(n302) );
  OAI21X1 U331 ( .A(n272), .B(n873), .C(n234), .Y(n518) );
  AOI22X1 U332 ( .A(dataIn1[35]), .B(n762), .C(dataIn0[35]), .D(n761), .Y(n303) );
  OAI21X1 U333 ( .A(n272), .B(n874), .C(n233), .Y(n519) );
  AOI22X1 U334 ( .A(dataIn1[34]), .B(n762), .C(dataIn0[34]), .D(n761), .Y(n304) );
  OAI21X1 U335 ( .A(n272), .B(n875), .C(n232), .Y(n520) );
  AOI22X1 U336 ( .A(dataIn1[33]), .B(n762), .C(dataIn0[33]), .D(n761), .Y(n305) );
  OAI21X1 U337 ( .A(n272), .B(n876), .C(n231), .Y(n521) );
  AOI22X1 U338 ( .A(dataIn1[32]), .B(n762), .C(dataIn0[32]), .D(n761), .Y(n306) );
  OAI21X1 U339 ( .A(n272), .B(n877), .C(n230), .Y(n522) );
  AOI22X1 U340 ( .A(dataIn1[31]), .B(n762), .C(dataIn0[31]), .D(n761), .Y(n307) );
  OAI21X1 U341 ( .A(n272), .B(n878), .C(n229), .Y(n523) );
  AOI22X1 U342 ( .A(dataIn1[30]), .B(n762), .C(dataIn0[30]), .D(n761), .Y(n308) );
  OAI21X1 U343 ( .A(n272), .B(n879), .C(n228), .Y(n524) );
  AOI22X1 U344 ( .A(dataIn1[29]), .B(n762), .C(dataIn0[29]), .D(n761), .Y(n309) );
  OAI21X1 U345 ( .A(n272), .B(n880), .C(n227), .Y(n525) );
  AOI22X1 U346 ( .A(dataIn1[28]), .B(n762), .C(dataIn0[28]), .D(n761), .Y(n310) );
  OAI21X1 U347 ( .A(n272), .B(n881), .C(n226), .Y(n526) );
  AOI22X1 U348 ( .A(dataIn1[27]), .B(n762), .C(dataIn0[27]), .D(n761), .Y(n311) );
  OAI21X1 U349 ( .A(n272), .B(n882), .C(n225), .Y(n527) );
  AOI22X1 U350 ( .A(dataIn1[26]), .B(n762), .C(dataIn0[26]), .D(n761), .Y(n312) );
  OAI21X1 U351 ( .A(n272), .B(n883), .C(n224), .Y(n528) );
  AOI22X1 U352 ( .A(dataIn1[25]), .B(n762), .C(dataIn0[25]), .D(n761), .Y(n313) );
  OAI21X1 U353 ( .A(n272), .B(n884), .C(n223), .Y(n529) );
  AOI22X1 U354 ( .A(dataIn1[24]), .B(n762), .C(dataIn0[24]), .D(n761), .Y(n314) );
  OAI21X1 U355 ( .A(n272), .B(n885), .C(n222), .Y(n530) );
  AOI22X1 U356 ( .A(dataIn1[23]), .B(n762), .C(dataIn0[23]), .D(n761), .Y(n315) );
  OAI21X1 U357 ( .A(n272), .B(n886), .C(n221), .Y(n531) );
  AOI22X1 U358 ( .A(dataIn1[22]), .B(n762), .C(dataIn0[22]), .D(n761), .Y(n316) );
  OAI21X1 U359 ( .A(n272), .B(n887), .C(n220), .Y(n532) );
  AOI22X1 U360 ( .A(dataIn1[21]), .B(n762), .C(dataIn0[21]), .D(n761), .Y(n317) );
  OAI21X1 U361 ( .A(n272), .B(n888), .C(n219), .Y(n533) );
  AOI22X1 U362 ( .A(dataIn1[20]), .B(n762), .C(dataIn0[20]), .D(n761), .Y(n318) );
  OAI21X1 U363 ( .A(n272), .B(n889), .C(n218), .Y(n534) );
  AOI22X1 U364 ( .A(dataIn1[19]), .B(n762), .C(dataIn0[19]), .D(n761), .Y(n319) );
  OAI21X1 U365 ( .A(n272), .B(n890), .C(n217), .Y(n535) );
  AOI22X1 U366 ( .A(dataIn1[18]), .B(n762), .C(dataIn0[18]), .D(n761), .Y(n320) );
  OAI21X1 U367 ( .A(n272), .B(n891), .C(n216), .Y(n536) );
  AOI22X1 U368 ( .A(dataIn1[17]), .B(n762), .C(dataIn0[17]), .D(n761), .Y(n321) );
  OAI21X1 U369 ( .A(n272), .B(n892), .C(n215), .Y(n537) );
  AOI22X1 U370 ( .A(dataIn1[16]), .B(n762), .C(dataIn0[16]), .D(n761), .Y(n322) );
  OAI21X1 U371 ( .A(n272), .B(n893), .C(n214), .Y(n538) );
  AOI22X1 U372 ( .A(dataIn1[15]), .B(n762), .C(dataIn0[15]), .D(n761), .Y(n323) );
  OAI21X1 U373 ( .A(n272), .B(n894), .C(n213), .Y(n539) );
  AOI22X1 U374 ( .A(dataIn1[14]), .B(n762), .C(dataIn0[14]), .D(n761), .Y(n324) );
  OAI21X1 U375 ( .A(n272), .B(n895), .C(n212), .Y(n540) );
  AOI22X1 U376 ( .A(dataIn1[13]), .B(n762), .C(dataIn0[13]), .D(n761), .Y(n325) );
  OAI21X1 U377 ( .A(n272), .B(n896), .C(n211), .Y(n541) );
  AOI22X1 U378 ( .A(dataIn1[12]), .B(n762), .C(dataIn0[12]), .D(n761), .Y(n326) );
  OAI21X1 U379 ( .A(n272), .B(n897), .C(n210), .Y(n542) );
  AOI22X1 U380 ( .A(dataIn1[11]), .B(n762), .C(dataIn0[11]), .D(n761), .Y(n327) );
  OAI21X1 U381 ( .A(n272), .B(n898), .C(n209), .Y(n543) );
  AOI22X1 U382 ( .A(dataIn1[10]), .B(n762), .C(dataIn0[10]), .D(n761), .Y(n328) );
  OAI21X1 U383 ( .A(n272), .B(n899), .C(n208), .Y(n544) );
  AOI22X1 U384 ( .A(dataIn1[9]), .B(n762), .C(dataIn0[9]), .D(n761), .Y(n329)
         );
  OAI21X1 U385 ( .A(n272), .B(n900), .C(n207), .Y(n545) );
  AOI22X1 U386 ( .A(dataIn1[8]), .B(n762), .C(dataIn0[8]), .D(n761), .Y(n330)
         );
  OAI21X1 U387 ( .A(n272), .B(n901), .C(n206), .Y(n546) );
  AOI22X1 U388 ( .A(dataIn1[7]), .B(n762), .C(dataIn0[7]), .D(n761), .Y(n331)
         );
  OAI21X1 U389 ( .A(n272), .B(n902), .C(n205), .Y(n547) );
  AOI22X1 U390 ( .A(dataIn1[6]), .B(n762), .C(dataIn0[6]), .D(n761), .Y(n332)
         );
  OAI21X1 U391 ( .A(n272), .B(n903), .C(n204), .Y(n548) );
  AOI22X1 U392 ( .A(dataIn1[5]), .B(n762), .C(dataIn0[5]), .D(n761), .Y(n333)
         );
  OAI21X1 U393 ( .A(n272), .B(n904), .C(n203), .Y(n549) );
  AOI22X1 U394 ( .A(dataIn1[4]), .B(n762), .C(dataIn0[4]), .D(n761), .Y(n334)
         );
  OAI21X1 U395 ( .A(n272), .B(n905), .C(n202), .Y(n550) );
  AOI22X1 U396 ( .A(dataIn1[3]), .B(n762), .C(dataIn0[3]), .D(n761), .Y(n335)
         );
  OAI21X1 U397 ( .A(n272), .B(n906), .C(n201), .Y(n551) );
  AOI22X1 U398 ( .A(dataIn1[2]), .B(n762), .C(dataIn0[2]), .D(n761), .Y(n336)
         );
  OAI21X1 U399 ( .A(n272), .B(n907), .C(n200), .Y(n552) );
  AOI22X1 U400 ( .A(dataIn1[1]), .B(n762), .C(dataIn0[1]), .D(n761), .Y(n337)
         );
  OAI21X1 U401 ( .A(n272), .B(n908), .C(n199), .Y(n553) );
  AOI22X1 U402 ( .A(dataIn1[0]), .B(n762), .C(dataIn0[0]), .D(n761), .Y(n338)
         );
  OAI21X1 U405 ( .A(n342), .B(n781), .C(n198), .Y(n554) );
  AOI22X1 U406 ( .A(n760), .B(dataIn1[63]), .C(n759), .D(dataIn0[63]), .Y(n343) );
  OAI21X1 U407 ( .A(n342), .B(n782), .C(n197), .Y(n555) );
  AOI22X1 U408 ( .A(n760), .B(dataIn1[62]), .C(n759), .D(dataIn0[62]), .Y(n346) );
  OAI21X1 U409 ( .A(n342), .B(n783), .C(n196), .Y(n556) );
  AOI22X1 U410 ( .A(n760), .B(dataIn1[61]), .C(n759), .D(dataIn0[61]), .Y(n347) );
  OAI21X1 U411 ( .A(n342), .B(n784), .C(n195), .Y(n557) );
  AOI22X1 U412 ( .A(n760), .B(dataIn1[60]), .C(n759), .D(dataIn0[60]), .Y(n348) );
  OAI21X1 U413 ( .A(n342), .B(n785), .C(n194), .Y(n558) );
  AOI22X1 U414 ( .A(n760), .B(dataIn1[59]), .C(n759), .D(dataIn0[59]), .Y(n349) );
  OAI21X1 U415 ( .A(n342), .B(n786), .C(n193), .Y(n559) );
  AOI22X1 U416 ( .A(n760), .B(dataIn1[58]), .C(n759), .D(dataIn0[58]), .Y(n350) );
  OAI21X1 U417 ( .A(n342), .B(n787), .C(n192), .Y(n560) );
  AOI22X1 U418 ( .A(n760), .B(dataIn1[57]), .C(n759), .D(dataIn0[57]), .Y(n351) );
  OAI21X1 U419 ( .A(n342), .B(n788), .C(n191), .Y(n561) );
  AOI22X1 U420 ( .A(n760), .B(dataIn1[56]), .C(n759), .D(dataIn0[56]), .Y(n352) );
  OAI21X1 U421 ( .A(n342), .B(n789), .C(n190), .Y(n562) );
  AOI22X1 U422 ( .A(n760), .B(dataIn1[55]), .C(n759), .D(dataIn0[55]), .Y(n353) );
  OAI21X1 U423 ( .A(n342), .B(n790), .C(n189), .Y(n563) );
  AOI22X1 U424 ( .A(n760), .B(dataIn1[54]), .C(n759), .D(dataIn0[54]), .Y(n354) );
  OAI21X1 U425 ( .A(n342), .B(n791), .C(n188), .Y(n564) );
  AOI22X1 U426 ( .A(n760), .B(dataIn1[53]), .C(n759), .D(dataIn0[53]), .Y(n355) );
  OAI21X1 U427 ( .A(n342), .B(n792), .C(n187), .Y(n565) );
  AOI22X1 U428 ( .A(n760), .B(dataIn1[52]), .C(n759), .D(dataIn0[52]), .Y(n356) );
  OAI21X1 U429 ( .A(n342), .B(n793), .C(n186), .Y(n566) );
  AOI22X1 U430 ( .A(n760), .B(dataIn1[51]), .C(n759), .D(dataIn0[51]), .Y(n357) );
  OAI21X1 U431 ( .A(n342), .B(n794), .C(n185), .Y(n567) );
  AOI22X1 U432 ( .A(n760), .B(dataIn1[50]), .C(n759), .D(dataIn0[50]), .Y(n358) );
  OAI21X1 U433 ( .A(n342), .B(n795), .C(n184), .Y(n568) );
  AOI22X1 U434 ( .A(n760), .B(dataIn1[49]), .C(n759), .D(dataIn0[49]), .Y(n359) );
  OAI21X1 U435 ( .A(n342), .B(n796), .C(n183), .Y(n569) );
  AOI22X1 U436 ( .A(n760), .B(dataIn1[48]), .C(n759), .D(dataIn0[48]), .Y(n360) );
  OAI21X1 U437 ( .A(n342), .B(n797), .C(n182), .Y(n570) );
  AOI22X1 U438 ( .A(n760), .B(dataIn1[47]), .C(n759), .D(dataIn0[47]), .Y(n361) );
  OAI21X1 U439 ( .A(n342), .B(n798), .C(n181), .Y(n571) );
  AOI22X1 U440 ( .A(n760), .B(dataIn1[46]), .C(n759), .D(dataIn0[46]), .Y(n362) );
  OAI21X1 U441 ( .A(n342), .B(n799), .C(n180), .Y(n572) );
  AOI22X1 U442 ( .A(n760), .B(dataIn1[45]), .C(n759), .D(dataIn0[45]), .Y(n363) );
  OAI21X1 U443 ( .A(n342), .B(n800), .C(n179), .Y(n573) );
  AOI22X1 U444 ( .A(n760), .B(dataIn1[44]), .C(n759), .D(dataIn0[44]), .Y(n364) );
  OAI21X1 U445 ( .A(n342), .B(n801), .C(n178), .Y(n574) );
  AOI22X1 U446 ( .A(n760), .B(dataIn1[43]), .C(n759), .D(dataIn0[43]), .Y(n365) );
  OAI21X1 U447 ( .A(n342), .B(n802), .C(n177), .Y(n575) );
  AOI22X1 U448 ( .A(n760), .B(dataIn1[42]), .C(n759), .D(dataIn0[42]), .Y(n366) );
  OAI21X1 U449 ( .A(n342), .B(n803), .C(n176), .Y(n576) );
  AOI22X1 U450 ( .A(n760), .B(dataIn1[41]), .C(n759), .D(dataIn0[41]), .Y(n367) );
  OAI21X1 U451 ( .A(n342), .B(n804), .C(n175), .Y(n577) );
  AOI22X1 U452 ( .A(n760), .B(dataIn1[40]), .C(n759), .D(dataIn0[40]), .Y(n368) );
  OAI21X1 U453 ( .A(n342), .B(n805), .C(n174), .Y(n578) );
  AOI22X1 U454 ( .A(n760), .B(dataIn1[39]), .C(n759), .D(dataIn0[39]), .Y(n369) );
  OAI21X1 U455 ( .A(n342), .B(n806), .C(n173), .Y(n579) );
  AOI22X1 U456 ( .A(n760), .B(dataIn1[38]), .C(n759), .D(dataIn0[38]), .Y(n370) );
  OAI21X1 U457 ( .A(n342), .B(n807), .C(n172), .Y(n580) );
  AOI22X1 U458 ( .A(n760), .B(dataIn1[37]), .C(n759), .D(dataIn0[37]), .Y(n371) );
  OAI21X1 U459 ( .A(n342), .B(n808), .C(n171), .Y(n581) );
  AOI22X1 U460 ( .A(n760), .B(dataIn1[36]), .C(n759), .D(dataIn0[36]), .Y(n372) );
  OAI21X1 U461 ( .A(n342), .B(n809), .C(n170), .Y(n582) );
  AOI22X1 U462 ( .A(n760), .B(dataIn1[35]), .C(n759), .D(dataIn0[35]), .Y(n373) );
  OAI21X1 U463 ( .A(n342), .B(n810), .C(n169), .Y(n583) );
  AOI22X1 U464 ( .A(n760), .B(dataIn1[34]), .C(n759), .D(dataIn0[34]), .Y(n374) );
  OAI21X1 U465 ( .A(n342), .B(n811), .C(n168), .Y(n584) );
  AOI22X1 U466 ( .A(n760), .B(dataIn1[33]), .C(n759), .D(dataIn0[33]), .Y(n375) );
  OAI21X1 U467 ( .A(n342), .B(n812), .C(n167), .Y(n585) );
  AOI22X1 U468 ( .A(n760), .B(dataIn1[32]), .C(n759), .D(dataIn0[32]), .Y(n376) );
  OAI21X1 U469 ( .A(n342), .B(n813), .C(n166), .Y(n586) );
  AOI22X1 U470 ( .A(n760), .B(dataIn1[31]), .C(n759), .D(dataIn0[31]), .Y(n377) );
  OAI21X1 U471 ( .A(n342), .B(n814), .C(n165), .Y(n587) );
  AOI22X1 U472 ( .A(n760), .B(dataIn1[30]), .C(n759), .D(dataIn0[30]), .Y(n378) );
  OAI21X1 U473 ( .A(n342), .B(n815), .C(n164), .Y(n588) );
  AOI22X1 U474 ( .A(n760), .B(dataIn1[29]), .C(n759), .D(dataIn0[29]), .Y(n379) );
  OAI21X1 U475 ( .A(n342), .B(n816), .C(n163), .Y(n589) );
  AOI22X1 U476 ( .A(n760), .B(dataIn1[28]), .C(n759), .D(dataIn0[28]), .Y(n380) );
  OAI21X1 U477 ( .A(n342), .B(n817), .C(n162), .Y(n590) );
  AOI22X1 U478 ( .A(n760), .B(dataIn1[27]), .C(n759), .D(dataIn0[27]), .Y(n381) );
  OAI21X1 U479 ( .A(n342), .B(n818), .C(n161), .Y(n591) );
  AOI22X1 U480 ( .A(n760), .B(dataIn1[26]), .C(n759), .D(dataIn0[26]), .Y(n382) );
  OAI21X1 U481 ( .A(n342), .B(n819), .C(n160), .Y(n592) );
  AOI22X1 U482 ( .A(n760), .B(dataIn1[25]), .C(n759), .D(dataIn0[25]), .Y(n383) );
  OAI21X1 U483 ( .A(n342), .B(n820), .C(n159), .Y(n593) );
  AOI22X1 U484 ( .A(n760), .B(dataIn1[24]), .C(n759), .D(dataIn0[24]), .Y(n384) );
  OAI21X1 U485 ( .A(n342), .B(n821), .C(n158), .Y(n594) );
  AOI22X1 U486 ( .A(n760), .B(dataIn1[23]), .C(n759), .D(dataIn0[23]), .Y(n385) );
  OAI21X1 U487 ( .A(n342), .B(n822), .C(n157), .Y(n595) );
  AOI22X1 U488 ( .A(n760), .B(dataIn1[22]), .C(n759), .D(dataIn0[22]), .Y(n386) );
  OAI21X1 U489 ( .A(n342), .B(n823), .C(n156), .Y(n596) );
  AOI22X1 U490 ( .A(n760), .B(dataIn1[21]), .C(n759), .D(dataIn0[21]), .Y(n387) );
  OAI21X1 U491 ( .A(n342), .B(n824), .C(n155), .Y(n597) );
  AOI22X1 U492 ( .A(n760), .B(dataIn1[20]), .C(n759), .D(dataIn0[20]), .Y(n388) );
  OAI21X1 U493 ( .A(n342), .B(n825), .C(n154), .Y(n598) );
  AOI22X1 U494 ( .A(n760), .B(dataIn1[19]), .C(n759), .D(dataIn0[19]), .Y(n389) );
  OAI21X1 U495 ( .A(n342), .B(n826), .C(n153), .Y(n599) );
  AOI22X1 U496 ( .A(n760), .B(dataIn1[18]), .C(n759), .D(dataIn0[18]), .Y(n390) );
  OAI21X1 U497 ( .A(n342), .B(n827), .C(n152), .Y(n600) );
  AOI22X1 U498 ( .A(n760), .B(dataIn1[17]), .C(n759), .D(dataIn0[17]), .Y(n391) );
  OAI21X1 U499 ( .A(n342), .B(n828), .C(n151), .Y(n601) );
  AOI22X1 U500 ( .A(n760), .B(dataIn1[16]), .C(n759), .D(dataIn0[16]), .Y(n392) );
  OAI21X1 U501 ( .A(n342), .B(n829), .C(n150), .Y(n602) );
  AOI22X1 U502 ( .A(n760), .B(dataIn1[15]), .C(n759), .D(dataIn0[15]), .Y(n393) );
  OAI21X1 U503 ( .A(n342), .B(n830), .C(n149), .Y(n603) );
  AOI22X1 U504 ( .A(n760), .B(dataIn1[14]), .C(n759), .D(dataIn0[14]), .Y(n394) );
  OAI21X1 U505 ( .A(n342), .B(n831), .C(n148), .Y(n604) );
  AOI22X1 U506 ( .A(n760), .B(dataIn1[13]), .C(n759), .D(dataIn0[13]), .Y(n395) );
  OAI21X1 U507 ( .A(n342), .B(n832), .C(n147), .Y(n605) );
  AOI22X1 U508 ( .A(n760), .B(dataIn1[12]), .C(n759), .D(dataIn0[12]), .Y(n396) );
  OAI21X1 U509 ( .A(n342), .B(n833), .C(n146), .Y(n606) );
  AOI22X1 U510 ( .A(n760), .B(dataIn1[11]), .C(n759), .D(dataIn0[11]), .Y(n397) );
  OAI21X1 U511 ( .A(n342), .B(n834), .C(n145), .Y(n607) );
  AOI22X1 U512 ( .A(n760), .B(dataIn1[10]), .C(n759), .D(dataIn0[10]), .Y(n398) );
  OAI21X1 U513 ( .A(n342), .B(n835), .C(n144), .Y(n608) );
  AOI22X1 U514 ( .A(n760), .B(dataIn1[9]), .C(n759), .D(dataIn0[9]), .Y(n399)
         );
  OAI21X1 U515 ( .A(n342), .B(n836), .C(n143), .Y(n609) );
  AOI22X1 U516 ( .A(n760), .B(dataIn1[8]), .C(n759), .D(dataIn0[8]), .Y(n400)
         );
  OAI21X1 U517 ( .A(n342), .B(n837), .C(n142), .Y(n610) );
  AOI22X1 U518 ( .A(n760), .B(dataIn1[7]), .C(n759), .D(dataIn0[7]), .Y(n401)
         );
  OAI21X1 U519 ( .A(n342), .B(n838), .C(n141), .Y(n611) );
  AOI22X1 U520 ( .A(n760), .B(dataIn1[6]), .C(n759), .D(dataIn0[6]), .Y(n402)
         );
  OAI21X1 U521 ( .A(n342), .B(n839), .C(n140), .Y(n612) );
  AOI22X1 U522 ( .A(n760), .B(dataIn1[5]), .C(n759), .D(dataIn0[5]), .Y(n403)
         );
  OAI21X1 U523 ( .A(n342), .B(n840), .C(n139), .Y(n613) );
  AOI22X1 U524 ( .A(n760), .B(dataIn1[4]), .C(n759), .D(dataIn0[4]), .Y(n404)
         );
  OAI21X1 U525 ( .A(n342), .B(n841), .C(n138), .Y(n614) );
  AOI22X1 U526 ( .A(n760), .B(dataIn1[3]), .C(n759), .D(dataIn0[3]), .Y(n405)
         );
  OAI21X1 U527 ( .A(n342), .B(n842), .C(n137), .Y(n615) );
  AOI22X1 U528 ( .A(n760), .B(dataIn1[2]), .C(n759), .D(dataIn0[2]), .Y(n406)
         );
  OAI21X1 U529 ( .A(n342), .B(n843), .C(n136), .Y(n616) );
  AOI22X1 U530 ( .A(n760), .B(dataIn1[1]), .C(n759), .D(dataIn0[1]), .Y(n407)
         );
  OAI21X1 U531 ( .A(n342), .B(n844), .C(n135), .Y(n617) );
  AOI22X1 U532 ( .A(n760), .B(dataIn1[0]), .C(n759), .D(dataIn0[0]), .Y(n408)
         );
  XNOR2X1 U535 ( .A(n755), .B(n684), .Y(n618) );
  XNOR2X1 U537 ( .A(n687), .B(n688), .Y(n619) );
  NAND3X1 U539 ( .A(inputBufferRequest[1]), .B(n631), .C(inputBufferRequest[0]), .Y(n412) );
  OAI21X1 U540 ( .A(n780), .B(n342), .C(n753), .Y(n620) );
  OAI21X1 U542 ( .A(n765), .B(n685), .C(n629), .Y(n342) );
  OAI21X1 U544 ( .A(n777), .B(n272), .C(n754), .Y(n621) );
  OAI21X1 U546 ( .A(n765), .B(n413), .C(n628), .Y(n272) );
  OAI21X1 U549 ( .A(n765), .B(n780), .C(n686), .Y(n417) );
  OAI21X1 U552 ( .A(n765), .B(n835), .C(n661), .Y(dataOut[9]) );
  OAI21X1 U554 ( .A(n765), .B(n836), .C(n665), .Y(dataOut[8]) );
  OAI21X1 U556 ( .A(n765), .B(n837), .C(n670), .Y(dataOut[7]) );
  OAI21X1 U558 ( .A(n766), .B(n838), .C(n673), .Y(dataOut[6]) );
  OAI21X1 U560 ( .A(n766), .B(n781), .C(n637), .Y(dataOut[63]) );
  OAI21X1 U562 ( .A(n765), .B(n782), .C(n641), .Y(dataOut[62]) );
  OAI21X1 U564 ( .A(n766), .B(n783), .C(n645), .Y(dataOut[61]) );
  OAI21X1 U566 ( .A(n766), .B(n784), .C(n653), .Y(dataOut[60]) );
  OAI21X1 U568 ( .A(n766), .B(n839), .C(n677), .Y(dataOut[5]) );
  OAI21X1 U570 ( .A(n766), .B(n785), .C(n627), .Y(dataOut[59]) );
  OAI21X1 U572 ( .A(n767), .B(n786), .C(n626), .Y(dataOut[58]) );
  OAI21X1 U574 ( .A(n766), .B(n787), .C(n625), .Y(dataOut[57]) );
  OAI21X1 U576 ( .A(n767), .B(n788), .C(n624), .Y(dataOut[56]) );
  OAI21X1 U578 ( .A(n767), .B(n789), .C(n623), .Y(dataOut[55]) );
  OAI21X1 U580 ( .A(n765), .B(n790), .C(n634), .Y(dataOut[54]) );
  OAI21X1 U582 ( .A(n767), .B(n791), .C(n638), .Y(dataOut[53]) );
  OAI21X1 U584 ( .A(n767), .B(n792), .C(n646), .Y(dataOut[52]) );
  OAI21X1 U586 ( .A(n767), .B(n793), .C(n649), .Y(dataOut[51]) );
  OAI21X1 U588 ( .A(n767), .B(n794), .C(n642), .Y(dataOut[50]) );
  OAI21X1 U590 ( .A(n766), .B(n840), .C(n674), .Y(dataOut[4]) );
  OAI21X1 U592 ( .A(n767), .B(n795), .C(n657), .Y(dataOut[49]) );
  OAI21X1 U594 ( .A(n767), .B(n796), .C(n654), .Y(dataOut[48]) );
  OAI21X1 U596 ( .A(n768), .B(n797), .C(n666), .Y(dataOut[47]) );
  OAI21X1 U598 ( .A(n766), .B(n798), .C(n681), .Y(dataOut[46]) );
  OAI21X1 U600 ( .A(n768), .B(n799), .C(n662), .Y(dataOut[45]) );
  OAI21X1 U602 ( .A(n768), .B(n800), .C(n675), .Y(dataOut[44]) );
  OAI21X1 U604 ( .A(n767), .B(n801), .C(n622), .Y(dataOut[43]) );
  OAI21X1 U606 ( .A(n768), .B(n802), .C(n271), .Y(dataOut[42]) );
  OAI21X1 U608 ( .A(n768), .B(n803), .C(n270), .Y(dataOut[41]) );
  OAI21X1 U610 ( .A(n768), .B(n804), .C(n269), .Y(dataOut[40]) );
  OAI21X1 U612 ( .A(n768), .B(n841), .C(n682), .Y(dataOut[3]) );
  OAI21X1 U614 ( .A(n768), .B(n805), .C(n268), .Y(dataOut[39]) );
  OAI21X1 U616 ( .A(n767), .B(n806), .C(n635), .Y(dataOut[38]) );
  OAI21X1 U618 ( .A(n768), .B(n807), .C(n658), .Y(dataOut[37]) );
  OAI21X1 U620 ( .A(n769), .B(n808), .C(n639), .Y(dataOut[36]) );
  OAI21X1 U622 ( .A(n768), .B(n809), .C(n650), .Y(dataOut[35]) );
  OAI21X1 U624 ( .A(n769), .B(n810), .C(n643), .Y(dataOut[34]) );
  OAI21X1 U626 ( .A(n769), .B(n811), .C(n647), .Y(dataOut[33]) );
  OAI21X1 U628 ( .A(n768), .B(n812), .C(n667), .Y(dataOut[32]) );
  OAI21X1 U630 ( .A(n769), .B(n813), .C(n655), .Y(dataOut[31]) );
  OAI21X1 U632 ( .A(n769), .B(n814), .C(n663), .Y(dataOut[30]) );
  OAI21X1 U634 ( .A(n766), .B(n842), .C(n678), .Y(dataOut[2]) );
  OAI21X1 U636 ( .A(n768), .B(n815), .C(n267), .Y(dataOut[29]) );
  OAI21X1 U638 ( .A(n769), .B(n816), .C(n266), .Y(dataOut[28]) );
  OAI21X1 U640 ( .A(n769), .B(n817), .C(n265), .Y(dataOut[27]) );
  OAI21X1 U642 ( .A(n768), .B(n818), .C(n264), .Y(dataOut[26]) );
  OAI21X1 U644 ( .A(n768), .B(n819), .C(n263), .Y(dataOut[25]) );
  OAI21X1 U646 ( .A(n768), .B(n820), .C(n636), .Y(dataOut[24]) );
  OAI21X1 U648 ( .A(n768), .B(n821), .C(n640), .Y(dataOut[23]) );
  OAI21X1 U650 ( .A(n768), .B(n822), .C(n644), .Y(dataOut[22]) );
  OAI21X1 U652 ( .A(n768), .B(n823), .C(n648), .Y(dataOut[21]) );
  OAI21X1 U654 ( .A(n767), .B(n824), .C(n671), .Y(dataOut[20]) );
  OAI21X1 U656 ( .A(n767), .B(n843), .C(n683), .Y(dataOut[1]) );
  OAI21X1 U658 ( .A(n766), .B(n825), .C(n659), .Y(dataOut[19]) );
  OAI21X1 U660 ( .A(n766), .B(n826), .C(n651), .Y(dataOut[18]) );
  OAI21X1 U662 ( .A(n767), .B(n827), .C(n668), .Y(dataOut[17]) );
  OAI21X1 U664 ( .A(n767), .B(n828), .C(n676), .Y(dataOut[16]) );
  OAI21X1 U666 ( .A(n766), .B(n829), .C(n660), .Y(dataOut[15]) );
  OAI21X1 U668 ( .A(n766), .B(n830), .C(n664), .Y(dataOut[14]) );
  OAI21X1 U670 ( .A(n766), .B(n831), .C(n669), .Y(dataOut[13]) );
  OAI21X1 U672 ( .A(n765), .B(n832), .C(n652), .Y(dataOut[12]) );
  OAI21X1 U674 ( .A(n765), .B(n833), .C(n656), .Y(dataOut[11]) );
  OAI21X1 U676 ( .A(n765), .B(n834), .C(n672), .Y(dataOut[10]) );
  OAI21X1 U678 ( .A(n765), .B(n844), .C(n679), .Y(dataOut[0]) );
  OAI21X1 U681 ( .A(inputBufferRequest[0]), .B(n630), .C(n134), .Y(n483) );
  AOI22X1 U682 ( .A(n687), .B(n486), .C(n755), .D(n487), .Y(n485) );
  OAI21X1 U684 ( .A(inputBufferRequest[1]), .B(n630), .C(n132), .Y(n488) );
  AOI22X1 U685 ( .A(n486), .B(n778), .C(n487), .D(n779), .Y(n489) );
  AND2X1 U133 ( .A(n769), .B(n680), .Y(n418) );
  AND2X1 U135 ( .A(inputBufferRequest[1]), .B(n483), .Y(InputBufferGrant[1])
         );
  AND2X1 U136 ( .A(inputBufferRequest[0]), .B(n488), .Y(InputBufferGrant[0])
         );
  OR2X1 U137 ( .A(n753), .B(n633), .Y(n344) );
  OR2X1 U138 ( .A(n753), .B(n632), .Y(n345) );
  OR2X1 U139 ( .A(n754), .B(n633), .Y(n274) );
  OR2X1 U140 ( .A(n632), .B(n754), .Y(n275) );
  BUFX2 U141 ( .A(n489), .Y(n132) );
  BUFX2 U142 ( .A(n485), .Y(n134) );
  BUFX2 U143 ( .A(n408), .Y(n135) );
  BUFX2 U144 ( .A(n407), .Y(n136) );
  BUFX2 U145 ( .A(n406), .Y(n137) );
  BUFX2 U146 ( .A(n405), .Y(n138) );
  BUFX2 U147 ( .A(n404), .Y(n139) );
  BUFX2 U148 ( .A(n403), .Y(n140) );
  BUFX2 U149 ( .A(n402), .Y(n141) );
  BUFX2 U150 ( .A(n401), .Y(n142) );
  BUFX2 U151 ( .A(n400), .Y(n143) );
  BUFX2 U152 ( .A(n399), .Y(n144) );
  BUFX2 U153 ( .A(n398), .Y(n145) );
  BUFX2 U154 ( .A(n397), .Y(n146) );
  BUFX2 U155 ( .A(n396), .Y(n147) );
  BUFX2 U156 ( .A(n395), .Y(n148) );
  BUFX2 U157 ( .A(n394), .Y(n149) );
  BUFX2 U158 ( .A(n393), .Y(n150) );
  BUFX2 U159 ( .A(n392), .Y(n151) );
  BUFX2 U160 ( .A(n391), .Y(n152) );
  BUFX2 U161 ( .A(n390), .Y(n153) );
  BUFX2 U162 ( .A(n389), .Y(n154) );
  BUFX2 U163 ( .A(n388), .Y(n155) );
  BUFX2 U164 ( .A(n387), .Y(n156) );
  BUFX2 U165 ( .A(n386), .Y(n157) );
  BUFX2 U166 ( .A(n385), .Y(n158) );
  BUFX2 U167 ( .A(n384), .Y(n159) );
  BUFX2 U168 ( .A(n383), .Y(n160) );
  BUFX2 U169 ( .A(n382), .Y(n161) );
  BUFX2 U170 ( .A(n381), .Y(n162) );
  BUFX2 U171 ( .A(n380), .Y(n163) );
  BUFX2 U172 ( .A(n379), .Y(n164) );
  BUFX2 U173 ( .A(n378), .Y(n165) );
  BUFX2 U174 ( .A(n377), .Y(n166) );
  BUFX2 U175 ( .A(n376), .Y(n167) );
  BUFX2 U176 ( .A(n375), .Y(n168) );
  BUFX2 U177 ( .A(n374), .Y(n169) );
  BUFX2 U178 ( .A(n373), .Y(n170) );
  BUFX2 U179 ( .A(n372), .Y(n171) );
  BUFX2 U180 ( .A(n371), .Y(n172) );
  BUFX2 U181 ( .A(n370), .Y(n173) );
  BUFX2 U182 ( .A(n369), .Y(n174) );
  BUFX2 U183 ( .A(n368), .Y(n175) );
  BUFX2 U184 ( .A(n367), .Y(n176) );
  BUFX2 U185 ( .A(n366), .Y(n177) );
  BUFX2 U186 ( .A(n365), .Y(n178) );
  BUFX2 U187 ( .A(n364), .Y(n179) );
  BUFX2 U188 ( .A(n363), .Y(n180) );
  BUFX2 U189 ( .A(n362), .Y(n181) );
  BUFX2 U190 ( .A(n361), .Y(n182) );
  BUFX2 U191 ( .A(n360), .Y(n183) );
  BUFX2 U192 ( .A(n359), .Y(n184) );
  BUFX2 U193 ( .A(n358), .Y(n185) );
  BUFX2 U194 ( .A(n357), .Y(n186) );
  BUFX2 U195 ( .A(n356), .Y(n187) );
  BUFX2 U196 ( .A(n355), .Y(n188) );
  BUFX2 U197 ( .A(n354), .Y(n189) );
  BUFX2 U198 ( .A(n353), .Y(n190) );
  BUFX2 U199 ( .A(n352), .Y(n191) );
  BUFX2 U200 ( .A(n351), .Y(n192) );
  BUFX2 U201 ( .A(n350), .Y(n193) );
  BUFX2 U202 ( .A(n349), .Y(n194) );
  BUFX2 U203 ( .A(n348), .Y(n195) );
  BUFX2 U204 ( .A(n347), .Y(n196) );
  BUFX2 U205 ( .A(n346), .Y(n197) );
  BUFX2 U206 ( .A(n343), .Y(n198) );
  BUFX2 U207 ( .A(n338), .Y(n199) );
  BUFX2 U208 ( .A(n337), .Y(n200) );
  BUFX2 U209 ( .A(n336), .Y(n201) );
  BUFX2 U210 ( .A(n335), .Y(n202) );
  BUFX2 U211 ( .A(n334), .Y(n203) );
  BUFX2 U212 ( .A(n333), .Y(n204) );
  BUFX2 U213 ( .A(n332), .Y(n205) );
  BUFX2 U214 ( .A(n331), .Y(n206) );
  BUFX2 U215 ( .A(n330), .Y(n207) );
  BUFX2 U216 ( .A(n329), .Y(n208) );
  BUFX2 U217 ( .A(n328), .Y(n209) );
  BUFX2 U218 ( .A(n327), .Y(n210) );
  BUFX2 U219 ( .A(n326), .Y(n211) );
  BUFX2 U220 ( .A(n325), .Y(n212) );
  BUFX2 U221 ( .A(n324), .Y(n213) );
  BUFX2 U222 ( .A(n323), .Y(n214) );
  BUFX2 U223 ( .A(n322), .Y(n215) );
  BUFX2 U224 ( .A(n321), .Y(n216) );
  BUFX2 U225 ( .A(n320), .Y(n217) );
  BUFX2 U226 ( .A(n319), .Y(n218) );
  BUFX2 U227 ( .A(n318), .Y(n219) );
  BUFX2 U228 ( .A(n317), .Y(n220) );
  BUFX2 U229 ( .A(n316), .Y(n221) );
  BUFX2 U230 ( .A(n315), .Y(n222) );
  BUFX2 U231 ( .A(n314), .Y(n223) );
  BUFX2 U232 ( .A(n313), .Y(n224) );
  BUFX2 U233 ( .A(n312), .Y(n225) );
  BUFX2 U234 ( .A(n311), .Y(n226) );
  BUFX2 U235 ( .A(n310), .Y(n227) );
  BUFX2 U236 ( .A(n309), .Y(n228) );
  BUFX2 U237 ( .A(n308), .Y(n229) );
  BUFX2 U238 ( .A(n307), .Y(n230) );
  BUFX2 U239 ( .A(n306), .Y(n231) );
  BUFX2 U240 ( .A(n305), .Y(n232) );
  BUFX2 U241 ( .A(n304), .Y(n233) );
  BUFX2 U242 ( .A(n303), .Y(n234) );
  BUFX2 U243 ( .A(n302), .Y(n235) );
  BUFX2 U244 ( .A(n301), .Y(n236) );
  BUFX2 U245 ( .A(n300), .Y(n237) );
  BUFX2 U246 ( .A(n299), .Y(n238) );
  BUFX2 U247 ( .A(n298), .Y(n239) );
  BUFX2 U248 ( .A(n297), .Y(n240) );
  BUFX2 U249 ( .A(n296), .Y(n241) );
  BUFX2 U250 ( .A(n295), .Y(n242) );
  BUFX2 U251 ( .A(n294), .Y(n243) );
  BUFX2 U252 ( .A(n293), .Y(n244) );
  BUFX2 U253 ( .A(n292), .Y(n245) );
  BUFX2 U254 ( .A(n291), .Y(n246) );
  BUFX2 U255 ( .A(n290), .Y(n247) );
  BUFX2 U256 ( .A(n289), .Y(n248) );
  BUFX2 U257 ( .A(n288), .Y(n249) );
  BUFX2 U258 ( .A(n287), .Y(n250) );
  BUFX2 U259 ( .A(n286), .Y(n251) );
  BUFX2 U260 ( .A(n285), .Y(n252) );
  BUFX2 U261 ( .A(n284), .Y(n253) );
  BUFX2 U262 ( .A(n283), .Y(n254) );
  BUFX2 U263 ( .A(n282), .Y(n255) );
  BUFX2 U264 ( .A(n281), .Y(n256) );
  BUFX2 U265 ( .A(n280), .Y(n257) );
  BUFX2 U266 ( .A(n279), .Y(n258) );
  BUFX2 U267 ( .A(n278), .Y(n259) );
  BUFX2 U268 ( .A(n277), .Y(n260) );
  BUFX2 U269 ( .A(n276), .Y(n261) );
  BUFX2 U270 ( .A(n273), .Y(n262) );
  AND2X1 U271 ( .A(n727), .B(n770), .Y(n465) );
  INVX1 U272 ( .A(n465), .Y(n263) );
  AND2X1 U273 ( .A(n726), .B(n770), .Y(n464) );
  INVX1 U274 ( .A(n464), .Y(n264) );
  AND2X1 U403 ( .A(n725), .B(n770), .Y(n463) );
  INVX1 U404 ( .A(n463), .Y(n265) );
  AND2X1 U533 ( .A(n724), .B(n770), .Y(n462) );
  INVX1 U534 ( .A(n462), .Y(n266) );
  AND2X1 U536 ( .A(n723), .B(n770), .Y(n461) );
  INVX1 U538 ( .A(n461), .Y(n267) );
  AND2X1 U541 ( .A(n713), .B(n771), .Y(n450) );
  INVX1 U543 ( .A(n450), .Y(n268) );
  AND2X1 U545 ( .A(n712), .B(n771), .Y(n448) );
  INVX1 U547 ( .A(n448), .Y(n269) );
  AND2X1 U548 ( .A(n711), .B(n771), .Y(n447) );
  INVX1 U550 ( .A(n447), .Y(n270) );
  AND2X1 U551 ( .A(n710), .B(n771), .Y(n446) );
  INVX1 U553 ( .A(n446), .Y(n271) );
  AND2X1 U555 ( .A(n709), .B(n771), .Y(n445) );
  INVX1 U557 ( .A(n445), .Y(n622) );
  AND2X1 U559 ( .A(n697), .B(n772), .Y(n432) );
  INVX1 U561 ( .A(n432), .Y(n623) );
  AND2X1 U563 ( .A(n696), .B(n772), .Y(n431) );
  INVX1 U565 ( .A(n431), .Y(n624) );
  AND2X1 U567 ( .A(n695), .B(n772), .Y(n430) );
  INVX1 U569 ( .A(n430), .Y(n625) );
  AND2X1 U571 ( .A(n694), .B(n772), .Y(n429) );
  INVX1 U573 ( .A(n429), .Y(n626) );
  AND2X1 U575 ( .A(n693), .B(n772), .Y(n428) );
  INVX1 U577 ( .A(n428), .Y(n627) );
  AND2X1 U579 ( .A(sendOut), .B(n773), .Y(n416) );
  INVX1 U581 ( .A(n416), .Y(n628) );
  AND2X1 U583 ( .A(n769), .B(n631), .Y(n415) );
  INVX1 U585 ( .A(n415), .Y(n629) );
  OR2X1 U587 ( .A(n487), .B(n486), .Y(n484) );
  INVX1 U589 ( .A(n484), .Y(n630) );
  AND2X1 U591 ( .A(n633), .B(n632), .Y(n413) );
  INVX1 U593 ( .A(n413), .Y(n631) );
  INVX1 U595 ( .A(InputBufferGrant[0]), .Y(n632) );
  INVX1 U597 ( .A(InputBufferGrant[1]), .Y(n633) );
  AND2X1 U599 ( .A(n698), .B(n772), .Y(n433) );
  INVX1 U601 ( .A(n433), .Y(n634) );
  AND2X1 U603 ( .A(n714), .B(n771), .Y(n451) );
  INVX1 U605 ( .A(n451), .Y(n635) );
  AND2X1 U607 ( .A(n728), .B(n770), .Y(n466) );
  INVX1 U609 ( .A(n466), .Y(n636) );
  AND2X1 U611 ( .A(n689), .B(n773), .Y(n423) );
  INVX1 U613 ( .A(n423), .Y(n637) );
  AND2X1 U615 ( .A(n699), .B(n772), .Y(n434) );
  INVX1 U617 ( .A(n434), .Y(n638) );
  AND2X1 U619 ( .A(n716), .B(n771), .Y(n453) );
  INVX1 U621 ( .A(n453), .Y(n639) );
  AND2X1 U623 ( .A(n729), .B(n770), .Y(n467) );
  INVX1 U625 ( .A(n467), .Y(n640) );
  AND2X1 U627 ( .A(n690), .B(n773), .Y(n424) );
  INVX1 U629 ( .A(n424), .Y(n641) );
  AND2X1 U631 ( .A(n702), .B(n772), .Y(n437) );
  INVX1 U633 ( .A(n437), .Y(n642) );
  AND2X1 U635 ( .A(n718), .B(n771), .Y(n455) );
  INVX1 U637 ( .A(n455), .Y(n643) );
  AND2X1 U639 ( .A(n730), .B(n770), .Y(n468) );
  INVX1 U641 ( .A(n468), .Y(n644) );
  AND2X1 U643 ( .A(n691), .B(n773), .Y(n425) );
  INVX1 U645 ( .A(n425), .Y(n645) );
  AND2X1 U647 ( .A(n700), .B(n772), .Y(n435) );
  INVX1 U649 ( .A(n435), .Y(n646) );
  AND2X1 U651 ( .A(n719), .B(n771), .Y(n456) );
  INVX1 U653 ( .A(n456), .Y(n647) );
  AND2X1 U655 ( .A(n731), .B(n770), .Y(n469) );
  INVX1 U657 ( .A(n469), .Y(n648) );
  AND2X1 U659 ( .A(n701), .B(n772), .Y(n436) );
  INVX1 U661 ( .A(n436), .Y(n649) );
  AND2X1 U663 ( .A(n717), .B(n771), .Y(n454) );
  INVX1 U665 ( .A(n454), .Y(n650) );
  AND2X1 U667 ( .A(n734), .B(n770), .Y(n473) );
  INVX1 U669 ( .A(n473), .Y(n651) );
  AND2X1 U671 ( .A(n740), .B(n769), .Y(n479) );
  INVX1 U673 ( .A(n479), .Y(n652) );
  AND2X1 U675 ( .A(n692), .B(n773), .Y(n426) );
  INVX1 U677 ( .A(n426), .Y(n653) );
  AND2X1 U679 ( .A(n704), .B(n772), .Y(n440) );
  INVX1 U680 ( .A(n440), .Y(n654) );
  AND2X1 U683 ( .A(n721), .B(n771), .Y(n458) );
  INVX1 U686 ( .A(n458), .Y(n655) );
  AND2X1 U687 ( .A(n741), .B(n770), .Y(n480) );
  INVX1 U688 ( .A(n480), .Y(n656) );
  AND2X1 U689 ( .A(n703), .B(n772), .Y(n439) );
  INVX1 U690 ( .A(n439), .Y(n657) );
  AND2X1 U691 ( .A(n715), .B(n771), .Y(n452) );
  INVX1 U692 ( .A(n452), .Y(n658) );
  AND2X1 U693 ( .A(n733), .B(n770), .Y(n472) );
  INVX1 U694 ( .A(n472), .Y(n659) );
  AND2X1 U695 ( .A(n737), .B(n769), .Y(n476) );
  INVX1 U696 ( .A(n476), .Y(n660) );
  AND2X1 U697 ( .A(n743), .B(n773), .Y(n419) );
  INVX1 U698 ( .A(n419), .Y(n661) );
  AND2X1 U699 ( .A(n707), .B(n772), .Y(n443) );
  INVX1 U700 ( .A(n443), .Y(n662) );
  AND2X1 U701 ( .A(n722), .B(n771), .Y(n459) );
  INVX1 U702 ( .A(n459), .Y(n663) );
  AND2X1 U703 ( .A(n738), .B(n770), .Y(n477) );
  INVX1 U704 ( .A(n477), .Y(n664) );
  AND2X1 U705 ( .A(n744), .B(n773), .Y(n420) );
  INVX1 U706 ( .A(n420), .Y(n665) );
  AND2X1 U707 ( .A(n705), .B(n772), .Y(n441) );
  INVX1 U708 ( .A(n441), .Y(n666) );
  AND2X1 U709 ( .A(n720), .B(n771), .Y(n457) );
  INVX1 U710 ( .A(n457), .Y(n667) );
  AND2X1 U711 ( .A(n735), .B(n770), .Y(n474) );
  INVX1 U712 ( .A(n474), .Y(n668) );
  AND2X1 U713 ( .A(n739), .B(n769), .Y(n478) );
  INVX1 U714 ( .A(n478), .Y(n669) );
  AND2X1 U715 ( .A(n745), .B(n773), .Y(n421) );
  INVX1 U716 ( .A(n421), .Y(n670) );
  AND2X1 U717 ( .A(n732), .B(n771), .Y(n470) );
  INVX1 U718 ( .A(n470), .Y(n671) );
  AND2X1 U719 ( .A(n742), .B(n770), .Y(n481) );
  INVX1 U720 ( .A(n481), .Y(n672) );
  AND2X1 U721 ( .A(n746), .B(n773), .Y(n422) );
  INVX1 U722 ( .A(n422), .Y(n673) );
  AND2X1 U723 ( .A(n748), .B(n772), .Y(n438) );
  INVX1 U724 ( .A(n438), .Y(n674) );
  AND2X1 U725 ( .A(n708), .B(n772), .Y(n444) );
  INVX1 U726 ( .A(n444), .Y(n675) );
  AND2X1 U727 ( .A(n736), .B(n769), .Y(n475) );
  INVX1 U728 ( .A(n475), .Y(n676) );
  AND2X1 U729 ( .A(n747), .B(n773), .Y(n427) );
  INVX1 U730 ( .A(n427), .Y(n677) );
  AND2X1 U731 ( .A(n750), .B(n770), .Y(n460) );
  INVX1 U732 ( .A(n460), .Y(n678) );
  AND2X1 U733 ( .A(n752), .B(n771), .Y(n482) );
  INVX1 U734 ( .A(n482), .Y(n679) );
  BUFX2 U735 ( .A(evenBufferFull), .Y(n680) );
  AND2X1 U736 ( .A(n706), .B(n772), .Y(n442) );
  INVX1 U737 ( .A(n442), .Y(n681) );
  AND2X1 U738 ( .A(n749), .B(n771), .Y(n449) );
  INVX1 U739 ( .A(n449), .Y(n682) );
  AND2X1 U740 ( .A(n751), .B(n770), .Y(n471) );
  INVX1 U741 ( .A(n471), .Y(n683) );
  AND2X1 U742 ( .A(n776), .B(n773), .Y(n410) );
  INVX1 U743 ( .A(n410), .Y(n684) );
  AND2X1 U744 ( .A(readyOut), .B(n417), .Y(sendOut) );
  INVX1 U745 ( .A(sendOut), .Y(n685) );
  INVX1 U746 ( .A(n418), .Y(n686) );
  BUFX2 U747 ( .A(priorityRegEven), .Y(n687) );
  AND2X1 U748 ( .A(n776), .B(n775), .Y(n411) );
  INVX1 U749 ( .A(n411), .Y(n688) );
  BUFX2 U750 ( .A(evenBuffer[63]), .Y(n689) );
  BUFX2 U751 ( .A(evenBuffer[62]), .Y(n690) );
  BUFX2 U752 ( .A(evenBuffer[61]), .Y(n691) );
  BUFX2 U753 ( .A(evenBuffer[60]), .Y(n692) );
  BUFX2 U754 ( .A(evenBuffer[59]), .Y(n693) );
  BUFX2 U755 ( .A(evenBuffer[58]), .Y(n694) );
  BUFX2 U756 ( .A(evenBuffer[57]), .Y(n695) );
  BUFX2 U757 ( .A(evenBuffer[56]), .Y(n696) );
  BUFX2 U758 ( .A(evenBuffer[55]), .Y(n697) );
  BUFX2 U759 ( .A(evenBuffer[54]), .Y(n698) );
  BUFX2 U760 ( .A(evenBuffer[53]), .Y(n699) );
  BUFX2 U761 ( .A(evenBuffer[52]), .Y(n700) );
  BUFX2 U762 ( .A(evenBuffer[51]), .Y(n701) );
  BUFX2 U763 ( .A(evenBuffer[50]), .Y(n702) );
  BUFX2 U764 ( .A(evenBuffer[49]), .Y(n703) );
  BUFX2 U765 ( .A(evenBuffer[48]), .Y(n704) );
  BUFX2 U766 ( .A(evenBuffer[47]), .Y(n705) );
  BUFX2 U767 ( .A(evenBuffer[46]), .Y(n706) );
  BUFX2 U768 ( .A(evenBuffer[45]), .Y(n707) );
  BUFX2 U769 ( .A(evenBuffer[44]), .Y(n708) );
  BUFX2 U770 ( .A(evenBuffer[43]), .Y(n709) );
  BUFX2 U771 ( .A(evenBuffer[42]), .Y(n710) );
  BUFX2 U772 ( .A(evenBuffer[41]), .Y(n711) );
  BUFX2 U773 ( .A(evenBuffer[40]), .Y(n712) );
  BUFX2 U774 ( .A(evenBuffer[39]), .Y(n713) );
  BUFX2 U775 ( .A(evenBuffer[38]), .Y(n714) );
  BUFX2 U776 ( .A(evenBuffer[37]), .Y(n715) );
  BUFX2 U777 ( .A(evenBuffer[36]), .Y(n716) );
  BUFX2 U778 ( .A(evenBuffer[35]), .Y(n717) );
  BUFX2 U779 ( .A(evenBuffer[34]), .Y(n718) );
  BUFX2 U780 ( .A(evenBuffer[33]), .Y(n719) );
  BUFX2 U781 ( .A(evenBuffer[32]), .Y(n720) );
  BUFX2 U782 ( .A(evenBuffer[31]), .Y(n721) );
  BUFX2 U783 ( .A(evenBuffer[30]), .Y(n722) );
  BUFX2 U784 ( .A(evenBuffer[29]), .Y(n723) );
  BUFX2 U785 ( .A(evenBuffer[28]), .Y(n724) );
  BUFX2 U786 ( .A(evenBuffer[27]), .Y(n725) );
  BUFX2 U787 ( .A(evenBuffer[26]), .Y(n726) );
  BUFX2 U788 ( .A(evenBuffer[25]), .Y(n727) );
  BUFX2 U789 ( .A(evenBuffer[24]), .Y(n728) );
  BUFX2 U790 ( .A(evenBuffer[23]), .Y(n729) );
  BUFX2 U791 ( .A(evenBuffer[22]), .Y(n730) );
  BUFX2 U792 ( .A(evenBuffer[21]), .Y(n731) );
  BUFX2 U793 ( .A(evenBuffer[20]), .Y(n732) );
  BUFX2 U794 ( .A(evenBuffer[19]), .Y(n733) );
  BUFX2 U795 ( .A(evenBuffer[18]), .Y(n734) );
  BUFX2 U796 ( .A(evenBuffer[17]), .Y(n735) );
  BUFX2 U797 ( .A(evenBuffer[16]), .Y(n736) );
  BUFX2 U798 ( .A(evenBuffer[15]), .Y(n737) );
  BUFX2 U799 ( .A(evenBuffer[14]), .Y(n738) );
  BUFX2 U800 ( .A(evenBuffer[13]), .Y(n739) );
  BUFX2 U801 ( .A(evenBuffer[12]), .Y(n740) );
  BUFX2 U802 ( .A(evenBuffer[11]), .Y(n741) );
  BUFX2 U803 ( .A(evenBuffer[10]), .Y(n742) );
  BUFX2 U804 ( .A(evenBuffer[9]), .Y(n743) );
  BUFX2 U805 ( .A(evenBuffer[8]), .Y(n744) );
  BUFX2 U806 ( .A(evenBuffer[7]), .Y(n745) );
  BUFX2 U807 ( .A(evenBuffer[6]), .Y(n746) );
  BUFX2 U808 ( .A(evenBuffer[5]), .Y(n747) );
  BUFX2 U809 ( .A(evenBuffer[4]), .Y(n748) );
  BUFX2 U810 ( .A(evenBuffer[3]), .Y(n749) );
  BUFX2 U811 ( .A(evenBuffer[2]), .Y(n750) );
  BUFX2 U812 ( .A(evenBuffer[1]), .Y(n751) );
  BUFX2 U813 ( .A(evenBuffer[0]), .Y(n752) );
  AND2X1 U814 ( .A(n769), .B(n342), .Y(n409) );
  INVX1 U815 ( .A(n409), .Y(n753) );
  AND2X1 U816 ( .A(n272), .B(n774), .Y(n340) );
  INVX1 U817 ( .A(n340), .Y(n754) );
  BUFX2 U818 ( .A(priorityRegOdd), .Y(n755) );
  INVX1 U819 ( .A(n775), .Y(n770) );
  INVX1 U820 ( .A(n775), .Y(n771) );
  INVX1 U821 ( .A(n775), .Y(n769) );
  INVX1 U822 ( .A(n774), .Y(n768) );
  INVX1 U823 ( .A(n775), .Y(n767) );
  INVX1 U824 ( .A(n775), .Y(n765) );
  INVX1 U825 ( .A(n775), .Y(n766) );
  INVX1 U826 ( .A(n774), .Y(n773) );
  INVX1 U827 ( .A(n763), .Y(n774) );
  INVX1 U828 ( .A(n763), .Y(n775) );
  INVX1 U829 ( .A(n275), .Y(n761) );
  INVX1 U830 ( .A(n344), .Y(n760) );
  INVX1 U831 ( .A(n764), .Y(n763) );
  INVX1 U832 ( .A(n345), .Y(n759) );
  INVX1 U833 ( .A(n274), .Y(n762) );
  INVX1 U834 ( .A(n775), .Y(n772) );
  INVX1 U835 ( .A(polarity), .Y(n764) );
  INVX1 U836 ( .A(reset), .Y(n758) );
  INVX1 U837 ( .A(reset), .Y(n756) );
  INVX1 U838 ( .A(reset), .Y(n757) );
  AND2X1 U839 ( .A(n773), .B(n780), .Y(n487) );
  AND2X1 U840 ( .A(n777), .B(n775), .Y(n486) );
  INVX1 U841 ( .A(n412), .Y(n776) );
  INVX1 U842 ( .A(n755), .Y(n779) );
  INVX1 U843 ( .A(n741), .Y(n897) );
  INVX1 U844 ( .A(n740), .Y(n896) );
  INVX1 U845 ( .A(n739), .Y(n895) );
  INVX1 U846 ( .A(n738), .Y(n894) );
  INVX1 U847 ( .A(n737), .Y(n893) );
  INVX1 U848 ( .A(n736), .Y(n892) );
  INVX1 U849 ( .A(n735), .Y(n891) );
  INVX1 U850 ( .A(n734), .Y(n890) );
  INVX1 U851 ( .A(n733), .Y(n889) );
  INVX1 U852 ( .A(n732), .Y(n888) );
  INVX1 U853 ( .A(n731), .Y(n887) );
  INVX1 U854 ( .A(n730), .Y(n886) );
  INVX1 U855 ( .A(n729), .Y(n885) );
  INVX1 U856 ( .A(n727), .Y(n883) );
  INVX1 U857 ( .A(n728), .Y(n884) );
  INVX1 U858 ( .A(n726), .Y(n882) );
  INVX1 U859 ( .A(n725), .Y(n881) );
  INVX1 U860 ( .A(n724), .Y(n880) );
  INVX1 U861 ( .A(n723), .Y(n879) );
  INVX1 U862 ( .A(n722), .Y(n878) );
  INVX1 U863 ( .A(n721), .Y(n877) );
  INVX1 U864 ( .A(n720), .Y(n876) );
  INVX1 U865 ( .A(n719), .Y(n875) );
  INVX1 U866 ( .A(n718), .Y(n874) );
  INVX1 U867 ( .A(n717), .Y(n873) );
  INVX1 U868 ( .A(n716), .Y(n872) );
  INVX1 U869 ( .A(n715), .Y(n871) );
  INVX1 U870 ( .A(n714), .Y(n870) );
  INVX1 U871 ( .A(n713), .Y(n869) );
  INVX1 U872 ( .A(n712), .Y(n868) );
  INVX1 U873 ( .A(n711), .Y(n867) );
  INVX1 U874 ( .A(n710), .Y(n866) );
  INVX1 U875 ( .A(n709), .Y(n865) );
  INVX1 U876 ( .A(n708), .Y(n864) );
  INVX1 U877 ( .A(n707), .Y(n863) );
  INVX1 U878 ( .A(n706), .Y(n862) );
  INVX1 U879 ( .A(n705), .Y(n861) );
  INVX1 U880 ( .A(n704), .Y(n860) );
  INVX1 U881 ( .A(n703), .Y(n859) );
  INVX1 U882 ( .A(n702), .Y(n858) );
  INVX1 U883 ( .A(n701), .Y(n857) );
  INVX1 U884 ( .A(n700), .Y(n856) );
  INVX1 U885 ( .A(n699), .Y(n855) );
  INVX1 U886 ( .A(n698), .Y(n854) );
  INVX1 U887 ( .A(n697), .Y(n853) );
  INVX1 U888 ( .A(n696), .Y(n852) );
  INVX1 U889 ( .A(n695), .Y(n851) );
  INVX1 U890 ( .A(n694), .Y(n850) );
  INVX1 U891 ( .A(n693), .Y(n849) );
  INVX1 U892 ( .A(n692), .Y(n848) );
  INVX1 U893 ( .A(n691), .Y(n847) );
  INVX1 U894 ( .A(n690), .Y(n846) );
  INVX1 U895 ( .A(n752), .Y(n908) );
  INVX1 U896 ( .A(n751), .Y(n907) );
  INVX1 U897 ( .A(n750), .Y(n906) );
  INVX1 U898 ( .A(n749), .Y(n905) );
  INVX1 U899 ( .A(n748), .Y(n904) );
  INVX1 U900 ( .A(n747), .Y(n903) );
  INVX1 U901 ( .A(n746), .Y(n902) );
  INVX1 U902 ( .A(n745), .Y(n901) );
  INVX1 U903 ( .A(n744), .Y(n900) );
  INVX1 U904 ( .A(n743), .Y(n899) );
  INVX1 U905 ( .A(n742), .Y(n898) );
  INVX1 U906 ( .A(n689), .Y(n845) );
  INVX1 U907 ( .A(n687), .Y(n778) );
  INVX1 U908 ( .A(n680), .Y(n777) );
  INVX1 U909 ( .A(oddBufferFull), .Y(n780) );
  INVX1 U910 ( .A(oddBuffer[0]), .Y(n844) );
  INVX1 U911 ( .A(oddBuffer[1]), .Y(n843) );
  INVX1 U912 ( .A(oddBuffer[2]), .Y(n842) );
  INVX1 U913 ( .A(oddBuffer[3]), .Y(n841) );
  INVX1 U914 ( .A(oddBuffer[4]), .Y(n840) );
  INVX1 U915 ( .A(oddBuffer[5]), .Y(n839) );
  INVX1 U916 ( .A(oddBuffer[6]), .Y(n838) );
  INVX1 U917 ( .A(oddBuffer[7]), .Y(n837) );
  INVX1 U918 ( .A(oddBuffer[8]), .Y(n836) );
  INVX1 U919 ( .A(oddBuffer[9]), .Y(n835) );
  INVX1 U920 ( .A(oddBuffer[10]), .Y(n834) );
  INVX1 U921 ( .A(oddBuffer[11]), .Y(n833) );
  INVX1 U922 ( .A(oddBuffer[12]), .Y(n832) );
  INVX1 U923 ( .A(oddBuffer[13]), .Y(n831) );
  INVX1 U924 ( .A(oddBuffer[14]), .Y(n830) );
  INVX1 U925 ( .A(oddBuffer[15]), .Y(n829) );
  INVX1 U926 ( .A(oddBuffer[16]), .Y(n828) );
  INVX1 U927 ( .A(oddBuffer[17]), .Y(n827) );
  INVX1 U928 ( .A(oddBuffer[18]), .Y(n826) );
  INVX1 U929 ( .A(oddBuffer[19]), .Y(n825) );
  INVX1 U930 ( .A(oddBuffer[20]), .Y(n824) );
  INVX1 U931 ( .A(oddBuffer[21]), .Y(n823) );
  INVX1 U932 ( .A(oddBuffer[22]), .Y(n822) );
  INVX1 U933 ( .A(oddBuffer[23]), .Y(n821) );
  INVX1 U934 ( .A(oddBuffer[24]), .Y(n820) );
  INVX1 U935 ( .A(oddBuffer[25]), .Y(n819) );
  INVX1 U936 ( .A(oddBuffer[26]), .Y(n818) );
  INVX1 U937 ( .A(oddBuffer[27]), .Y(n817) );
  INVX1 U938 ( .A(oddBuffer[28]), .Y(n816) );
  INVX1 U939 ( .A(oddBuffer[29]), .Y(n815) );
  INVX1 U940 ( .A(oddBuffer[30]), .Y(n814) );
  INVX1 U941 ( .A(oddBuffer[31]), .Y(n813) );
  INVX1 U942 ( .A(oddBuffer[32]), .Y(n812) );
  INVX1 U943 ( .A(oddBuffer[33]), .Y(n811) );
  INVX1 U944 ( .A(oddBuffer[34]), .Y(n810) );
  INVX1 U945 ( .A(oddBuffer[35]), .Y(n809) );
  INVX1 U946 ( .A(oddBuffer[36]), .Y(n808) );
  INVX1 U947 ( .A(oddBuffer[37]), .Y(n807) );
  INVX1 U948 ( .A(oddBuffer[38]), .Y(n806) );
  INVX1 U949 ( .A(oddBuffer[39]), .Y(n805) );
  INVX1 U950 ( .A(oddBuffer[40]), .Y(n804) );
  INVX1 U951 ( .A(oddBuffer[41]), .Y(n803) );
  INVX1 U952 ( .A(oddBuffer[42]), .Y(n802) );
  INVX1 U953 ( .A(oddBuffer[43]), .Y(n801) );
  INVX1 U954 ( .A(oddBuffer[44]), .Y(n800) );
  INVX1 U955 ( .A(oddBuffer[45]), .Y(n799) );
  INVX1 U956 ( .A(oddBuffer[46]), .Y(n798) );
  INVX1 U957 ( .A(oddBuffer[47]), .Y(n797) );
  INVX1 U958 ( .A(oddBuffer[48]), .Y(n796) );
  INVX1 U959 ( .A(oddBuffer[49]), .Y(n795) );
  INVX1 U960 ( .A(oddBuffer[50]), .Y(n794) );
  INVX1 U961 ( .A(oddBuffer[51]), .Y(n793) );
  INVX1 U962 ( .A(oddBuffer[52]), .Y(n792) );
  INVX1 U963 ( .A(oddBuffer[53]), .Y(n791) );
  INVX1 U964 ( .A(oddBuffer[54]), .Y(n790) );
  INVX1 U965 ( .A(oddBuffer[55]), .Y(n789) );
  INVX1 U966 ( .A(oddBuffer[56]), .Y(n788) );
  INVX1 U967 ( .A(oddBuffer[57]), .Y(n787) );
  INVX1 U968 ( .A(oddBuffer[58]), .Y(n786) );
  INVX1 U969 ( .A(oddBuffer[59]), .Y(n785) );
  INVX1 U970 ( .A(oddBuffer[60]), .Y(n784) );
  INVX1 U971 ( .A(oddBuffer[61]), .Y(n783) );
  INVX1 U972 ( .A(oddBuffer[62]), .Y(n782) );
  INVX1 U973 ( .A(oddBuffer[63]), .Y(n781) );
endmodule


module outputBuffer_1 ( clk, reset, polarity, inputBufferRequest, dataIn0, 
        dataIn1, sendOut, readyOut, dataOut, InputBufferGrant );
  input [1:0] inputBufferRequest;
  input [63:0] dataIn0;
  input [63:0] dataIn1;
  output [63:0] dataOut;
  output [1:0] InputBufferGrant;
  input clk, reset, polarity, readyOut;
  output sendOut;
  wire   evenBufferFull, oddBufferFull, priorityRegEven, priorityRegOdd, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1191, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259;
  wire   [63:0] evenBuffer;
  wire   [63:0] oddBuffer;

  OAI21X1 U275 ( .A(n1259), .B(n845), .C(n130), .Y(n1041) );
  AOI22X1 U276 ( .A(dataIn1[63]), .B(n759), .C(dataIn0[63]), .D(n758), .Y(
        n1258) );
  OAI21X1 U277 ( .A(n1259), .B(n846), .C(n129), .Y(n1040) );
  AOI22X1 U278 ( .A(dataIn1[62]), .B(n759), .C(dataIn0[62]), .D(n758), .Y(
        n1255) );
  OAI21X1 U279 ( .A(n1259), .B(n847), .C(n128), .Y(n1039) );
  AOI22X1 U280 ( .A(dataIn1[61]), .B(n759), .C(dataIn0[61]), .D(n758), .Y(
        n1254) );
  OAI21X1 U281 ( .A(n1259), .B(n848), .C(n127), .Y(n1038) );
  AOI22X1 U282 ( .A(dataIn1[60]), .B(n759), .C(dataIn0[60]), .D(n758), .Y(
        n1253) );
  OAI21X1 U283 ( .A(n1259), .B(n849), .C(n126), .Y(n1037) );
  AOI22X1 U284 ( .A(dataIn1[59]), .B(n759), .C(dataIn0[59]), .D(n758), .Y(
        n1252) );
  OAI21X1 U285 ( .A(n1259), .B(n850), .C(n125), .Y(n1036) );
  AOI22X1 U286 ( .A(dataIn1[58]), .B(n759), .C(dataIn0[58]), .D(n758), .Y(
        n1251) );
  OAI21X1 U287 ( .A(n1259), .B(n851), .C(n124), .Y(n1035) );
  AOI22X1 U288 ( .A(dataIn1[57]), .B(n759), .C(dataIn0[57]), .D(n758), .Y(
        n1250) );
  OAI21X1 U289 ( .A(n1259), .B(n852), .C(n123), .Y(n1034) );
  AOI22X1 U290 ( .A(dataIn1[56]), .B(n759), .C(dataIn0[56]), .D(n758), .Y(
        n1249) );
  OAI21X1 U291 ( .A(n1259), .B(n853), .C(n122), .Y(n1033) );
  AOI22X1 U292 ( .A(dataIn1[55]), .B(n759), .C(dataIn0[55]), .D(n758), .Y(
        n1248) );
  OAI21X1 U293 ( .A(n1259), .B(n854), .C(n121), .Y(n1032) );
  AOI22X1 U294 ( .A(dataIn1[54]), .B(n759), .C(dataIn0[54]), .D(n758), .Y(
        n1247) );
  OAI21X1 U295 ( .A(n1259), .B(n855), .C(n120), .Y(n1031) );
  AOI22X1 U296 ( .A(dataIn1[53]), .B(n759), .C(dataIn0[53]), .D(n758), .Y(
        n1246) );
  OAI21X1 U297 ( .A(n1259), .B(n856), .C(n119), .Y(n1030) );
  AOI22X1 U298 ( .A(dataIn1[52]), .B(n759), .C(dataIn0[52]), .D(n758), .Y(
        n1245) );
  OAI21X1 U299 ( .A(n1259), .B(n857), .C(n118), .Y(n1029) );
  AOI22X1 U300 ( .A(dataIn1[51]), .B(n759), .C(dataIn0[51]), .D(n758), .Y(
        n1244) );
  OAI21X1 U301 ( .A(n1259), .B(n858), .C(n117), .Y(n1028) );
  AOI22X1 U302 ( .A(dataIn1[50]), .B(n759), .C(dataIn0[50]), .D(n758), .Y(
        n1243) );
  OAI21X1 U303 ( .A(n1259), .B(n859), .C(n116), .Y(n1027) );
  AOI22X1 U304 ( .A(dataIn1[49]), .B(n759), .C(dataIn0[49]), .D(n758), .Y(
        n1242) );
  OAI21X1 U305 ( .A(n1259), .B(n860), .C(n115), .Y(n1026) );
  AOI22X1 U306 ( .A(dataIn1[48]), .B(n759), .C(dataIn0[48]), .D(n758), .Y(
        n1241) );
  OAI21X1 U307 ( .A(n1259), .B(n861), .C(n114), .Y(n1025) );
  AOI22X1 U308 ( .A(dataIn1[47]), .B(n759), .C(dataIn0[47]), .D(n758), .Y(
        n1240) );
  OAI21X1 U309 ( .A(n1259), .B(n862), .C(n113), .Y(n1024) );
  AOI22X1 U310 ( .A(dataIn1[46]), .B(n759), .C(dataIn0[46]), .D(n758), .Y(
        n1239) );
  OAI21X1 U311 ( .A(n1259), .B(n863), .C(n112), .Y(n1023) );
  AOI22X1 U312 ( .A(dataIn1[45]), .B(n759), .C(dataIn0[45]), .D(n758), .Y(
        n1238) );
  OAI21X1 U313 ( .A(n1259), .B(n864), .C(n111), .Y(n1022) );
  AOI22X1 U314 ( .A(dataIn1[44]), .B(n759), .C(dataIn0[44]), .D(n758), .Y(
        n1237) );
  OAI21X1 U315 ( .A(n1259), .B(n865), .C(n110), .Y(n1021) );
  AOI22X1 U316 ( .A(dataIn1[43]), .B(n759), .C(dataIn0[43]), .D(n758), .Y(
        n1236) );
  OAI21X1 U317 ( .A(n1259), .B(n866), .C(n109), .Y(n1020) );
  AOI22X1 U318 ( .A(dataIn1[42]), .B(n759), .C(dataIn0[42]), .D(n758), .Y(
        n1235) );
  OAI21X1 U319 ( .A(n1259), .B(n867), .C(n108), .Y(n1019) );
  AOI22X1 U320 ( .A(dataIn1[41]), .B(n759), .C(dataIn0[41]), .D(n758), .Y(
        n1234) );
  OAI21X1 U321 ( .A(n1259), .B(n868), .C(n107), .Y(n1018) );
  AOI22X1 U322 ( .A(dataIn1[40]), .B(n759), .C(dataIn0[40]), .D(n758), .Y(
        n1233) );
  OAI21X1 U323 ( .A(n1259), .B(n869), .C(n106), .Y(n1017) );
  AOI22X1 U324 ( .A(dataIn1[39]), .B(n759), .C(dataIn0[39]), .D(n758), .Y(
        n1232) );
  OAI21X1 U325 ( .A(n1259), .B(n870), .C(n105), .Y(n1016) );
  AOI22X1 U326 ( .A(dataIn1[38]), .B(n759), .C(dataIn0[38]), .D(n758), .Y(
        n1231) );
  OAI21X1 U327 ( .A(n1259), .B(n871), .C(n104), .Y(n1015) );
  AOI22X1 U328 ( .A(dataIn1[37]), .B(n759), .C(dataIn0[37]), .D(n758), .Y(
        n1230) );
  OAI21X1 U329 ( .A(n1259), .B(n872), .C(n103), .Y(n1014) );
  AOI22X1 U330 ( .A(dataIn1[36]), .B(n759), .C(dataIn0[36]), .D(n758), .Y(
        n1229) );
  OAI21X1 U331 ( .A(n1259), .B(n873), .C(n102), .Y(n1013) );
  AOI22X1 U332 ( .A(dataIn1[35]), .B(n759), .C(dataIn0[35]), .D(n758), .Y(
        n1228) );
  OAI21X1 U333 ( .A(n1259), .B(n874), .C(n101), .Y(n1012) );
  AOI22X1 U334 ( .A(dataIn1[34]), .B(n759), .C(dataIn0[34]), .D(n758), .Y(
        n1227) );
  OAI21X1 U335 ( .A(n1259), .B(n875), .C(n100), .Y(n1011) );
  AOI22X1 U336 ( .A(dataIn1[33]), .B(n759), .C(dataIn0[33]), .D(n758), .Y(
        n1226) );
  OAI21X1 U337 ( .A(n1259), .B(n876), .C(n99), .Y(n1010) );
  AOI22X1 U338 ( .A(dataIn1[32]), .B(n759), .C(dataIn0[32]), .D(n758), .Y(
        n1225) );
  OAI21X1 U339 ( .A(n1259), .B(n877), .C(n98), .Y(n1009) );
  AOI22X1 U340 ( .A(dataIn1[31]), .B(n759), .C(dataIn0[31]), .D(n758), .Y(
        n1224) );
  OAI21X1 U341 ( .A(n1259), .B(n878), .C(n97), .Y(n1008) );
  AOI22X1 U342 ( .A(dataIn1[30]), .B(n759), .C(dataIn0[30]), .D(n758), .Y(
        n1223) );
  OAI21X1 U343 ( .A(n1259), .B(n879), .C(n96), .Y(n1007) );
  AOI22X1 U344 ( .A(dataIn1[29]), .B(n759), .C(dataIn0[29]), .D(n758), .Y(
        n1222) );
  OAI21X1 U345 ( .A(n1259), .B(n880), .C(n95), .Y(n1006) );
  AOI22X1 U346 ( .A(dataIn1[28]), .B(n759), .C(dataIn0[28]), .D(n758), .Y(
        n1221) );
  OAI21X1 U347 ( .A(n1259), .B(n881), .C(n94), .Y(n1005) );
  AOI22X1 U348 ( .A(dataIn1[27]), .B(n759), .C(dataIn0[27]), .D(n758), .Y(
        n1220) );
  OAI21X1 U349 ( .A(n1259), .B(n882), .C(n93), .Y(n1004) );
  AOI22X1 U350 ( .A(dataIn1[26]), .B(n759), .C(dataIn0[26]), .D(n758), .Y(
        n1219) );
  OAI21X1 U351 ( .A(n1259), .B(n883), .C(n92), .Y(n1003) );
  AOI22X1 U352 ( .A(dataIn1[25]), .B(n759), .C(dataIn0[25]), .D(n758), .Y(
        n1218) );
  OAI21X1 U353 ( .A(n1259), .B(n884), .C(n91), .Y(n1002) );
  AOI22X1 U354 ( .A(dataIn1[24]), .B(n759), .C(dataIn0[24]), .D(n758), .Y(
        n1217) );
  OAI21X1 U355 ( .A(n1259), .B(n885), .C(n90), .Y(n1001) );
  AOI22X1 U356 ( .A(dataIn1[23]), .B(n759), .C(dataIn0[23]), .D(n758), .Y(
        n1216) );
  OAI21X1 U357 ( .A(n1259), .B(n886), .C(n89), .Y(n1000) );
  AOI22X1 U358 ( .A(dataIn1[22]), .B(n759), .C(dataIn0[22]), .D(n758), .Y(
        n1215) );
  OAI21X1 U359 ( .A(n1259), .B(n887), .C(n88), .Y(n999) );
  AOI22X1 U360 ( .A(dataIn1[21]), .B(n759), .C(dataIn0[21]), .D(n758), .Y(
        n1214) );
  OAI21X1 U361 ( .A(n1259), .B(n888), .C(n87), .Y(n998) );
  AOI22X1 U362 ( .A(dataIn1[20]), .B(n759), .C(dataIn0[20]), .D(n758), .Y(
        n1213) );
  OAI21X1 U363 ( .A(n1259), .B(n889), .C(n86), .Y(n997) );
  AOI22X1 U364 ( .A(dataIn1[19]), .B(n759), .C(dataIn0[19]), .D(n758), .Y(
        n1212) );
  OAI21X1 U365 ( .A(n1259), .B(n890), .C(n85), .Y(n996) );
  AOI22X1 U366 ( .A(dataIn1[18]), .B(n759), .C(dataIn0[18]), .D(n758), .Y(
        n1211) );
  OAI21X1 U367 ( .A(n1259), .B(n891), .C(n84), .Y(n995) );
  AOI22X1 U368 ( .A(dataIn1[17]), .B(n759), .C(dataIn0[17]), .D(n758), .Y(
        n1210) );
  OAI21X1 U369 ( .A(n1259), .B(n892), .C(n83), .Y(n994) );
  AOI22X1 U370 ( .A(dataIn1[16]), .B(n759), .C(dataIn0[16]), .D(n758), .Y(
        n1209) );
  OAI21X1 U371 ( .A(n1259), .B(n893), .C(n82), .Y(n993) );
  AOI22X1 U372 ( .A(dataIn1[15]), .B(n759), .C(dataIn0[15]), .D(n758), .Y(
        n1208) );
  OAI21X1 U373 ( .A(n1259), .B(n894), .C(n81), .Y(n992) );
  AOI22X1 U374 ( .A(dataIn1[14]), .B(n759), .C(dataIn0[14]), .D(n758), .Y(
        n1207) );
  OAI21X1 U375 ( .A(n1259), .B(n895), .C(n80), .Y(n991) );
  AOI22X1 U376 ( .A(dataIn1[13]), .B(n759), .C(dataIn0[13]), .D(n758), .Y(
        n1206) );
  OAI21X1 U377 ( .A(n1259), .B(n896), .C(n79), .Y(n990) );
  AOI22X1 U378 ( .A(dataIn1[12]), .B(n759), .C(dataIn0[12]), .D(n758), .Y(
        n1205) );
  OAI21X1 U379 ( .A(n1259), .B(n897), .C(n78), .Y(n989) );
  AOI22X1 U380 ( .A(dataIn1[11]), .B(n759), .C(dataIn0[11]), .D(n758), .Y(
        n1204) );
  OAI21X1 U381 ( .A(n1259), .B(n898), .C(n77), .Y(n988) );
  AOI22X1 U382 ( .A(dataIn1[10]), .B(n759), .C(dataIn0[10]), .D(n758), .Y(
        n1203) );
  OAI21X1 U383 ( .A(n1259), .B(n899), .C(n76), .Y(n987) );
  AOI22X1 U384 ( .A(dataIn1[9]), .B(n759), .C(dataIn0[9]), .D(n758), .Y(n1202)
         );
  OAI21X1 U385 ( .A(n1259), .B(n900), .C(n75), .Y(n986) );
  AOI22X1 U386 ( .A(dataIn1[8]), .B(n759), .C(dataIn0[8]), .D(n758), .Y(n1201)
         );
  OAI21X1 U387 ( .A(n1259), .B(n901), .C(n74), .Y(n985) );
  AOI22X1 U388 ( .A(dataIn1[7]), .B(n759), .C(dataIn0[7]), .D(n758), .Y(n1200)
         );
  OAI21X1 U389 ( .A(n1259), .B(n902), .C(n73), .Y(n984) );
  AOI22X1 U390 ( .A(dataIn1[6]), .B(n759), .C(dataIn0[6]), .D(n758), .Y(n1199)
         );
  OAI21X1 U391 ( .A(n1259), .B(n903), .C(n72), .Y(n983) );
  AOI22X1 U392 ( .A(dataIn1[5]), .B(n759), .C(dataIn0[5]), .D(n758), .Y(n1198)
         );
  OAI21X1 U393 ( .A(n1259), .B(n904), .C(n71), .Y(n982) );
  AOI22X1 U394 ( .A(dataIn1[4]), .B(n759), .C(dataIn0[4]), .D(n758), .Y(n1197)
         );
  OAI21X1 U395 ( .A(n1259), .B(n905), .C(n70), .Y(n981) );
  AOI22X1 U396 ( .A(dataIn1[3]), .B(n759), .C(dataIn0[3]), .D(n758), .Y(n1196)
         );
  OAI21X1 U397 ( .A(n1259), .B(n906), .C(n69), .Y(n980) );
  AOI22X1 U398 ( .A(dataIn1[2]), .B(n759), .C(dataIn0[2]), .D(n758), .Y(n1195)
         );
  OAI21X1 U399 ( .A(n1259), .B(n907), .C(n68), .Y(n979) );
  AOI22X1 U400 ( .A(dataIn1[1]), .B(n759), .C(dataIn0[1]), .D(n758), .Y(n1194)
         );
  OAI21X1 U401 ( .A(n1259), .B(n908), .C(n67), .Y(n978) );
  AOI22X1 U402 ( .A(dataIn1[0]), .B(n759), .C(dataIn0[0]), .D(n758), .Y(n1193)
         );
  OAI21X1 U405 ( .A(n1189), .B(n781), .C(n66), .Y(n977) );
  AOI22X1 U406 ( .A(n757), .B(dataIn1[63]), .C(n756), .D(dataIn0[63]), .Y(
        n1188) );
  OAI21X1 U407 ( .A(n1189), .B(n782), .C(n65), .Y(n976) );
  AOI22X1 U408 ( .A(n757), .B(dataIn1[62]), .C(n756), .D(dataIn0[62]), .Y(
        n1185) );
  OAI21X1 U409 ( .A(n1189), .B(n783), .C(n64), .Y(n975) );
  AOI22X1 U410 ( .A(n757), .B(dataIn1[61]), .C(n756), .D(dataIn0[61]), .Y(
        n1184) );
  OAI21X1 U411 ( .A(n1189), .B(n784), .C(n63), .Y(n974) );
  AOI22X1 U412 ( .A(n757), .B(dataIn1[60]), .C(n756), .D(dataIn0[60]), .Y(
        n1183) );
  OAI21X1 U413 ( .A(n1189), .B(n785), .C(n62), .Y(n973) );
  AOI22X1 U414 ( .A(n757), .B(dataIn1[59]), .C(n756), .D(dataIn0[59]), .Y(
        n1182) );
  OAI21X1 U415 ( .A(n1189), .B(n786), .C(n61), .Y(n972) );
  AOI22X1 U416 ( .A(n757), .B(dataIn1[58]), .C(n756), .D(dataIn0[58]), .Y(
        n1181) );
  OAI21X1 U417 ( .A(n1189), .B(n787), .C(n60), .Y(n971) );
  AOI22X1 U418 ( .A(n757), .B(dataIn1[57]), .C(n756), .D(dataIn0[57]), .Y(
        n1180) );
  OAI21X1 U419 ( .A(n1189), .B(n788), .C(n59), .Y(n970) );
  AOI22X1 U420 ( .A(n757), .B(dataIn1[56]), .C(n756), .D(dataIn0[56]), .Y(
        n1179) );
  OAI21X1 U421 ( .A(n1189), .B(n789), .C(n58), .Y(n969) );
  AOI22X1 U422 ( .A(n757), .B(dataIn1[55]), .C(n756), .D(dataIn0[55]), .Y(
        n1178) );
  OAI21X1 U423 ( .A(n1189), .B(n790), .C(n57), .Y(n968) );
  AOI22X1 U424 ( .A(n757), .B(dataIn1[54]), .C(n756), .D(dataIn0[54]), .Y(
        n1177) );
  OAI21X1 U425 ( .A(n1189), .B(n791), .C(n56), .Y(n967) );
  AOI22X1 U426 ( .A(n757), .B(dataIn1[53]), .C(n756), .D(dataIn0[53]), .Y(
        n1176) );
  OAI21X1 U427 ( .A(n1189), .B(n792), .C(n55), .Y(n966) );
  AOI22X1 U428 ( .A(n757), .B(dataIn1[52]), .C(n756), .D(dataIn0[52]), .Y(
        n1175) );
  OAI21X1 U429 ( .A(n1189), .B(n793), .C(n54), .Y(n965) );
  AOI22X1 U430 ( .A(n757), .B(dataIn1[51]), .C(n756), .D(dataIn0[51]), .Y(
        n1174) );
  OAI21X1 U431 ( .A(n1189), .B(n794), .C(n53), .Y(n964) );
  AOI22X1 U432 ( .A(n757), .B(dataIn1[50]), .C(n756), .D(dataIn0[50]), .Y(
        n1173) );
  OAI21X1 U433 ( .A(n1189), .B(n795), .C(n52), .Y(n963) );
  AOI22X1 U434 ( .A(n757), .B(dataIn1[49]), .C(n756), .D(dataIn0[49]), .Y(
        n1172) );
  OAI21X1 U435 ( .A(n1189), .B(n796), .C(n51), .Y(n962) );
  AOI22X1 U436 ( .A(n757), .B(dataIn1[48]), .C(n756), .D(dataIn0[48]), .Y(
        n1171) );
  OAI21X1 U437 ( .A(n1189), .B(n797), .C(n50), .Y(n961) );
  AOI22X1 U438 ( .A(n757), .B(dataIn1[47]), .C(n756), .D(dataIn0[47]), .Y(
        n1170) );
  OAI21X1 U439 ( .A(n1189), .B(n798), .C(n49), .Y(n960) );
  AOI22X1 U440 ( .A(n757), .B(dataIn1[46]), .C(n756), .D(dataIn0[46]), .Y(
        n1169) );
  OAI21X1 U441 ( .A(n1189), .B(n799), .C(n48), .Y(n959) );
  AOI22X1 U442 ( .A(n757), .B(dataIn1[45]), .C(n756), .D(dataIn0[45]), .Y(
        n1168) );
  OAI21X1 U443 ( .A(n1189), .B(n800), .C(n47), .Y(n958) );
  AOI22X1 U444 ( .A(n757), .B(dataIn1[44]), .C(n756), .D(dataIn0[44]), .Y(
        n1167) );
  OAI21X1 U445 ( .A(n1189), .B(n801), .C(n46), .Y(n957) );
  AOI22X1 U446 ( .A(n757), .B(dataIn1[43]), .C(n756), .D(dataIn0[43]), .Y(
        n1166) );
  OAI21X1 U447 ( .A(n1189), .B(n802), .C(n45), .Y(n956) );
  AOI22X1 U448 ( .A(n757), .B(dataIn1[42]), .C(n756), .D(dataIn0[42]), .Y(
        n1165) );
  OAI21X1 U449 ( .A(n1189), .B(n803), .C(n44), .Y(n955) );
  AOI22X1 U450 ( .A(n757), .B(dataIn1[41]), .C(n756), .D(dataIn0[41]), .Y(
        n1164) );
  OAI21X1 U451 ( .A(n1189), .B(n804), .C(n43), .Y(n954) );
  AOI22X1 U452 ( .A(n757), .B(dataIn1[40]), .C(n756), .D(dataIn0[40]), .Y(
        n1163) );
  OAI21X1 U453 ( .A(n1189), .B(n805), .C(n42), .Y(n953) );
  AOI22X1 U454 ( .A(n757), .B(dataIn1[39]), .C(n756), .D(dataIn0[39]), .Y(
        n1162) );
  OAI21X1 U455 ( .A(n1189), .B(n806), .C(n41), .Y(n952) );
  AOI22X1 U456 ( .A(n757), .B(dataIn1[38]), .C(n756), .D(dataIn0[38]), .Y(
        n1161) );
  OAI21X1 U457 ( .A(n1189), .B(n807), .C(n40), .Y(n951) );
  AOI22X1 U458 ( .A(n757), .B(dataIn1[37]), .C(n756), .D(dataIn0[37]), .Y(
        n1160) );
  OAI21X1 U459 ( .A(n1189), .B(n808), .C(n39), .Y(n950) );
  AOI22X1 U460 ( .A(n757), .B(dataIn1[36]), .C(n756), .D(dataIn0[36]), .Y(
        n1159) );
  OAI21X1 U461 ( .A(n1189), .B(n809), .C(n38), .Y(n949) );
  AOI22X1 U462 ( .A(n757), .B(dataIn1[35]), .C(n756), .D(dataIn0[35]), .Y(
        n1158) );
  OAI21X1 U463 ( .A(n1189), .B(n810), .C(n37), .Y(n948) );
  AOI22X1 U464 ( .A(n757), .B(dataIn1[34]), .C(n756), .D(dataIn0[34]), .Y(
        n1157) );
  OAI21X1 U465 ( .A(n1189), .B(n811), .C(n36), .Y(n947) );
  AOI22X1 U466 ( .A(n757), .B(dataIn1[33]), .C(n756), .D(dataIn0[33]), .Y(
        n1156) );
  OAI21X1 U467 ( .A(n1189), .B(n812), .C(n35), .Y(n946) );
  AOI22X1 U468 ( .A(n757), .B(dataIn1[32]), .C(n756), .D(dataIn0[32]), .Y(
        n1155) );
  OAI21X1 U469 ( .A(n1189), .B(n813), .C(n34), .Y(n945) );
  AOI22X1 U470 ( .A(n757), .B(dataIn1[31]), .C(n756), .D(dataIn0[31]), .Y(
        n1154) );
  OAI21X1 U471 ( .A(n1189), .B(n814), .C(n33), .Y(n944) );
  AOI22X1 U472 ( .A(n757), .B(dataIn1[30]), .C(n756), .D(dataIn0[30]), .Y(
        n1153) );
  OAI21X1 U473 ( .A(n1189), .B(n815), .C(n32), .Y(n943) );
  AOI22X1 U474 ( .A(n757), .B(dataIn1[29]), .C(n756), .D(dataIn0[29]), .Y(
        n1152) );
  OAI21X1 U475 ( .A(n1189), .B(n816), .C(n31), .Y(n942) );
  AOI22X1 U476 ( .A(n757), .B(dataIn1[28]), .C(n756), .D(dataIn0[28]), .Y(
        n1151) );
  OAI21X1 U477 ( .A(n1189), .B(n817), .C(n30), .Y(n941) );
  AOI22X1 U478 ( .A(n757), .B(dataIn1[27]), .C(n756), .D(dataIn0[27]), .Y(
        n1150) );
  OAI21X1 U479 ( .A(n1189), .B(n818), .C(n29), .Y(n940) );
  AOI22X1 U480 ( .A(n757), .B(dataIn1[26]), .C(n756), .D(dataIn0[26]), .Y(
        n1149) );
  OAI21X1 U481 ( .A(n1189), .B(n819), .C(n28), .Y(n939) );
  AOI22X1 U482 ( .A(n757), .B(dataIn1[25]), .C(n756), .D(dataIn0[25]), .Y(
        n1148) );
  OAI21X1 U483 ( .A(n1189), .B(n820), .C(n27), .Y(n938) );
  AOI22X1 U484 ( .A(n757), .B(dataIn1[24]), .C(n756), .D(dataIn0[24]), .Y(
        n1147) );
  OAI21X1 U485 ( .A(n1189), .B(n821), .C(n26), .Y(n937) );
  AOI22X1 U486 ( .A(n757), .B(dataIn1[23]), .C(n756), .D(dataIn0[23]), .Y(
        n1146) );
  OAI21X1 U487 ( .A(n1189), .B(n822), .C(n25), .Y(n936) );
  AOI22X1 U488 ( .A(n757), .B(dataIn1[22]), .C(n756), .D(dataIn0[22]), .Y(
        n1145) );
  OAI21X1 U489 ( .A(n1189), .B(n823), .C(n24), .Y(n935) );
  AOI22X1 U490 ( .A(n757), .B(dataIn1[21]), .C(n756), .D(dataIn0[21]), .Y(
        n1144) );
  OAI21X1 U491 ( .A(n1189), .B(n824), .C(n23), .Y(n934) );
  AOI22X1 U492 ( .A(n757), .B(dataIn1[20]), .C(n756), .D(dataIn0[20]), .Y(
        n1143) );
  OAI21X1 U493 ( .A(n1189), .B(n825), .C(n22), .Y(n933) );
  AOI22X1 U494 ( .A(n757), .B(dataIn1[19]), .C(n756), .D(dataIn0[19]), .Y(
        n1142) );
  OAI21X1 U495 ( .A(n1189), .B(n826), .C(n21), .Y(n932) );
  AOI22X1 U496 ( .A(n757), .B(dataIn1[18]), .C(n756), .D(dataIn0[18]), .Y(
        n1141) );
  OAI21X1 U497 ( .A(n1189), .B(n827), .C(n20), .Y(n931) );
  AOI22X1 U498 ( .A(n757), .B(dataIn1[17]), .C(n756), .D(dataIn0[17]), .Y(
        n1140) );
  OAI21X1 U499 ( .A(n1189), .B(n828), .C(n19), .Y(n930) );
  AOI22X1 U500 ( .A(n757), .B(dataIn1[16]), .C(n756), .D(dataIn0[16]), .Y(
        n1139) );
  OAI21X1 U501 ( .A(n1189), .B(n829), .C(n18), .Y(n929) );
  AOI22X1 U502 ( .A(n757), .B(dataIn1[15]), .C(n756), .D(dataIn0[15]), .Y(
        n1138) );
  OAI21X1 U503 ( .A(n1189), .B(n830), .C(n17), .Y(n928) );
  AOI22X1 U504 ( .A(n757), .B(dataIn1[14]), .C(n756), .D(dataIn0[14]), .Y(
        n1137) );
  OAI21X1 U505 ( .A(n1189), .B(n831), .C(n16), .Y(n927) );
  AOI22X1 U506 ( .A(n757), .B(dataIn1[13]), .C(n756), .D(dataIn0[13]), .Y(
        n1136) );
  OAI21X1 U507 ( .A(n1189), .B(n832), .C(n15), .Y(n926) );
  AOI22X1 U508 ( .A(n757), .B(dataIn1[12]), .C(n756), .D(dataIn0[12]), .Y(
        n1135) );
  OAI21X1 U509 ( .A(n1189), .B(n833), .C(n14), .Y(n925) );
  AOI22X1 U510 ( .A(n757), .B(dataIn1[11]), .C(n756), .D(dataIn0[11]), .Y(
        n1134) );
  OAI21X1 U511 ( .A(n1189), .B(n834), .C(n13), .Y(n924) );
  AOI22X1 U512 ( .A(n757), .B(dataIn1[10]), .C(n756), .D(dataIn0[10]), .Y(
        n1133) );
  OAI21X1 U513 ( .A(n1189), .B(n835), .C(n12), .Y(n923) );
  AOI22X1 U514 ( .A(n757), .B(dataIn1[9]), .C(n756), .D(dataIn0[9]), .Y(n1132)
         );
  OAI21X1 U515 ( .A(n1189), .B(n836), .C(n11), .Y(n922) );
  AOI22X1 U516 ( .A(n757), .B(dataIn1[8]), .C(n756), .D(dataIn0[8]), .Y(n1131)
         );
  OAI21X1 U517 ( .A(n1189), .B(n837), .C(n10), .Y(n921) );
  AOI22X1 U518 ( .A(n757), .B(dataIn1[7]), .C(n756), .D(dataIn0[7]), .Y(n1130)
         );
  OAI21X1 U519 ( .A(n1189), .B(n838), .C(n9), .Y(n920) );
  AOI22X1 U520 ( .A(n757), .B(dataIn1[6]), .C(n756), .D(dataIn0[6]), .Y(n1129)
         );
  OAI21X1 U521 ( .A(n1189), .B(n839), .C(n8), .Y(n919) );
  AOI22X1 U522 ( .A(n757), .B(dataIn1[5]), .C(n756), .D(dataIn0[5]), .Y(n1128)
         );
  OAI21X1 U523 ( .A(n1189), .B(n840), .C(n7), .Y(n918) );
  AOI22X1 U524 ( .A(n757), .B(dataIn1[4]), .C(n756), .D(dataIn0[4]), .Y(n1127)
         );
  OAI21X1 U525 ( .A(n1189), .B(n841), .C(n6), .Y(n917) );
  AOI22X1 U526 ( .A(n757), .B(dataIn1[3]), .C(n756), .D(dataIn0[3]), .Y(n1126)
         );
  OAI21X1 U527 ( .A(n1189), .B(n842), .C(n5), .Y(n916) );
  AOI22X1 U528 ( .A(n757), .B(dataIn1[2]), .C(n756), .D(dataIn0[2]), .Y(n1125)
         );
  OAI21X1 U529 ( .A(n1189), .B(n843), .C(n4), .Y(n915) );
  AOI22X1 U530 ( .A(n757), .B(dataIn1[1]), .C(n756), .D(dataIn0[1]), .Y(n1124)
         );
  OAI21X1 U531 ( .A(n1189), .B(n844), .C(n3), .Y(n914) );
  AOI22X1 U532 ( .A(n757), .B(dataIn1[0]), .C(n756), .D(dataIn0[0]), .Y(n1123)
         );
  XNOR2X1 U535 ( .A(n755), .B(n684), .Y(n913) );
  XNOR2X1 U537 ( .A(n687), .B(n688), .Y(n912) );
  NAND3X1 U539 ( .A(inputBufferRequest[1]), .B(n149), .C(inputBufferRequest[0]), .Y(n1119) );
  OAI21X1 U540 ( .A(n780), .B(n1189), .C(n753), .Y(n911) );
  OAI21X1 U542 ( .A(n763), .B(n685), .C(n147), .Y(n1189) );
  OAI21X1 U544 ( .A(n777), .B(n1259), .C(n754), .Y(n910) );
  OAI21X1 U546 ( .A(n763), .B(n1118), .C(n146), .Y(n1259) );
  OAI21X1 U549 ( .A(n763), .B(n780), .C(n686), .Y(n1114) );
  OAI21X1 U552 ( .A(n763), .B(n835), .C(n661), .Y(dataOut[9]) );
  OAI21X1 U554 ( .A(n763), .B(n836), .C(n665), .Y(dataOut[8]) );
  OAI21X1 U556 ( .A(n763), .B(n837), .C(n670), .Y(dataOut[7]) );
  OAI21X1 U558 ( .A(n764), .B(n838), .C(n673), .Y(dataOut[6]) );
  OAI21X1 U560 ( .A(n764), .B(n781), .C(n637), .Y(dataOut[63]) );
  OAI21X1 U562 ( .A(n763), .B(n782), .C(n641), .Y(dataOut[62]) );
  OAI21X1 U564 ( .A(n764), .B(n783), .C(n645), .Y(dataOut[61]) );
  OAI21X1 U566 ( .A(n764), .B(n784), .C(n653), .Y(dataOut[60]) );
  OAI21X1 U568 ( .A(n764), .B(n839), .C(n677), .Y(dataOut[5]) );
  OAI21X1 U570 ( .A(n764), .B(n785), .C(n145), .Y(dataOut[59]) );
  OAI21X1 U572 ( .A(n765), .B(n786), .C(n144), .Y(dataOut[58]) );
  OAI21X1 U574 ( .A(n764), .B(n787), .C(n143), .Y(dataOut[57]) );
  OAI21X1 U576 ( .A(n765), .B(n788), .C(n142), .Y(dataOut[56]) );
  OAI21X1 U578 ( .A(n765), .B(n789), .C(n141), .Y(dataOut[55]) );
  OAI21X1 U580 ( .A(n763), .B(n790), .C(n634), .Y(dataOut[54]) );
  OAI21X1 U582 ( .A(n765), .B(n791), .C(n638), .Y(dataOut[53]) );
  OAI21X1 U584 ( .A(n765), .B(n792), .C(n646), .Y(dataOut[52]) );
  OAI21X1 U586 ( .A(n765), .B(n793), .C(n649), .Y(dataOut[51]) );
  OAI21X1 U588 ( .A(n766), .B(n794), .C(n642), .Y(dataOut[50]) );
  OAI21X1 U590 ( .A(n766), .B(n840), .C(n674), .Y(dataOut[4]) );
  OAI21X1 U592 ( .A(n765), .B(n795), .C(n657), .Y(dataOut[49]) );
  OAI21X1 U594 ( .A(n766), .B(n796), .C(n654), .Y(dataOut[48]) );
  OAI21X1 U596 ( .A(n766), .B(n797), .C(n666), .Y(dataOut[47]) );
  OAI21X1 U598 ( .A(n764), .B(n798), .C(n681), .Y(dataOut[46]) );
  OAI21X1 U600 ( .A(n767), .B(n799), .C(n662), .Y(dataOut[45]) );
  OAI21X1 U602 ( .A(n767), .B(n800), .C(n675), .Y(dataOut[44]) );
  OAI21X1 U604 ( .A(n765), .B(n801), .C(n140), .Y(dataOut[43]) );
  OAI21X1 U606 ( .A(n767), .B(n802), .C(n139), .Y(dataOut[42]) );
  OAI21X1 U608 ( .A(n767), .B(n803), .C(n138), .Y(dataOut[41]) );
  OAI21X1 U610 ( .A(n766), .B(n804), .C(n137), .Y(dataOut[40]) );
  OAI21X1 U612 ( .A(n767), .B(n841), .C(n682), .Y(dataOut[3]) );
  OAI21X1 U614 ( .A(n767), .B(n805), .C(n136), .Y(dataOut[39]) );
  OAI21X1 U616 ( .A(n765), .B(n806), .C(n635), .Y(dataOut[38]) );
  OAI21X1 U618 ( .A(n767), .B(n807), .C(n658), .Y(dataOut[37]) );
  OAI21X1 U620 ( .A(n768), .B(n808), .C(n639), .Y(dataOut[36]) );
  OAI21X1 U622 ( .A(n766), .B(n809), .C(n650), .Y(dataOut[35]) );
  OAI21X1 U624 ( .A(n768), .B(n810), .C(n643), .Y(dataOut[34]) );
  OAI21X1 U626 ( .A(n768), .B(n811), .C(n647), .Y(dataOut[33]) );
  OAI21X1 U628 ( .A(n767), .B(n812), .C(n667), .Y(dataOut[32]) );
  OAI21X1 U630 ( .A(n768), .B(n813), .C(n655), .Y(dataOut[31]) );
  OAI21X1 U632 ( .A(n768), .B(n814), .C(n663), .Y(dataOut[30]) );
  OAI21X1 U634 ( .A(n766), .B(n842), .C(n678), .Y(dataOut[2]) );
  OAI21X1 U636 ( .A(n767), .B(n815), .C(n135), .Y(dataOut[29]) );
  OAI21X1 U638 ( .A(n768), .B(n816), .C(n134), .Y(dataOut[28]) );
  OAI21X1 U640 ( .A(n768), .B(n817), .C(n133), .Y(dataOut[27]) );
  OAI21X1 U642 ( .A(n766), .B(n818), .C(n132), .Y(dataOut[26]) );
  OAI21X1 U644 ( .A(n767), .B(n819), .C(n131), .Y(dataOut[25]) );
  OAI21X1 U646 ( .A(n767), .B(n820), .C(n636), .Y(dataOut[24]) );
  OAI21X1 U648 ( .A(n766), .B(n821), .C(n640), .Y(dataOut[23]) );
  OAI21X1 U650 ( .A(n767), .B(n822), .C(n644), .Y(dataOut[22]) );
  OAI21X1 U652 ( .A(n766), .B(n823), .C(n648), .Y(dataOut[21]) );
  OAI21X1 U654 ( .A(n765), .B(n824), .C(n671), .Y(dataOut[20]) );
  OAI21X1 U656 ( .A(n766), .B(n843), .C(n683), .Y(dataOut[1]) );
  OAI21X1 U658 ( .A(n766), .B(n825), .C(n659), .Y(dataOut[19]) );
  OAI21X1 U660 ( .A(n764), .B(n826), .C(n651), .Y(dataOut[18]) );
  OAI21X1 U662 ( .A(n765), .B(n827), .C(n668), .Y(dataOut[17]) );
  OAI21X1 U664 ( .A(n765), .B(n828), .C(n676), .Y(dataOut[16]) );
  OAI21X1 U666 ( .A(n764), .B(n829), .C(n660), .Y(dataOut[15]) );
  OAI21X1 U668 ( .A(n764), .B(n830), .C(n664), .Y(dataOut[14]) );
  OAI21X1 U670 ( .A(n764), .B(n831), .C(n669), .Y(dataOut[13]) );
  OAI21X1 U672 ( .A(n763), .B(n832), .C(n652), .Y(dataOut[12]) );
  OAI21X1 U674 ( .A(n763), .B(n833), .C(n656), .Y(dataOut[11]) );
  OAI21X1 U676 ( .A(n763), .B(n834), .C(n672), .Y(dataOut[10]) );
  OAI21X1 U678 ( .A(n763), .B(n844), .C(n679), .Y(dataOut[0]) );
  OAI21X1 U681 ( .A(inputBufferRequest[0]), .B(n148), .C(n2), .Y(n1048) );
  AOI22X1 U682 ( .A(n687), .B(n1045), .C(n755), .D(n1044), .Y(n1046) );
  OAI21X1 U684 ( .A(inputBufferRequest[1]), .B(n148), .C(n1), .Y(n1043) );
  AOI22X1 U685 ( .A(n1045), .B(n778), .C(n1044), .D(n779), .Y(n1042) );
  DFFSR priorityRegOdd_reg ( .D(n913), .CLK(clk), .R(n909), .S(1'b1), .Q(
        priorityRegOdd) );
  DFFSR priorityRegEven_reg ( .D(n912), .CLK(clk), .R(n909), .S(1'b1), .Q(
        priorityRegEven) );
  DFFSR oddBufferFull_reg ( .D(n911), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBufferFull) );
  DFFSR evenBufferFull_reg ( .D(n910), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBufferFull) );
  DFFSR oddBuffer_reg_63_ ( .D(n977), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[63]) );
  DFFSR oddBuffer_reg_62_ ( .D(n976), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[62]) );
  DFFSR oddBuffer_reg_61_ ( .D(n975), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[61]) );
  DFFSR oddBuffer_reg_60_ ( .D(n974), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[60]) );
  DFFSR oddBuffer_reg_59_ ( .D(n973), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[59]) );
  DFFSR oddBuffer_reg_58_ ( .D(n972), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[58]) );
  DFFSR oddBuffer_reg_57_ ( .D(n971), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[57]) );
  DFFSR oddBuffer_reg_56_ ( .D(n970), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[56]) );
  DFFSR oddBuffer_reg_55_ ( .D(n969), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[55]) );
  DFFSR oddBuffer_reg_54_ ( .D(n968), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[54]) );
  DFFSR oddBuffer_reg_53_ ( .D(n967), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[53]) );
  DFFSR oddBuffer_reg_52_ ( .D(n966), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[52]) );
  DFFSR oddBuffer_reg_10_ ( .D(n924), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[10]) );
  DFFSR oddBuffer_reg_8_ ( .D(n922), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[8]) );
  DFFSR oddBuffer_reg_7_ ( .D(n921), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[7]) );
  DFFSR oddBuffer_reg_6_ ( .D(n920), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[6]) );
  DFFSR oddBuffer_reg_5_ ( .D(n919), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[5]) );
  DFFSR oddBuffer_reg_4_ ( .D(n918), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[4]) );
  DFFSR oddBuffer_reg_3_ ( .D(n917), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[3]) );
  DFFSR oddBuffer_reg_2_ ( .D(n916), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[2]) );
  DFFSR oddBuffer_reg_1_ ( .D(n915), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[1]) );
  DFFSR oddBuffer_reg_0_ ( .D(n914), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[0]) );
  DFFSR oddBuffer_reg_9_ ( .D(n923), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[9]) );
  DFFSR oddBuffer_reg_25_ ( .D(n939), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[25]) );
  DFFSR oddBuffer_reg_23_ ( .D(n937), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[23]) );
  DFFSR oddBuffer_reg_22_ ( .D(n936), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[22]) );
  DFFSR oddBuffer_reg_21_ ( .D(n935), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[21]) );
  DFFSR oddBuffer_reg_20_ ( .D(n934), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[20]) );
  DFFSR oddBuffer_reg_19_ ( .D(n933), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[19]) );
  DFFSR oddBuffer_reg_18_ ( .D(n932), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[18]) );
  DFFSR oddBuffer_reg_17_ ( .D(n931), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[17]) );
  DFFSR oddBuffer_reg_16_ ( .D(n930), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[16]) );
  DFFSR oddBuffer_reg_15_ ( .D(n929), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[15]) );
  DFFSR oddBuffer_reg_14_ ( .D(n928), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[14]) );
  DFFSR oddBuffer_reg_13_ ( .D(n927), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[13]) );
  DFFSR oddBuffer_reg_12_ ( .D(n926), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[12]) );
  DFFSR oddBuffer_reg_11_ ( .D(n925), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[11]) );
  DFFSR oddBuffer_reg_24_ ( .D(n938), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[24]) );
  DFFSR evenBuffer_reg_63_ ( .D(n1041), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[63]) );
  DFFSR evenBuffer_reg_62_ ( .D(n1040), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[62]) );
  DFFSR evenBuffer_reg_61_ ( .D(n1039), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[61]) );
  DFFSR evenBuffer_reg_60_ ( .D(n1038), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[60]) );
  DFFSR evenBuffer_reg_59_ ( .D(n1037), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[59]) );
  DFFSR evenBuffer_reg_58_ ( .D(n1036), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[58]) );
  DFFSR evenBuffer_reg_57_ ( .D(n1035), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[57]) );
  DFFSR evenBuffer_reg_56_ ( .D(n1034), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[56]) );
  DFFSR evenBuffer_reg_55_ ( .D(n1033), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[55]) );
  DFFSR evenBuffer_reg_54_ ( .D(n1032), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[54]) );
  DFFSR evenBuffer_reg_53_ ( .D(n1031), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[53]) );
  DFFSR evenBuffer_reg_52_ ( .D(n1030), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[52]) );
  DFFSR oddBuffer_reg_47_ ( .D(n961), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[47]) );
  DFFSR oddBuffer_reg_46_ ( .D(n960), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[46]) );
  DFFSR oddBuffer_reg_45_ ( .D(n959), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[45]) );
  DFFSR oddBuffer_reg_44_ ( .D(n958), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[44]) );
  DFFSR oddBuffer_reg_43_ ( .D(n957), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[43]) );
  DFFSR oddBuffer_reg_42_ ( .D(n956), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[42]) );
  DFFSR oddBuffer_reg_41_ ( .D(n955), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[41]) );
  DFFSR oddBuffer_reg_40_ ( .D(n954), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[40]) );
  DFFSR oddBuffer_reg_39_ ( .D(n953), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[39]) );
  DFFSR oddBuffer_reg_38_ ( .D(n952), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[38]) );
  DFFSR oddBuffer_reg_37_ ( .D(n951), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[37]) );
  DFFSR oddBuffer_reg_36_ ( .D(n950), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[36]) );
  DFFSR oddBuffer_reg_35_ ( .D(n949), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[35]) );
  DFFSR oddBuffer_reg_34_ ( .D(n948), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[34]) );
  DFFSR oddBuffer_reg_33_ ( .D(n947), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[33]) );
  DFFSR oddBuffer_reg_32_ ( .D(n946), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[32]) );
  DFFSR oddBuffer_reg_31_ ( .D(n945), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[31]) );
  DFFSR oddBuffer_reg_30_ ( .D(n944), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[30]) );
  DFFSR oddBuffer_reg_29_ ( .D(n943), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[29]) );
  DFFSR oddBuffer_reg_26_ ( .D(n940), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[26]) );
  DFFSR oddBuffer_reg_28_ ( .D(n942), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[28]) );
  DFFSR oddBuffer_reg_27_ ( .D(n941), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[27]) );
  DFFSR oddBuffer_reg_51_ ( .D(n965), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[51]) );
  DFFSR oddBuffer_reg_50_ ( .D(n964), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[50]) );
  DFFSR oddBuffer_reg_49_ ( .D(n963), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[49]) );
  DFFSR oddBuffer_reg_48_ ( .D(n962), .CLK(clk), .R(n909), .S(1'b1), .Q(
        oddBuffer[48]) );
  DFFSR evenBuffer_reg_10_ ( .D(n988), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[10]) );
  DFFSR evenBuffer_reg_9_ ( .D(n987), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[9]) );
  DFFSR evenBuffer_reg_8_ ( .D(n986), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[8]) );
  DFFSR evenBuffer_reg_7_ ( .D(n985), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[7]) );
  DFFSR evenBuffer_reg_6_ ( .D(n984), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[6]) );
  DFFSR evenBuffer_reg_5_ ( .D(n983), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[5]) );
  DFFSR evenBuffer_reg_4_ ( .D(n982), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[4]) );
  DFFSR evenBuffer_reg_3_ ( .D(n981), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[3]) );
  DFFSR evenBuffer_reg_2_ ( .D(n980), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[2]) );
  DFFSR evenBuffer_reg_1_ ( .D(n979), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[1]) );
  DFFSR evenBuffer_reg_0_ ( .D(n978), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[0]) );
  DFFSR evenBuffer_reg_25_ ( .D(n1003), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[25]) );
  DFFSR evenBuffer_reg_24_ ( .D(n1002), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[24]) );
  DFFSR evenBuffer_reg_23_ ( .D(n1001), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[23]) );
  DFFSR evenBuffer_reg_22_ ( .D(n1000), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[22]) );
  DFFSR evenBuffer_reg_21_ ( .D(n999), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[21]) );
  DFFSR evenBuffer_reg_20_ ( .D(n998), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[20]) );
  DFFSR evenBuffer_reg_19_ ( .D(n997), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[19]) );
  DFFSR evenBuffer_reg_18_ ( .D(n996), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[18]) );
  DFFSR evenBuffer_reg_17_ ( .D(n995), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[17]) );
  DFFSR evenBuffer_reg_16_ ( .D(n994), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[16]) );
  DFFSR evenBuffer_reg_15_ ( .D(n993), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[15]) );
  DFFSR evenBuffer_reg_14_ ( .D(n992), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[14]) );
  DFFSR evenBuffer_reg_13_ ( .D(n991), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[13]) );
  DFFSR evenBuffer_reg_12_ ( .D(n990), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[12]) );
  DFFSR evenBuffer_reg_11_ ( .D(n989), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[11]) );
  DFFSR evenBuffer_reg_51_ ( .D(n1029), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[51]) );
  DFFSR evenBuffer_reg_50_ ( .D(n1028), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[50]) );
  DFFSR evenBuffer_reg_49_ ( .D(n1027), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[49]) );
  DFFSR evenBuffer_reg_48_ ( .D(n1026), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[48]) );
  DFFSR evenBuffer_reg_47_ ( .D(n1025), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[47]) );
  DFFSR evenBuffer_reg_46_ ( .D(n1024), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[46]) );
  DFFSR evenBuffer_reg_45_ ( .D(n1023), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[45]) );
  DFFSR evenBuffer_reg_44_ ( .D(n1022), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[44]) );
  DFFSR evenBuffer_reg_43_ ( .D(n1021), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[43]) );
  DFFSR evenBuffer_reg_42_ ( .D(n1020), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[42]) );
  DFFSR evenBuffer_reg_41_ ( .D(n1019), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[41]) );
  DFFSR evenBuffer_reg_40_ ( .D(n1018), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[40]) );
  DFFSR evenBuffer_reg_39_ ( .D(n1017), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[39]) );
  DFFSR evenBuffer_reg_38_ ( .D(n1016), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[38]) );
  DFFSR evenBuffer_reg_37_ ( .D(n1015), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[37]) );
  DFFSR evenBuffer_reg_36_ ( .D(n1014), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[36]) );
  DFFSR evenBuffer_reg_35_ ( .D(n1013), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[35]) );
  DFFSR evenBuffer_reg_34_ ( .D(n1012), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[34]) );
  DFFSR evenBuffer_reg_33_ ( .D(n1011), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[33]) );
  DFFSR evenBuffer_reg_32_ ( .D(n1010), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[32]) );
  DFFSR evenBuffer_reg_31_ ( .D(n1009), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[31]) );
  DFFSR evenBuffer_reg_30_ ( .D(n1008), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[30]) );
  DFFSR evenBuffer_reg_29_ ( .D(n1007), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[29]) );
  DFFSR evenBuffer_reg_28_ ( .D(n1006), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[28]) );
  DFFSR evenBuffer_reg_27_ ( .D(n1005), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[27]) );
  DFFSR evenBuffer_reg_26_ ( .D(n1004), .CLK(clk), .R(n909), .S(1'b1), .Q(
        evenBuffer[26]) );
  AND2X1 U2 ( .A(n768), .B(n680), .Y(n1113) );
  AND2X1 U3 ( .A(inputBufferRequest[1]), .B(n1048), .Y(InputBufferGrant[1]) );
  AND2X1 U4 ( .A(inputBufferRequest[0]), .B(n1043), .Y(InputBufferGrant[0]) );
  OR2X1 U5 ( .A(n753), .B(n151), .Y(n1187) );
  OR2X1 U6 ( .A(n753), .B(n150), .Y(n1186) );
  OR2X1 U7 ( .A(n754), .B(n151), .Y(n1257) );
  OR2X1 U8 ( .A(n150), .B(n754), .Y(n1256) );
  BUFX2 U9 ( .A(n1042), .Y(n1) );
  BUFX2 U10 ( .A(n1046), .Y(n2) );
  BUFX2 U11 ( .A(n1123), .Y(n3) );
  BUFX2 U12 ( .A(n1124), .Y(n4) );
  BUFX2 U13 ( .A(n1125), .Y(n5) );
  BUFX2 U14 ( .A(n1126), .Y(n6) );
  BUFX2 U15 ( .A(n1127), .Y(n7) );
  BUFX2 U16 ( .A(n1128), .Y(n8) );
  BUFX2 U17 ( .A(n1129), .Y(n9) );
  BUFX2 U18 ( .A(n1130), .Y(n10) );
  BUFX2 U19 ( .A(n1131), .Y(n11) );
  BUFX2 U20 ( .A(n1132), .Y(n12) );
  BUFX2 U21 ( .A(n1133), .Y(n13) );
  BUFX2 U22 ( .A(n1134), .Y(n14) );
  BUFX2 U23 ( .A(n1135), .Y(n15) );
  BUFX2 U24 ( .A(n1136), .Y(n16) );
  BUFX2 U25 ( .A(n1137), .Y(n17) );
  BUFX2 U26 ( .A(n1138), .Y(n18) );
  BUFX2 U27 ( .A(n1139), .Y(n19) );
  BUFX2 U28 ( .A(n1140), .Y(n20) );
  BUFX2 U29 ( .A(n1141), .Y(n21) );
  BUFX2 U30 ( .A(n1142), .Y(n22) );
  BUFX2 U31 ( .A(n1143), .Y(n23) );
  BUFX2 U32 ( .A(n1144), .Y(n24) );
  BUFX2 U33 ( .A(n1145), .Y(n25) );
  BUFX2 U34 ( .A(n1146), .Y(n26) );
  BUFX2 U35 ( .A(n1147), .Y(n27) );
  BUFX2 U36 ( .A(n1148), .Y(n28) );
  BUFX2 U37 ( .A(n1149), .Y(n29) );
  BUFX2 U38 ( .A(n1150), .Y(n30) );
  BUFX2 U39 ( .A(n1151), .Y(n31) );
  BUFX2 U40 ( .A(n1152), .Y(n32) );
  BUFX2 U41 ( .A(n1153), .Y(n33) );
  BUFX2 U42 ( .A(n1154), .Y(n34) );
  BUFX2 U43 ( .A(n1155), .Y(n35) );
  BUFX2 U44 ( .A(n1156), .Y(n36) );
  BUFX2 U45 ( .A(n1157), .Y(n37) );
  BUFX2 U46 ( .A(n1158), .Y(n38) );
  BUFX2 U47 ( .A(n1159), .Y(n39) );
  BUFX2 U48 ( .A(n1160), .Y(n40) );
  BUFX2 U49 ( .A(n1161), .Y(n41) );
  BUFX2 U50 ( .A(n1162), .Y(n42) );
  BUFX2 U51 ( .A(n1163), .Y(n43) );
  BUFX2 U52 ( .A(n1164), .Y(n44) );
  BUFX2 U53 ( .A(n1165), .Y(n45) );
  BUFX2 U54 ( .A(n1166), .Y(n46) );
  BUFX2 U55 ( .A(n1167), .Y(n47) );
  BUFX2 U56 ( .A(n1168), .Y(n48) );
  BUFX2 U57 ( .A(n1169), .Y(n49) );
  BUFX2 U58 ( .A(n1170), .Y(n50) );
  BUFX2 U59 ( .A(n1171), .Y(n51) );
  BUFX2 U60 ( .A(n1172), .Y(n52) );
  BUFX2 U61 ( .A(n1173), .Y(n53) );
  BUFX2 U62 ( .A(n1174), .Y(n54) );
  BUFX2 U63 ( .A(n1175), .Y(n55) );
  BUFX2 U64 ( .A(n1176), .Y(n56) );
  BUFX2 U65 ( .A(n1177), .Y(n57) );
  BUFX2 U66 ( .A(n1178), .Y(n58) );
  BUFX2 U67 ( .A(n1179), .Y(n59) );
  BUFX2 U68 ( .A(n1180), .Y(n60) );
  BUFX2 U69 ( .A(n1181), .Y(n61) );
  BUFX2 U70 ( .A(n1182), .Y(n62) );
  BUFX2 U71 ( .A(n1183), .Y(n63) );
  BUFX2 U72 ( .A(n1184), .Y(n64) );
  BUFX2 U73 ( .A(n1185), .Y(n65) );
  BUFX2 U74 ( .A(n1188), .Y(n66) );
  BUFX2 U75 ( .A(n1193), .Y(n67) );
  BUFX2 U76 ( .A(n1194), .Y(n68) );
  BUFX2 U77 ( .A(n1195), .Y(n69) );
  BUFX2 U78 ( .A(n1196), .Y(n70) );
  BUFX2 U79 ( .A(n1197), .Y(n71) );
  BUFX2 U80 ( .A(n1198), .Y(n72) );
  BUFX2 U81 ( .A(n1199), .Y(n73) );
  BUFX2 U82 ( .A(n1200), .Y(n74) );
  BUFX2 U83 ( .A(n1201), .Y(n75) );
  BUFX2 U84 ( .A(n1202), .Y(n76) );
  BUFX2 U85 ( .A(n1203), .Y(n77) );
  BUFX2 U86 ( .A(n1204), .Y(n78) );
  BUFX2 U87 ( .A(n1205), .Y(n79) );
  BUFX2 U88 ( .A(n1206), .Y(n80) );
  BUFX2 U89 ( .A(n1207), .Y(n81) );
  BUFX2 U90 ( .A(n1208), .Y(n82) );
  BUFX2 U91 ( .A(n1209), .Y(n83) );
  BUFX2 U92 ( .A(n1210), .Y(n84) );
  BUFX2 U93 ( .A(n1211), .Y(n85) );
  BUFX2 U94 ( .A(n1212), .Y(n86) );
  BUFX2 U95 ( .A(n1213), .Y(n87) );
  BUFX2 U96 ( .A(n1214), .Y(n88) );
  BUFX2 U97 ( .A(n1215), .Y(n89) );
  BUFX2 U98 ( .A(n1216), .Y(n90) );
  BUFX2 U99 ( .A(n1217), .Y(n91) );
  BUFX2 U100 ( .A(n1218), .Y(n92) );
  BUFX2 U101 ( .A(n1219), .Y(n93) );
  BUFX2 U102 ( .A(n1220), .Y(n94) );
  BUFX2 U103 ( .A(n1221), .Y(n95) );
  BUFX2 U104 ( .A(n1222), .Y(n96) );
  BUFX2 U105 ( .A(n1223), .Y(n97) );
  BUFX2 U106 ( .A(n1224), .Y(n98) );
  BUFX2 U107 ( .A(n1225), .Y(n99) );
  BUFX2 U108 ( .A(n1226), .Y(n100) );
  BUFX2 U109 ( .A(n1227), .Y(n101) );
  BUFX2 U110 ( .A(n1228), .Y(n102) );
  BUFX2 U111 ( .A(n1229), .Y(n103) );
  BUFX2 U112 ( .A(n1230), .Y(n104) );
  BUFX2 U113 ( .A(n1231), .Y(n105) );
  BUFX2 U114 ( .A(n1232), .Y(n106) );
  BUFX2 U115 ( .A(n1233), .Y(n107) );
  BUFX2 U116 ( .A(n1234), .Y(n108) );
  BUFX2 U117 ( .A(n1235), .Y(n109) );
  BUFX2 U118 ( .A(n1236), .Y(n110) );
  BUFX2 U119 ( .A(n1237), .Y(n111) );
  BUFX2 U120 ( .A(n1238), .Y(n112) );
  BUFX2 U121 ( .A(n1239), .Y(n113) );
  BUFX2 U122 ( .A(n1240), .Y(n114) );
  BUFX2 U123 ( .A(n1241), .Y(n115) );
  BUFX2 U124 ( .A(n1242), .Y(n116) );
  BUFX2 U125 ( .A(n1243), .Y(n117) );
  BUFX2 U126 ( .A(n1244), .Y(n118) );
  BUFX2 U127 ( .A(n1245), .Y(n119) );
  BUFX2 U128 ( .A(n1246), .Y(n120) );
  BUFX2 U129 ( .A(n1247), .Y(n121) );
  BUFX2 U130 ( .A(n1248), .Y(n122) );
  BUFX2 U131 ( .A(n1249), .Y(n123) );
  BUFX2 U132 ( .A(n1250), .Y(n124) );
  BUFX2 U133 ( .A(n1251), .Y(n125) );
  BUFX2 U134 ( .A(n1252), .Y(n126) );
  BUFX2 U135 ( .A(n1253), .Y(n127) );
  BUFX2 U136 ( .A(n1254), .Y(n128) );
  BUFX2 U137 ( .A(n1255), .Y(n129) );
  BUFX2 U138 ( .A(n1258), .Y(n130) );
  AND2X1 U139 ( .A(n727), .B(n769), .Y(n1066) );
  INVX1 U140 ( .A(n1066), .Y(n131) );
  AND2X1 U141 ( .A(n726), .B(n769), .Y(n1067) );
  INVX1 U142 ( .A(n1067), .Y(n132) );
  AND2X1 U143 ( .A(n725), .B(n769), .Y(n1068) );
  INVX1 U144 ( .A(n1068), .Y(n133) );
  AND2X1 U145 ( .A(n724), .B(n769), .Y(n1069) );
  INVX1 U146 ( .A(n1069), .Y(n134) );
  AND2X1 U147 ( .A(n723), .B(n769), .Y(n1070) );
  INVX1 U148 ( .A(n1070), .Y(n135) );
  AND2X1 U149 ( .A(n713), .B(n770), .Y(n1081) );
  INVX1 U150 ( .A(n1081), .Y(n136) );
  AND2X1 U151 ( .A(n712), .B(n770), .Y(n1083) );
  INVX1 U152 ( .A(n1083), .Y(n137) );
  AND2X1 U153 ( .A(n711), .B(n770), .Y(n1084) );
  INVX1 U154 ( .A(n1084), .Y(n138) );
  AND2X1 U155 ( .A(n710), .B(n770), .Y(n1085) );
  INVX1 U156 ( .A(n1085), .Y(n139) );
  AND2X1 U157 ( .A(n709), .B(n770), .Y(n1086) );
  INVX1 U158 ( .A(n1086), .Y(n140) );
  AND2X1 U159 ( .A(n697), .B(n771), .Y(n1099) );
  INVX1 U160 ( .A(n1099), .Y(n141) );
  AND2X1 U161 ( .A(n696), .B(n771), .Y(n1100) );
  INVX1 U162 ( .A(n1100), .Y(n142) );
  AND2X1 U163 ( .A(n695), .B(n771), .Y(n1101) );
  INVX1 U164 ( .A(n1101), .Y(n143) );
  AND2X1 U165 ( .A(n694), .B(n771), .Y(n1102) );
  INVX1 U166 ( .A(n1102), .Y(n144) );
  AND2X1 U167 ( .A(n693), .B(n771), .Y(n1103) );
  INVX1 U168 ( .A(n1103), .Y(n145) );
  AND2X1 U169 ( .A(sendOut), .B(n772), .Y(n1115) );
  INVX1 U170 ( .A(n1115), .Y(n146) );
  AND2X1 U171 ( .A(n768), .B(n149), .Y(n1116) );
  INVX1 U172 ( .A(n1116), .Y(n147) );
  OR2X1 U173 ( .A(n1044), .B(n1045), .Y(n1047) );
  INVX1 U174 ( .A(n1047), .Y(n148) );
  AND2X1 U175 ( .A(n151), .B(n150), .Y(n1118) );
  INVX1 U176 ( .A(n1118), .Y(n149) );
  INVX1 U177 ( .A(InputBufferGrant[0]), .Y(n150) );
  INVX1 U178 ( .A(InputBufferGrant[1]), .Y(n151) );
  INVX8 U179 ( .A(reset), .Y(n909) );
  AND2X1 U601 ( .A(n698), .B(n771), .Y(n1098) );
  INVX1 U603 ( .A(n1098), .Y(n634) );
  AND2X1 U605 ( .A(n714), .B(n770), .Y(n1080) );
  INVX1 U607 ( .A(n1080), .Y(n635) );
  AND2X1 U609 ( .A(n728), .B(n769), .Y(n1065) );
  INVX1 U611 ( .A(n1065), .Y(n636) );
  AND2X1 U613 ( .A(n689), .B(n772), .Y(n1108) );
  INVX1 U615 ( .A(n1108), .Y(n637) );
  AND2X1 U617 ( .A(n699), .B(n771), .Y(n1097) );
  INVX1 U619 ( .A(n1097), .Y(n638) );
  AND2X1 U621 ( .A(n716), .B(n770), .Y(n1078) );
  INVX1 U623 ( .A(n1078), .Y(n639) );
  AND2X1 U625 ( .A(n729), .B(n769), .Y(n1064) );
  INVX1 U627 ( .A(n1064), .Y(n640) );
  AND2X1 U629 ( .A(n690), .B(n772), .Y(n1107) );
  INVX1 U631 ( .A(n1107), .Y(n641) );
  AND2X1 U633 ( .A(n702), .B(n771), .Y(n1094) );
  INVX1 U635 ( .A(n1094), .Y(n642) );
  AND2X1 U637 ( .A(n718), .B(n770), .Y(n1076) );
  INVX1 U639 ( .A(n1076), .Y(n643) );
  AND2X1 U641 ( .A(n730), .B(n769), .Y(n1063) );
  INVX1 U643 ( .A(n1063), .Y(n644) );
  AND2X1 U645 ( .A(n691), .B(n772), .Y(n1106) );
  INVX1 U647 ( .A(n1106), .Y(n645) );
  AND2X1 U649 ( .A(n700), .B(n771), .Y(n1096) );
  INVX1 U651 ( .A(n1096), .Y(n646) );
  AND2X1 U653 ( .A(n719), .B(n770), .Y(n1075) );
  INVX1 U655 ( .A(n1075), .Y(n647) );
  AND2X1 U657 ( .A(n731), .B(n769), .Y(n1062) );
  INVX1 U659 ( .A(n1062), .Y(n648) );
  AND2X1 U661 ( .A(n701), .B(n771), .Y(n1095) );
  INVX1 U663 ( .A(n1095), .Y(n649) );
  AND2X1 U665 ( .A(n717), .B(n770), .Y(n1077) );
  INVX1 U667 ( .A(n1077), .Y(n650) );
  AND2X1 U669 ( .A(n734), .B(n769), .Y(n1058) );
  INVX1 U671 ( .A(n1058), .Y(n651) );
  AND2X1 U673 ( .A(n740), .B(n768), .Y(n1052) );
  INVX1 U675 ( .A(n1052), .Y(n652) );
  AND2X1 U677 ( .A(n692), .B(n772), .Y(n1105) );
  INVX1 U679 ( .A(n1105), .Y(n653) );
  AND2X1 U680 ( .A(n704), .B(n771), .Y(n1091) );
  INVX1 U683 ( .A(n1091), .Y(n654) );
  AND2X1 U686 ( .A(n721), .B(n770), .Y(n1073) );
  INVX1 U687 ( .A(n1073), .Y(n655) );
  AND2X1 U688 ( .A(n741), .B(n769), .Y(n1051) );
  INVX1 U689 ( .A(n1051), .Y(n656) );
  AND2X1 U690 ( .A(n703), .B(n771), .Y(n1092) );
  INVX1 U691 ( .A(n1092), .Y(n657) );
  AND2X1 U692 ( .A(n715), .B(n770), .Y(n1079) );
  INVX1 U693 ( .A(n1079), .Y(n658) );
  AND2X1 U694 ( .A(n733), .B(n769), .Y(n1059) );
  INVX1 U695 ( .A(n1059), .Y(n659) );
  AND2X1 U696 ( .A(n737), .B(n768), .Y(n1055) );
  INVX1 U697 ( .A(n1055), .Y(n660) );
  AND2X1 U698 ( .A(n743), .B(n772), .Y(n1112) );
  INVX1 U699 ( .A(n1112), .Y(n661) );
  AND2X1 U700 ( .A(n707), .B(n771), .Y(n1088) );
  INVX1 U701 ( .A(n1088), .Y(n662) );
  AND2X1 U702 ( .A(n722), .B(n770), .Y(n1072) );
  INVX1 U703 ( .A(n1072), .Y(n663) );
  AND2X1 U704 ( .A(n738), .B(n769), .Y(n1054) );
  INVX1 U705 ( .A(n1054), .Y(n664) );
  AND2X1 U706 ( .A(n744), .B(n772), .Y(n1111) );
  INVX1 U707 ( .A(n1111), .Y(n665) );
  AND2X1 U708 ( .A(n705), .B(n771), .Y(n1090) );
  INVX1 U709 ( .A(n1090), .Y(n666) );
  AND2X1 U710 ( .A(n720), .B(n770), .Y(n1074) );
  INVX1 U711 ( .A(n1074), .Y(n667) );
  AND2X1 U712 ( .A(n735), .B(n769), .Y(n1057) );
  INVX1 U713 ( .A(n1057), .Y(n668) );
  AND2X1 U714 ( .A(n739), .B(n768), .Y(n1053) );
  INVX1 U715 ( .A(n1053), .Y(n669) );
  AND2X1 U716 ( .A(n745), .B(n772), .Y(n1110) );
  INVX1 U717 ( .A(n1110), .Y(n670) );
  AND2X1 U718 ( .A(n732), .B(n770), .Y(n1061) );
  INVX1 U719 ( .A(n1061), .Y(n671) );
  AND2X1 U720 ( .A(n742), .B(n769), .Y(n1050) );
  INVX1 U721 ( .A(n1050), .Y(n672) );
  AND2X1 U722 ( .A(n746), .B(n772), .Y(n1109) );
  INVX1 U723 ( .A(n1109), .Y(n673) );
  AND2X1 U724 ( .A(n748), .B(n771), .Y(n1093) );
  INVX1 U725 ( .A(n1093), .Y(n674) );
  AND2X1 U726 ( .A(n708), .B(n771), .Y(n1087) );
  INVX1 U727 ( .A(n1087), .Y(n675) );
  AND2X1 U728 ( .A(n736), .B(n768), .Y(n1056) );
  INVX1 U729 ( .A(n1056), .Y(n676) );
  AND2X1 U730 ( .A(n747), .B(n772), .Y(n1104) );
  INVX1 U731 ( .A(n1104), .Y(n677) );
  AND2X1 U732 ( .A(n750), .B(n769), .Y(n1071) );
  INVX1 U733 ( .A(n1071), .Y(n678) );
  AND2X1 U734 ( .A(n752), .B(n770), .Y(n1049) );
  INVX1 U735 ( .A(n1049), .Y(n679) );
  BUFX2 U736 ( .A(evenBufferFull), .Y(n680) );
  AND2X1 U737 ( .A(n706), .B(n771), .Y(n1089) );
  INVX1 U738 ( .A(n1089), .Y(n681) );
  AND2X1 U739 ( .A(n749), .B(n770), .Y(n1082) );
  INVX1 U740 ( .A(n1082), .Y(n682) );
  AND2X1 U741 ( .A(n751), .B(n769), .Y(n1060) );
  INVX1 U742 ( .A(n1060), .Y(n683) );
  AND2X1 U743 ( .A(n776), .B(n772), .Y(n1121) );
  INVX1 U744 ( .A(n1121), .Y(n684) );
  AND2X1 U745 ( .A(readyOut), .B(n1114), .Y(sendOut) );
  INVX1 U746 ( .A(sendOut), .Y(n685) );
  INVX1 U747 ( .A(n1113), .Y(n686) );
  BUFX2 U748 ( .A(priorityRegEven), .Y(n687) );
  AND2X1 U749 ( .A(n776), .B(n775), .Y(n1120) );
  INVX1 U750 ( .A(n1120), .Y(n688) );
  BUFX2 U751 ( .A(evenBuffer[63]), .Y(n689) );
  BUFX2 U752 ( .A(evenBuffer[62]), .Y(n690) );
  BUFX2 U753 ( .A(evenBuffer[61]), .Y(n691) );
  BUFX2 U754 ( .A(evenBuffer[60]), .Y(n692) );
  BUFX2 U755 ( .A(evenBuffer[59]), .Y(n693) );
  BUFX2 U756 ( .A(evenBuffer[58]), .Y(n694) );
  BUFX2 U757 ( .A(evenBuffer[57]), .Y(n695) );
  BUFX2 U758 ( .A(evenBuffer[56]), .Y(n696) );
  BUFX2 U759 ( .A(evenBuffer[55]), .Y(n697) );
  BUFX2 U760 ( .A(evenBuffer[54]), .Y(n698) );
  BUFX2 U761 ( .A(evenBuffer[53]), .Y(n699) );
  BUFX2 U762 ( .A(evenBuffer[52]), .Y(n700) );
  BUFX2 U763 ( .A(evenBuffer[51]), .Y(n701) );
  BUFX2 U764 ( .A(evenBuffer[50]), .Y(n702) );
  BUFX2 U765 ( .A(evenBuffer[49]), .Y(n703) );
  BUFX2 U766 ( .A(evenBuffer[48]), .Y(n704) );
  BUFX2 U767 ( .A(evenBuffer[47]), .Y(n705) );
  BUFX2 U768 ( .A(evenBuffer[46]), .Y(n706) );
  BUFX2 U769 ( .A(evenBuffer[45]), .Y(n707) );
  BUFX2 U770 ( .A(evenBuffer[44]), .Y(n708) );
  BUFX2 U771 ( .A(evenBuffer[43]), .Y(n709) );
  BUFX2 U772 ( .A(evenBuffer[42]), .Y(n710) );
  BUFX2 U773 ( .A(evenBuffer[41]), .Y(n711) );
  BUFX2 U774 ( .A(evenBuffer[40]), .Y(n712) );
  BUFX2 U775 ( .A(evenBuffer[39]), .Y(n713) );
  BUFX2 U776 ( .A(evenBuffer[38]), .Y(n714) );
  BUFX2 U777 ( .A(evenBuffer[37]), .Y(n715) );
  BUFX2 U778 ( .A(evenBuffer[36]), .Y(n716) );
  BUFX2 U779 ( .A(evenBuffer[35]), .Y(n717) );
  BUFX2 U780 ( .A(evenBuffer[34]), .Y(n718) );
  BUFX2 U781 ( .A(evenBuffer[33]), .Y(n719) );
  BUFX2 U782 ( .A(evenBuffer[32]), .Y(n720) );
  BUFX2 U783 ( .A(evenBuffer[31]), .Y(n721) );
  BUFX2 U784 ( .A(evenBuffer[30]), .Y(n722) );
  BUFX2 U785 ( .A(evenBuffer[29]), .Y(n723) );
  BUFX2 U786 ( .A(evenBuffer[28]), .Y(n724) );
  BUFX2 U787 ( .A(evenBuffer[27]), .Y(n725) );
  BUFX2 U788 ( .A(evenBuffer[26]), .Y(n726) );
  BUFX2 U789 ( .A(evenBuffer[25]), .Y(n727) );
  BUFX2 U790 ( .A(evenBuffer[24]), .Y(n728) );
  BUFX2 U791 ( .A(evenBuffer[23]), .Y(n729) );
  BUFX2 U792 ( .A(evenBuffer[22]), .Y(n730) );
  BUFX2 U793 ( .A(evenBuffer[21]), .Y(n731) );
  BUFX2 U794 ( .A(evenBuffer[20]), .Y(n732) );
  BUFX2 U795 ( .A(evenBuffer[19]), .Y(n733) );
  BUFX2 U796 ( .A(evenBuffer[18]), .Y(n734) );
  BUFX2 U797 ( .A(evenBuffer[17]), .Y(n735) );
  BUFX2 U798 ( .A(evenBuffer[16]), .Y(n736) );
  BUFX2 U799 ( .A(evenBuffer[15]), .Y(n737) );
  BUFX2 U800 ( .A(evenBuffer[14]), .Y(n738) );
  BUFX2 U801 ( .A(evenBuffer[13]), .Y(n739) );
  BUFX2 U802 ( .A(evenBuffer[12]), .Y(n740) );
  BUFX2 U803 ( .A(evenBuffer[11]), .Y(n741) );
  BUFX2 U804 ( .A(evenBuffer[10]), .Y(n742) );
  BUFX2 U805 ( .A(evenBuffer[9]), .Y(n743) );
  BUFX2 U806 ( .A(evenBuffer[8]), .Y(n744) );
  BUFX2 U807 ( .A(evenBuffer[7]), .Y(n745) );
  BUFX2 U808 ( .A(evenBuffer[6]), .Y(n746) );
  BUFX2 U809 ( .A(evenBuffer[5]), .Y(n747) );
  BUFX2 U810 ( .A(evenBuffer[4]), .Y(n748) );
  BUFX2 U811 ( .A(evenBuffer[3]), .Y(n749) );
  BUFX2 U812 ( .A(evenBuffer[2]), .Y(n750) );
  BUFX2 U813 ( .A(evenBuffer[1]), .Y(n751) );
  BUFX2 U814 ( .A(evenBuffer[0]), .Y(n752) );
  AND2X1 U815 ( .A(n768), .B(n1189), .Y(n1122) );
  INVX1 U816 ( .A(n1122), .Y(n753) );
  AND2X1 U817 ( .A(n1259), .B(n773), .Y(n1191) );
  INVX1 U818 ( .A(n1191), .Y(n754) );
  BUFX2 U819 ( .A(priorityRegOdd), .Y(n755) );
  INVX1 U820 ( .A(n774), .Y(n769) );
  INVX1 U821 ( .A(n774), .Y(n770) );
  INVX1 U822 ( .A(n774), .Y(n768) );
  INVX1 U823 ( .A(n773), .Y(n767) );
  INVX1 U824 ( .A(n773), .Y(n766) );
  INVX1 U825 ( .A(n775), .Y(n765) );
  INVX1 U826 ( .A(n775), .Y(n763) );
  INVX1 U827 ( .A(n775), .Y(n764) );
  INVX1 U828 ( .A(n773), .Y(n772) );
  INVX1 U829 ( .A(n760), .Y(n773) );
  INVX1 U830 ( .A(n760), .Y(n774) );
  INVX1 U831 ( .A(n1256), .Y(n758) );
  INVX1 U832 ( .A(n1187), .Y(n757) );
  INVX1 U833 ( .A(n762), .Y(n760) );
  INVX1 U834 ( .A(n1186), .Y(n756) );
  INVX1 U835 ( .A(n1257), .Y(n759) );
  INVX1 U836 ( .A(n775), .Y(n771) );
  INVX1 U837 ( .A(n761), .Y(n775) );
  INVX1 U838 ( .A(n762), .Y(n761) );
  INVX1 U839 ( .A(polarity), .Y(n762) );
  AND2X1 U840 ( .A(n772), .B(n780), .Y(n1044) );
  AND2X1 U841 ( .A(n777), .B(n774), .Y(n1045) );
  INVX1 U842 ( .A(n1119), .Y(n776) );
  INVX1 U843 ( .A(n755), .Y(n779) );
  INVX1 U844 ( .A(n741), .Y(n897) );
  INVX1 U845 ( .A(n740), .Y(n896) );
  INVX1 U846 ( .A(n739), .Y(n895) );
  INVX1 U847 ( .A(n738), .Y(n894) );
  INVX1 U848 ( .A(n737), .Y(n893) );
  INVX1 U849 ( .A(n736), .Y(n892) );
  INVX1 U850 ( .A(n735), .Y(n891) );
  INVX1 U851 ( .A(n734), .Y(n890) );
  INVX1 U852 ( .A(n733), .Y(n889) );
  INVX1 U853 ( .A(n732), .Y(n888) );
  INVX1 U854 ( .A(n731), .Y(n887) );
  INVX1 U855 ( .A(n730), .Y(n886) );
  INVX1 U856 ( .A(n729), .Y(n885) );
  INVX1 U857 ( .A(n727), .Y(n883) );
  INVX1 U858 ( .A(n728), .Y(n884) );
  INVX1 U859 ( .A(n726), .Y(n882) );
  INVX1 U860 ( .A(n725), .Y(n881) );
  INVX1 U861 ( .A(n724), .Y(n880) );
  INVX1 U862 ( .A(n723), .Y(n879) );
  INVX1 U863 ( .A(n722), .Y(n878) );
  INVX1 U864 ( .A(n721), .Y(n877) );
  INVX1 U865 ( .A(n720), .Y(n876) );
  INVX1 U866 ( .A(n719), .Y(n875) );
  INVX1 U867 ( .A(n718), .Y(n874) );
  INVX1 U868 ( .A(n717), .Y(n873) );
  INVX1 U869 ( .A(n716), .Y(n872) );
  INVX1 U870 ( .A(n715), .Y(n871) );
  INVX1 U871 ( .A(n714), .Y(n870) );
  INVX1 U872 ( .A(n713), .Y(n869) );
  INVX1 U873 ( .A(n712), .Y(n868) );
  INVX1 U874 ( .A(n711), .Y(n867) );
  INVX1 U875 ( .A(n710), .Y(n866) );
  INVX1 U876 ( .A(n709), .Y(n865) );
  INVX1 U877 ( .A(n708), .Y(n864) );
  INVX1 U878 ( .A(n707), .Y(n863) );
  INVX1 U879 ( .A(n706), .Y(n862) );
  INVX1 U880 ( .A(n705), .Y(n861) );
  INVX1 U881 ( .A(n704), .Y(n860) );
  INVX1 U882 ( .A(n703), .Y(n859) );
  INVX1 U883 ( .A(n702), .Y(n858) );
  INVX1 U884 ( .A(n701), .Y(n857) );
  INVX1 U885 ( .A(n700), .Y(n856) );
  INVX1 U886 ( .A(n699), .Y(n855) );
  INVX1 U887 ( .A(n698), .Y(n854) );
  INVX1 U888 ( .A(n697), .Y(n853) );
  INVX1 U889 ( .A(n696), .Y(n852) );
  INVX1 U890 ( .A(n695), .Y(n851) );
  INVX1 U891 ( .A(n694), .Y(n850) );
  INVX1 U892 ( .A(n693), .Y(n849) );
  INVX1 U893 ( .A(n692), .Y(n848) );
  INVX1 U894 ( .A(n691), .Y(n847) );
  INVX1 U895 ( .A(n690), .Y(n846) );
  INVX1 U896 ( .A(n752), .Y(n908) );
  INVX1 U897 ( .A(n751), .Y(n907) );
  INVX1 U898 ( .A(n750), .Y(n906) );
  INVX1 U899 ( .A(n749), .Y(n905) );
  INVX1 U900 ( .A(n748), .Y(n904) );
  INVX1 U901 ( .A(n747), .Y(n903) );
  INVX1 U902 ( .A(n746), .Y(n902) );
  INVX1 U903 ( .A(n745), .Y(n901) );
  INVX1 U904 ( .A(n744), .Y(n900) );
  INVX1 U905 ( .A(n743), .Y(n899) );
  INVX1 U906 ( .A(n742), .Y(n898) );
  INVX1 U907 ( .A(n689), .Y(n845) );
  INVX1 U908 ( .A(n687), .Y(n778) );
  INVX1 U909 ( .A(n680), .Y(n777) );
  INVX1 U910 ( .A(oddBufferFull), .Y(n780) );
  INVX1 U911 ( .A(oddBuffer[0]), .Y(n844) );
  INVX1 U912 ( .A(oddBuffer[1]), .Y(n843) );
  INVX1 U913 ( .A(oddBuffer[2]), .Y(n842) );
  INVX1 U914 ( .A(oddBuffer[3]), .Y(n841) );
  INVX1 U915 ( .A(oddBuffer[4]), .Y(n840) );
  INVX1 U916 ( .A(oddBuffer[5]), .Y(n839) );
  INVX1 U917 ( .A(oddBuffer[6]), .Y(n838) );
  INVX1 U918 ( .A(oddBuffer[7]), .Y(n837) );
  INVX1 U919 ( .A(oddBuffer[8]), .Y(n836) );
  INVX1 U920 ( .A(oddBuffer[9]), .Y(n835) );
  INVX1 U921 ( .A(oddBuffer[10]), .Y(n834) );
  INVX1 U922 ( .A(oddBuffer[11]), .Y(n833) );
  INVX1 U923 ( .A(oddBuffer[12]), .Y(n832) );
  INVX1 U924 ( .A(oddBuffer[13]), .Y(n831) );
  INVX1 U925 ( .A(oddBuffer[14]), .Y(n830) );
  INVX1 U926 ( .A(oddBuffer[15]), .Y(n829) );
  INVX1 U927 ( .A(oddBuffer[16]), .Y(n828) );
  INVX1 U928 ( .A(oddBuffer[17]), .Y(n827) );
  INVX1 U929 ( .A(oddBuffer[18]), .Y(n826) );
  INVX1 U930 ( .A(oddBuffer[19]), .Y(n825) );
  INVX1 U931 ( .A(oddBuffer[20]), .Y(n824) );
  INVX1 U932 ( .A(oddBuffer[21]), .Y(n823) );
  INVX1 U933 ( .A(oddBuffer[22]), .Y(n822) );
  INVX1 U934 ( .A(oddBuffer[23]), .Y(n821) );
  INVX1 U935 ( .A(oddBuffer[24]), .Y(n820) );
  INVX1 U936 ( .A(oddBuffer[25]), .Y(n819) );
  INVX1 U937 ( .A(oddBuffer[26]), .Y(n818) );
  INVX1 U938 ( .A(oddBuffer[27]), .Y(n817) );
  INVX1 U939 ( .A(oddBuffer[28]), .Y(n816) );
  INVX1 U940 ( .A(oddBuffer[29]), .Y(n815) );
  INVX1 U941 ( .A(oddBuffer[30]), .Y(n814) );
  INVX1 U942 ( .A(oddBuffer[31]), .Y(n813) );
  INVX1 U943 ( .A(oddBuffer[32]), .Y(n812) );
  INVX1 U944 ( .A(oddBuffer[33]), .Y(n811) );
  INVX1 U945 ( .A(oddBuffer[34]), .Y(n810) );
  INVX1 U946 ( .A(oddBuffer[35]), .Y(n809) );
  INVX1 U947 ( .A(oddBuffer[36]), .Y(n808) );
  INVX1 U948 ( .A(oddBuffer[37]), .Y(n807) );
  INVX1 U949 ( .A(oddBuffer[38]), .Y(n806) );
  INVX1 U950 ( .A(oddBuffer[39]), .Y(n805) );
  INVX1 U951 ( .A(oddBuffer[40]), .Y(n804) );
  INVX1 U952 ( .A(oddBuffer[41]), .Y(n803) );
  INVX1 U953 ( .A(oddBuffer[42]), .Y(n802) );
  INVX1 U954 ( .A(oddBuffer[43]), .Y(n801) );
  INVX1 U955 ( .A(oddBuffer[44]), .Y(n800) );
  INVX1 U956 ( .A(oddBuffer[45]), .Y(n799) );
  INVX1 U957 ( .A(oddBuffer[46]), .Y(n798) );
  INVX1 U958 ( .A(oddBuffer[47]), .Y(n797) );
  INVX1 U959 ( .A(oddBuffer[48]), .Y(n796) );
  INVX1 U960 ( .A(oddBuffer[49]), .Y(n795) );
  INVX1 U961 ( .A(oddBuffer[50]), .Y(n794) );
  INVX1 U962 ( .A(oddBuffer[51]), .Y(n793) );
  INVX1 U963 ( .A(oddBuffer[52]), .Y(n792) );
  INVX1 U964 ( .A(oddBuffer[53]), .Y(n791) );
  INVX1 U965 ( .A(oddBuffer[54]), .Y(n790) );
  INVX1 U966 ( .A(oddBuffer[55]), .Y(n789) );
  INVX1 U967 ( .A(oddBuffer[56]), .Y(n788) );
  INVX1 U968 ( .A(oddBuffer[57]), .Y(n787) );
  INVX1 U969 ( .A(oddBuffer[58]), .Y(n786) );
  INVX1 U970 ( .A(oddBuffer[59]), .Y(n785) );
  INVX1 U971 ( .A(oddBuffer[60]), .Y(n784) );
  INVX1 U972 ( .A(oddBuffer[61]), .Y(n783) );
  INVX1 U973 ( .A(oddBuffer[62]), .Y(n782) );
  INVX1 U974 ( .A(oddBuffer[63]), .Y(n781) );
endmodule


module outputBuffer_0 ( clk, reset, polarity, inputBufferRequest, dataIn0, 
        dataIn1, sendOut, readyOut, dataOut, InputBufferGrant );
  input [1:0] inputBufferRequest;
  input [63:0] dataIn0;
  input [63:0] dataIn1;
  output [63:0] dataOut;
  output [1:0] InputBufferGrant;
  input clk, reset, polarity, readyOut;
  output sendOut;
  wire   evenBufferFull, oddBufferFull, priorityRegEven, priorityRegOdd, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1189, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257;
  wire   [63:0] evenBuffer;
  wire   [63:0] oddBuffer;

  OAI21X1 U275 ( .A(n1257), .B(n843), .C(n130), .Y(n1039) );
  AOI22X1 U276 ( .A(dataIn1[63]), .B(n759), .C(dataIn0[63]), .D(n758), .Y(
        n1256) );
  OAI21X1 U277 ( .A(n1257), .B(n844), .C(n129), .Y(n1038) );
  AOI22X1 U278 ( .A(dataIn1[62]), .B(n759), .C(dataIn0[62]), .D(n758), .Y(
        n1253) );
  OAI21X1 U279 ( .A(n1257), .B(n845), .C(n128), .Y(n1037) );
  AOI22X1 U280 ( .A(dataIn1[61]), .B(n759), .C(dataIn0[61]), .D(n758), .Y(
        n1252) );
  OAI21X1 U281 ( .A(n1257), .B(n846), .C(n127), .Y(n1036) );
  AOI22X1 U282 ( .A(dataIn1[60]), .B(n759), .C(dataIn0[60]), .D(n758), .Y(
        n1251) );
  OAI21X1 U283 ( .A(n1257), .B(n847), .C(n126), .Y(n1035) );
  AOI22X1 U284 ( .A(dataIn1[59]), .B(n759), .C(dataIn0[59]), .D(n758), .Y(
        n1250) );
  OAI21X1 U285 ( .A(n1257), .B(n848), .C(n125), .Y(n1034) );
  AOI22X1 U286 ( .A(dataIn1[58]), .B(n759), .C(dataIn0[58]), .D(n758), .Y(
        n1249) );
  OAI21X1 U287 ( .A(n1257), .B(n849), .C(n124), .Y(n1033) );
  AOI22X1 U288 ( .A(dataIn1[57]), .B(n759), .C(dataIn0[57]), .D(n758), .Y(
        n1248) );
  OAI21X1 U289 ( .A(n1257), .B(n850), .C(n123), .Y(n1032) );
  AOI22X1 U290 ( .A(dataIn1[56]), .B(n759), .C(dataIn0[56]), .D(n758), .Y(
        n1247) );
  OAI21X1 U291 ( .A(n1257), .B(n851), .C(n122), .Y(n1031) );
  AOI22X1 U292 ( .A(dataIn1[55]), .B(n759), .C(dataIn0[55]), .D(n758), .Y(
        n1246) );
  OAI21X1 U293 ( .A(n1257), .B(n852), .C(n121), .Y(n1030) );
  AOI22X1 U294 ( .A(dataIn1[54]), .B(n759), .C(dataIn0[54]), .D(n758), .Y(
        n1245) );
  OAI21X1 U295 ( .A(n1257), .B(n853), .C(n120), .Y(n1029) );
  AOI22X1 U296 ( .A(dataIn1[53]), .B(n759), .C(dataIn0[53]), .D(n758), .Y(
        n1244) );
  OAI21X1 U297 ( .A(n1257), .B(n854), .C(n119), .Y(n1028) );
  AOI22X1 U298 ( .A(dataIn1[52]), .B(n759), .C(dataIn0[52]), .D(n758), .Y(
        n1243) );
  OAI21X1 U299 ( .A(n1257), .B(n855), .C(n118), .Y(n1027) );
  AOI22X1 U300 ( .A(dataIn1[51]), .B(n759), .C(dataIn0[51]), .D(n758), .Y(
        n1242) );
  OAI21X1 U301 ( .A(n1257), .B(n856), .C(n117), .Y(n1026) );
  AOI22X1 U302 ( .A(dataIn1[50]), .B(n759), .C(dataIn0[50]), .D(n758), .Y(
        n1241) );
  OAI21X1 U303 ( .A(n1257), .B(n857), .C(n116), .Y(n1025) );
  AOI22X1 U304 ( .A(dataIn1[49]), .B(n759), .C(dataIn0[49]), .D(n758), .Y(
        n1240) );
  OAI21X1 U305 ( .A(n1257), .B(n858), .C(n115), .Y(n1024) );
  AOI22X1 U306 ( .A(dataIn1[48]), .B(n759), .C(dataIn0[48]), .D(n758), .Y(
        n1239) );
  OAI21X1 U307 ( .A(n1257), .B(n859), .C(n114), .Y(n1023) );
  AOI22X1 U308 ( .A(dataIn1[47]), .B(n759), .C(dataIn0[47]), .D(n758), .Y(
        n1238) );
  OAI21X1 U309 ( .A(n1257), .B(n860), .C(n113), .Y(n1022) );
  AOI22X1 U310 ( .A(dataIn1[46]), .B(n759), .C(dataIn0[46]), .D(n758), .Y(
        n1237) );
  OAI21X1 U311 ( .A(n1257), .B(n861), .C(n112), .Y(n1021) );
  AOI22X1 U312 ( .A(dataIn1[45]), .B(n759), .C(dataIn0[45]), .D(n758), .Y(
        n1236) );
  OAI21X1 U313 ( .A(n1257), .B(n862), .C(n111), .Y(n1020) );
  AOI22X1 U314 ( .A(dataIn1[44]), .B(n759), .C(dataIn0[44]), .D(n758), .Y(
        n1235) );
  OAI21X1 U315 ( .A(n1257), .B(n863), .C(n110), .Y(n1019) );
  AOI22X1 U316 ( .A(dataIn1[43]), .B(n759), .C(dataIn0[43]), .D(n758), .Y(
        n1234) );
  OAI21X1 U317 ( .A(n1257), .B(n864), .C(n109), .Y(n1018) );
  AOI22X1 U318 ( .A(dataIn1[42]), .B(n759), .C(dataIn0[42]), .D(n758), .Y(
        n1233) );
  OAI21X1 U319 ( .A(n1257), .B(n865), .C(n108), .Y(n1017) );
  AOI22X1 U320 ( .A(dataIn1[41]), .B(n759), .C(dataIn0[41]), .D(n758), .Y(
        n1232) );
  OAI21X1 U321 ( .A(n1257), .B(n866), .C(n107), .Y(n1016) );
  AOI22X1 U322 ( .A(dataIn1[40]), .B(n759), .C(dataIn0[40]), .D(n758), .Y(
        n1231) );
  OAI21X1 U323 ( .A(n1257), .B(n867), .C(n106), .Y(n1015) );
  AOI22X1 U324 ( .A(dataIn1[39]), .B(n759), .C(dataIn0[39]), .D(n758), .Y(
        n1230) );
  OAI21X1 U325 ( .A(n1257), .B(n868), .C(n105), .Y(n1014) );
  AOI22X1 U326 ( .A(dataIn1[38]), .B(n759), .C(dataIn0[38]), .D(n758), .Y(
        n1229) );
  OAI21X1 U327 ( .A(n1257), .B(n869), .C(n104), .Y(n1013) );
  AOI22X1 U328 ( .A(dataIn1[37]), .B(n759), .C(dataIn0[37]), .D(n758), .Y(
        n1228) );
  OAI21X1 U329 ( .A(n1257), .B(n870), .C(n103), .Y(n1012) );
  AOI22X1 U330 ( .A(dataIn1[36]), .B(n759), .C(dataIn0[36]), .D(n758), .Y(
        n1227) );
  OAI21X1 U331 ( .A(n1257), .B(n871), .C(n102), .Y(n1011) );
  AOI22X1 U332 ( .A(dataIn1[35]), .B(n759), .C(dataIn0[35]), .D(n758), .Y(
        n1226) );
  OAI21X1 U333 ( .A(n1257), .B(n872), .C(n101), .Y(n1010) );
  AOI22X1 U334 ( .A(dataIn1[34]), .B(n759), .C(dataIn0[34]), .D(n758), .Y(
        n1225) );
  OAI21X1 U335 ( .A(n1257), .B(n873), .C(n100), .Y(n1009) );
  AOI22X1 U336 ( .A(dataIn1[33]), .B(n759), .C(dataIn0[33]), .D(n758), .Y(
        n1224) );
  OAI21X1 U337 ( .A(n1257), .B(n874), .C(n99), .Y(n1008) );
  AOI22X1 U338 ( .A(dataIn1[32]), .B(n759), .C(dataIn0[32]), .D(n758), .Y(
        n1223) );
  OAI21X1 U339 ( .A(n1257), .B(n875), .C(n98), .Y(n1007) );
  AOI22X1 U340 ( .A(dataIn1[31]), .B(n759), .C(dataIn0[31]), .D(n758), .Y(
        n1222) );
  OAI21X1 U341 ( .A(n1257), .B(n876), .C(n97), .Y(n1006) );
  AOI22X1 U342 ( .A(dataIn1[30]), .B(n759), .C(dataIn0[30]), .D(n758), .Y(
        n1221) );
  OAI21X1 U343 ( .A(n1257), .B(n877), .C(n96), .Y(n1005) );
  AOI22X1 U344 ( .A(dataIn1[29]), .B(n759), .C(dataIn0[29]), .D(n758), .Y(
        n1220) );
  OAI21X1 U345 ( .A(n1257), .B(n878), .C(n95), .Y(n1004) );
  AOI22X1 U346 ( .A(dataIn1[28]), .B(n759), .C(dataIn0[28]), .D(n758), .Y(
        n1219) );
  OAI21X1 U347 ( .A(n1257), .B(n879), .C(n94), .Y(n1003) );
  AOI22X1 U348 ( .A(dataIn1[27]), .B(n759), .C(dataIn0[27]), .D(n758), .Y(
        n1218) );
  OAI21X1 U349 ( .A(n1257), .B(n880), .C(n93), .Y(n1002) );
  AOI22X1 U350 ( .A(dataIn1[26]), .B(n759), .C(dataIn0[26]), .D(n758), .Y(
        n1217) );
  OAI21X1 U351 ( .A(n1257), .B(n881), .C(n92), .Y(n1001) );
  AOI22X1 U352 ( .A(dataIn1[25]), .B(n759), .C(dataIn0[25]), .D(n758), .Y(
        n1216) );
  OAI21X1 U353 ( .A(n1257), .B(n882), .C(n91), .Y(n1000) );
  AOI22X1 U354 ( .A(dataIn1[24]), .B(n759), .C(dataIn0[24]), .D(n758), .Y(
        n1215) );
  OAI21X1 U355 ( .A(n1257), .B(n883), .C(n90), .Y(n999) );
  AOI22X1 U356 ( .A(dataIn1[23]), .B(n759), .C(dataIn0[23]), .D(n758), .Y(
        n1214) );
  OAI21X1 U357 ( .A(n1257), .B(n884), .C(n89), .Y(n998) );
  AOI22X1 U358 ( .A(dataIn1[22]), .B(n759), .C(dataIn0[22]), .D(n758), .Y(
        n1213) );
  OAI21X1 U359 ( .A(n1257), .B(n885), .C(n88), .Y(n997) );
  AOI22X1 U360 ( .A(dataIn1[21]), .B(n759), .C(dataIn0[21]), .D(n758), .Y(
        n1212) );
  OAI21X1 U361 ( .A(n1257), .B(n886), .C(n87), .Y(n996) );
  AOI22X1 U362 ( .A(dataIn1[20]), .B(n759), .C(dataIn0[20]), .D(n758), .Y(
        n1211) );
  OAI21X1 U363 ( .A(n1257), .B(n887), .C(n86), .Y(n995) );
  AOI22X1 U364 ( .A(dataIn1[19]), .B(n759), .C(dataIn0[19]), .D(n758), .Y(
        n1210) );
  OAI21X1 U365 ( .A(n1257), .B(n888), .C(n85), .Y(n994) );
  AOI22X1 U366 ( .A(dataIn1[18]), .B(n759), .C(dataIn0[18]), .D(n758), .Y(
        n1209) );
  OAI21X1 U367 ( .A(n1257), .B(n889), .C(n84), .Y(n993) );
  AOI22X1 U368 ( .A(dataIn1[17]), .B(n759), .C(dataIn0[17]), .D(n758), .Y(
        n1208) );
  OAI21X1 U369 ( .A(n1257), .B(n890), .C(n83), .Y(n992) );
  AOI22X1 U370 ( .A(dataIn1[16]), .B(n759), .C(dataIn0[16]), .D(n758), .Y(
        n1207) );
  OAI21X1 U371 ( .A(n1257), .B(n891), .C(n82), .Y(n991) );
  AOI22X1 U372 ( .A(dataIn1[15]), .B(n759), .C(dataIn0[15]), .D(n758), .Y(
        n1206) );
  OAI21X1 U373 ( .A(n1257), .B(n892), .C(n81), .Y(n990) );
  AOI22X1 U374 ( .A(dataIn1[14]), .B(n759), .C(dataIn0[14]), .D(n758), .Y(
        n1205) );
  OAI21X1 U375 ( .A(n1257), .B(n893), .C(n80), .Y(n989) );
  AOI22X1 U376 ( .A(dataIn1[13]), .B(n759), .C(dataIn0[13]), .D(n758), .Y(
        n1204) );
  OAI21X1 U377 ( .A(n1257), .B(n894), .C(n79), .Y(n988) );
  AOI22X1 U378 ( .A(dataIn1[12]), .B(n759), .C(dataIn0[12]), .D(n758), .Y(
        n1203) );
  OAI21X1 U379 ( .A(n1257), .B(n895), .C(n78), .Y(n987) );
  AOI22X1 U380 ( .A(dataIn1[11]), .B(n759), .C(dataIn0[11]), .D(n758), .Y(
        n1202) );
  OAI21X1 U381 ( .A(n1257), .B(n896), .C(n77), .Y(n986) );
  AOI22X1 U382 ( .A(dataIn1[10]), .B(n759), .C(dataIn0[10]), .D(n758), .Y(
        n1201) );
  OAI21X1 U383 ( .A(n1257), .B(n897), .C(n76), .Y(n985) );
  AOI22X1 U384 ( .A(dataIn1[9]), .B(n759), .C(dataIn0[9]), .D(n758), .Y(n1200)
         );
  OAI21X1 U385 ( .A(n1257), .B(n898), .C(n75), .Y(n984) );
  AOI22X1 U386 ( .A(dataIn1[8]), .B(n759), .C(dataIn0[8]), .D(n758), .Y(n1199)
         );
  OAI21X1 U387 ( .A(n1257), .B(n899), .C(n74), .Y(n983) );
  AOI22X1 U388 ( .A(dataIn1[7]), .B(n759), .C(dataIn0[7]), .D(n758), .Y(n1198)
         );
  OAI21X1 U389 ( .A(n1257), .B(n900), .C(n73), .Y(n982) );
  AOI22X1 U390 ( .A(dataIn1[6]), .B(n759), .C(dataIn0[6]), .D(n758), .Y(n1197)
         );
  OAI21X1 U391 ( .A(n1257), .B(n901), .C(n72), .Y(n981) );
  AOI22X1 U392 ( .A(dataIn1[5]), .B(n759), .C(dataIn0[5]), .D(n758), .Y(n1196)
         );
  OAI21X1 U393 ( .A(n1257), .B(n902), .C(n71), .Y(n980) );
  AOI22X1 U394 ( .A(dataIn1[4]), .B(n759), .C(dataIn0[4]), .D(n758), .Y(n1195)
         );
  OAI21X1 U395 ( .A(n1257), .B(n903), .C(n70), .Y(n979) );
  AOI22X1 U396 ( .A(dataIn1[3]), .B(n759), .C(dataIn0[3]), .D(n758), .Y(n1194)
         );
  OAI21X1 U397 ( .A(n1257), .B(n904), .C(n69), .Y(n978) );
  AOI22X1 U398 ( .A(dataIn1[2]), .B(n759), .C(dataIn0[2]), .D(n758), .Y(n1193)
         );
  OAI21X1 U399 ( .A(n1257), .B(n905), .C(n68), .Y(n977) );
  AOI22X1 U400 ( .A(dataIn1[1]), .B(n759), .C(dataIn0[1]), .D(n758), .Y(n1192)
         );
  OAI21X1 U401 ( .A(n1257), .B(n906), .C(n67), .Y(n976) );
  AOI22X1 U402 ( .A(dataIn1[0]), .B(n759), .C(dataIn0[0]), .D(n758), .Y(n1191)
         );
  OAI21X1 U405 ( .A(n1187), .B(n779), .C(n66), .Y(n975) );
  AOI22X1 U406 ( .A(n757), .B(dataIn1[63]), .C(n756), .D(dataIn0[63]), .Y(
        n1186) );
  OAI21X1 U407 ( .A(n1187), .B(n780), .C(n65), .Y(n974) );
  AOI22X1 U408 ( .A(n757), .B(dataIn1[62]), .C(n756), .D(dataIn0[62]), .Y(
        n1183) );
  OAI21X1 U409 ( .A(n1187), .B(n781), .C(n64), .Y(n973) );
  AOI22X1 U410 ( .A(n757), .B(dataIn1[61]), .C(n756), .D(dataIn0[61]), .Y(
        n1182) );
  OAI21X1 U411 ( .A(n1187), .B(n782), .C(n63), .Y(n972) );
  AOI22X1 U412 ( .A(n757), .B(dataIn1[60]), .C(n756), .D(dataIn0[60]), .Y(
        n1181) );
  OAI21X1 U413 ( .A(n1187), .B(n783), .C(n62), .Y(n971) );
  AOI22X1 U414 ( .A(n757), .B(dataIn1[59]), .C(n756), .D(dataIn0[59]), .Y(
        n1180) );
  OAI21X1 U415 ( .A(n1187), .B(n784), .C(n61), .Y(n970) );
  AOI22X1 U416 ( .A(n757), .B(dataIn1[58]), .C(n756), .D(dataIn0[58]), .Y(
        n1179) );
  OAI21X1 U417 ( .A(n1187), .B(n785), .C(n60), .Y(n969) );
  AOI22X1 U418 ( .A(n757), .B(dataIn1[57]), .C(n756), .D(dataIn0[57]), .Y(
        n1178) );
  OAI21X1 U419 ( .A(n1187), .B(n786), .C(n59), .Y(n968) );
  AOI22X1 U420 ( .A(n757), .B(dataIn1[56]), .C(n756), .D(dataIn0[56]), .Y(
        n1177) );
  OAI21X1 U421 ( .A(n1187), .B(n787), .C(n58), .Y(n967) );
  AOI22X1 U422 ( .A(n757), .B(dataIn1[55]), .C(n756), .D(dataIn0[55]), .Y(
        n1176) );
  OAI21X1 U423 ( .A(n1187), .B(n788), .C(n57), .Y(n966) );
  AOI22X1 U424 ( .A(n757), .B(dataIn1[54]), .C(n756), .D(dataIn0[54]), .Y(
        n1175) );
  OAI21X1 U425 ( .A(n1187), .B(n789), .C(n56), .Y(n965) );
  AOI22X1 U426 ( .A(n757), .B(dataIn1[53]), .C(n756), .D(dataIn0[53]), .Y(
        n1174) );
  OAI21X1 U427 ( .A(n1187), .B(n790), .C(n55), .Y(n964) );
  AOI22X1 U428 ( .A(n757), .B(dataIn1[52]), .C(n756), .D(dataIn0[52]), .Y(
        n1173) );
  OAI21X1 U429 ( .A(n1187), .B(n791), .C(n54), .Y(n963) );
  AOI22X1 U430 ( .A(n757), .B(dataIn1[51]), .C(n756), .D(dataIn0[51]), .Y(
        n1172) );
  OAI21X1 U431 ( .A(n1187), .B(n792), .C(n53), .Y(n962) );
  AOI22X1 U432 ( .A(n757), .B(dataIn1[50]), .C(n756), .D(dataIn0[50]), .Y(
        n1171) );
  OAI21X1 U433 ( .A(n1187), .B(n793), .C(n52), .Y(n961) );
  AOI22X1 U434 ( .A(n757), .B(dataIn1[49]), .C(n756), .D(dataIn0[49]), .Y(
        n1170) );
  OAI21X1 U435 ( .A(n1187), .B(n794), .C(n51), .Y(n960) );
  AOI22X1 U436 ( .A(n757), .B(dataIn1[48]), .C(n756), .D(dataIn0[48]), .Y(
        n1169) );
  OAI21X1 U437 ( .A(n1187), .B(n795), .C(n50), .Y(n959) );
  AOI22X1 U438 ( .A(n757), .B(dataIn1[47]), .C(n756), .D(dataIn0[47]), .Y(
        n1168) );
  OAI21X1 U439 ( .A(n1187), .B(n796), .C(n49), .Y(n958) );
  AOI22X1 U440 ( .A(n757), .B(dataIn1[46]), .C(n756), .D(dataIn0[46]), .Y(
        n1167) );
  OAI21X1 U441 ( .A(n1187), .B(n797), .C(n48), .Y(n957) );
  AOI22X1 U442 ( .A(n757), .B(dataIn1[45]), .C(n756), .D(dataIn0[45]), .Y(
        n1166) );
  OAI21X1 U443 ( .A(n1187), .B(n798), .C(n47), .Y(n956) );
  AOI22X1 U444 ( .A(n757), .B(dataIn1[44]), .C(n756), .D(dataIn0[44]), .Y(
        n1165) );
  OAI21X1 U445 ( .A(n1187), .B(n799), .C(n46), .Y(n955) );
  AOI22X1 U446 ( .A(n757), .B(dataIn1[43]), .C(n756), .D(dataIn0[43]), .Y(
        n1164) );
  OAI21X1 U447 ( .A(n1187), .B(n800), .C(n45), .Y(n954) );
  AOI22X1 U448 ( .A(n757), .B(dataIn1[42]), .C(n756), .D(dataIn0[42]), .Y(
        n1163) );
  OAI21X1 U449 ( .A(n1187), .B(n801), .C(n44), .Y(n953) );
  AOI22X1 U450 ( .A(n757), .B(dataIn1[41]), .C(n756), .D(dataIn0[41]), .Y(
        n1162) );
  OAI21X1 U451 ( .A(n1187), .B(n802), .C(n43), .Y(n952) );
  AOI22X1 U452 ( .A(n757), .B(dataIn1[40]), .C(n756), .D(dataIn0[40]), .Y(
        n1161) );
  OAI21X1 U453 ( .A(n1187), .B(n803), .C(n42), .Y(n951) );
  AOI22X1 U454 ( .A(n757), .B(dataIn1[39]), .C(n756), .D(dataIn0[39]), .Y(
        n1160) );
  OAI21X1 U455 ( .A(n1187), .B(n804), .C(n41), .Y(n950) );
  AOI22X1 U456 ( .A(n757), .B(dataIn1[38]), .C(n756), .D(dataIn0[38]), .Y(
        n1159) );
  OAI21X1 U457 ( .A(n1187), .B(n805), .C(n40), .Y(n949) );
  AOI22X1 U458 ( .A(n757), .B(dataIn1[37]), .C(n756), .D(dataIn0[37]), .Y(
        n1158) );
  OAI21X1 U459 ( .A(n1187), .B(n806), .C(n39), .Y(n948) );
  AOI22X1 U460 ( .A(n757), .B(dataIn1[36]), .C(n756), .D(dataIn0[36]), .Y(
        n1157) );
  OAI21X1 U461 ( .A(n1187), .B(n807), .C(n38), .Y(n947) );
  AOI22X1 U462 ( .A(n757), .B(dataIn1[35]), .C(n756), .D(dataIn0[35]), .Y(
        n1156) );
  OAI21X1 U463 ( .A(n1187), .B(n808), .C(n37), .Y(n946) );
  AOI22X1 U464 ( .A(n757), .B(dataIn1[34]), .C(n756), .D(dataIn0[34]), .Y(
        n1155) );
  OAI21X1 U465 ( .A(n1187), .B(n809), .C(n36), .Y(n945) );
  AOI22X1 U466 ( .A(n757), .B(dataIn1[33]), .C(n756), .D(dataIn0[33]), .Y(
        n1154) );
  OAI21X1 U467 ( .A(n1187), .B(n810), .C(n35), .Y(n944) );
  AOI22X1 U468 ( .A(n757), .B(dataIn1[32]), .C(n756), .D(dataIn0[32]), .Y(
        n1153) );
  OAI21X1 U469 ( .A(n1187), .B(n811), .C(n34), .Y(n943) );
  AOI22X1 U470 ( .A(n757), .B(dataIn1[31]), .C(n756), .D(dataIn0[31]), .Y(
        n1152) );
  OAI21X1 U471 ( .A(n1187), .B(n812), .C(n33), .Y(n942) );
  AOI22X1 U472 ( .A(n757), .B(dataIn1[30]), .C(n756), .D(dataIn0[30]), .Y(
        n1151) );
  OAI21X1 U473 ( .A(n1187), .B(n813), .C(n32), .Y(n941) );
  AOI22X1 U474 ( .A(n757), .B(dataIn1[29]), .C(n756), .D(dataIn0[29]), .Y(
        n1150) );
  OAI21X1 U475 ( .A(n1187), .B(n814), .C(n31), .Y(n940) );
  AOI22X1 U476 ( .A(n757), .B(dataIn1[28]), .C(n756), .D(dataIn0[28]), .Y(
        n1149) );
  OAI21X1 U477 ( .A(n1187), .B(n815), .C(n30), .Y(n939) );
  AOI22X1 U478 ( .A(n757), .B(dataIn1[27]), .C(n756), .D(dataIn0[27]), .Y(
        n1148) );
  OAI21X1 U479 ( .A(n1187), .B(n816), .C(n29), .Y(n938) );
  AOI22X1 U480 ( .A(n757), .B(dataIn1[26]), .C(n756), .D(dataIn0[26]), .Y(
        n1147) );
  OAI21X1 U481 ( .A(n1187), .B(n817), .C(n28), .Y(n937) );
  AOI22X1 U482 ( .A(n757), .B(dataIn1[25]), .C(n756), .D(dataIn0[25]), .Y(
        n1146) );
  OAI21X1 U483 ( .A(n1187), .B(n818), .C(n27), .Y(n936) );
  AOI22X1 U484 ( .A(n757), .B(dataIn1[24]), .C(n756), .D(dataIn0[24]), .Y(
        n1145) );
  OAI21X1 U485 ( .A(n1187), .B(n819), .C(n26), .Y(n935) );
  AOI22X1 U486 ( .A(n757), .B(dataIn1[23]), .C(n756), .D(dataIn0[23]), .Y(
        n1144) );
  OAI21X1 U487 ( .A(n1187), .B(n820), .C(n25), .Y(n934) );
  AOI22X1 U488 ( .A(n757), .B(dataIn1[22]), .C(n756), .D(dataIn0[22]), .Y(
        n1143) );
  OAI21X1 U489 ( .A(n1187), .B(n821), .C(n24), .Y(n933) );
  AOI22X1 U490 ( .A(n757), .B(dataIn1[21]), .C(n756), .D(dataIn0[21]), .Y(
        n1142) );
  OAI21X1 U491 ( .A(n1187), .B(n822), .C(n23), .Y(n932) );
  AOI22X1 U492 ( .A(n757), .B(dataIn1[20]), .C(n756), .D(dataIn0[20]), .Y(
        n1141) );
  OAI21X1 U493 ( .A(n1187), .B(n823), .C(n22), .Y(n931) );
  AOI22X1 U494 ( .A(n757), .B(dataIn1[19]), .C(n756), .D(dataIn0[19]), .Y(
        n1140) );
  OAI21X1 U495 ( .A(n1187), .B(n824), .C(n21), .Y(n930) );
  AOI22X1 U496 ( .A(n757), .B(dataIn1[18]), .C(n756), .D(dataIn0[18]), .Y(
        n1139) );
  OAI21X1 U497 ( .A(n1187), .B(n825), .C(n20), .Y(n929) );
  AOI22X1 U498 ( .A(n757), .B(dataIn1[17]), .C(n756), .D(dataIn0[17]), .Y(
        n1138) );
  OAI21X1 U499 ( .A(n1187), .B(n826), .C(n19), .Y(n928) );
  AOI22X1 U500 ( .A(n757), .B(dataIn1[16]), .C(n756), .D(dataIn0[16]), .Y(
        n1137) );
  OAI21X1 U501 ( .A(n1187), .B(n827), .C(n18), .Y(n927) );
  AOI22X1 U502 ( .A(n757), .B(dataIn1[15]), .C(n756), .D(dataIn0[15]), .Y(
        n1136) );
  OAI21X1 U503 ( .A(n1187), .B(n828), .C(n17), .Y(n926) );
  AOI22X1 U504 ( .A(n757), .B(dataIn1[14]), .C(n756), .D(dataIn0[14]), .Y(
        n1135) );
  OAI21X1 U505 ( .A(n1187), .B(n829), .C(n16), .Y(n925) );
  AOI22X1 U506 ( .A(n757), .B(dataIn1[13]), .C(n756), .D(dataIn0[13]), .Y(
        n1134) );
  OAI21X1 U507 ( .A(n1187), .B(n830), .C(n15), .Y(n924) );
  AOI22X1 U508 ( .A(n757), .B(dataIn1[12]), .C(n756), .D(dataIn0[12]), .Y(
        n1133) );
  OAI21X1 U509 ( .A(n1187), .B(n831), .C(n14), .Y(n923) );
  AOI22X1 U510 ( .A(n757), .B(dataIn1[11]), .C(n756), .D(dataIn0[11]), .Y(
        n1132) );
  OAI21X1 U511 ( .A(n1187), .B(n832), .C(n13), .Y(n922) );
  AOI22X1 U512 ( .A(n757), .B(dataIn1[10]), .C(n756), .D(dataIn0[10]), .Y(
        n1131) );
  OAI21X1 U513 ( .A(n1187), .B(n833), .C(n12), .Y(n921) );
  AOI22X1 U514 ( .A(n757), .B(dataIn1[9]), .C(n756), .D(dataIn0[9]), .Y(n1130)
         );
  OAI21X1 U515 ( .A(n1187), .B(n834), .C(n11), .Y(n920) );
  AOI22X1 U516 ( .A(n757), .B(dataIn1[8]), .C(n756), .D(dataIn0[8]), .Y(n1129)
         );
  OAI21X1 U517 ( .A(n1187), .B(n835), .C(n10), .Y(n919) );
  AOI22X1 U518 ( .A(n757), .B(dataIn1[7]), .C(n756), .D(dataIn0[7]), .Y(n1128)
         );
  OAI21X1 U519 ( .A(n1187), .B(n836), .C(n9), .Y(n918) );
  AOI22X1 U520 ( .A(n757), .B(dataIn1[6]), .C(n756), .D(dataIn0[6]), .Y(n1127)
         );
  OAI21X1 U521 ( .A(n1187), .B(n837), .C(n8), .Y(n917) );
  AOI22X1 U522 ( .A(n757), .B(dataIn1[5]), .C(n756), .D(dataIn0[5]), .Y(n1126)
         );
  OAI21X1 U523 ( .A(n1187), .B(n838), .C(n7), .Y(n916) );
  AOI22X1 U524 ( .A(n757), .B(dataIn1[4]), .C(n756), .D(dataIn0[4]), .Y(n1125)
         );
  OAI21X1 U525 ( .A(n1187), .B(n839), .C(n6), .Y(n915) );
  AOI22X1 U526 ( .A(n757), .B(dataIn1[3]), .C(n756), .D(dataIn0[3]), .Y(n1124)
         );
  OAI21X1 U527 ( .A(n1187), .B(n840), .C(n5), .Y(n914) );
  AOI22X1 U528 ( .A(n757), .B(dataIn1[2]), .C(n756), .D(dataIn0[2]), .Y(n1123)
         );
  OAI21X1 U529 ( .A(n1187), .B(n841), .C(n4), .Y(n913) );
  AOI22X1 U530 ( .A(n757), .B(dataIn1[1]), .C(n756), .D(dataIn0[1]), .Y(n1122)
         );
  OAI21X1 U531 ( .A(n1187), .B(n842), .C(n3), .Y(n912) );
  AOI22X1 U532 ( .A(n757), .B(dataIn1[0]), .C(n756), .D(dataIn0[0]), .Y(n1121)
         );
  XNOR2X1 U535 ( .A(n755), .B(n684), .Y(n911) );
  XNOR2X1 U537 ( .A(n687), .B(n688), .Y(n910) );
  NAND3X1 U539 ( .A(inputBufferRequest[1]), .B(n149), .C(inputBufferRequest[0]), .Y(n1117) );
  OAI21X1 U540 ( .A(n778), .B(n1187), .C(n753), .Y(n909) );
  OAI21X1 U542 ( .A(n762), .B(n685), .C(n147), .Y(n1187) );
  OAI21X1 U544 ( .A(n775), .B(n1257), .C(n754), .Y(n908) );
  OAI21X1 U546 ( .A(n762), .B(n1116), .C(n146), .Y(n1257) );
  OAI21X1 U549 ( .A(n762), .B(n778), .C(n686), .Y(n1112) );
  OAI21X1 U552 ( .A(n762), .B(n833), .C(n661), .Y(dataOut[9]) );
  OAI21X1 U554 ( .A(n762), .B(n834), .C(n665), .Y(dataOut[8]) );
  OAI21X1 U556 ( .A(n762), .B(n835), .C(n670), .Y(dataOut[7]) );
  OAI21X1 U558 ( .A(n763), .B(n836), .C(n673), .Y(dataOut[6]) );
  OAI21X1 U560 ( .A(n763), .B(n779), .C(n637), .Y(dataOut[63]) );
  OAI21X1 U562 ( .A(n762), .B(n780), .C(n641), .Y(dataOut[62]) );
  OAI21X1 U564 ( .A(n763), .B(n781), .C(n645), .Y(dataOut[61]) );
  OAI21X1 U566 ( .A(n763), .B(n782), .C(n653), .Y(dataOut[60]) );
  OAI21X1 U568 ( .A(n763), .B(n837), .C(n677), .Y(dataOut[5]) );
  OAI21X1 U570 ( .A(n763), .B(n783), .C(n145), .Y(dataOut[59]) );
  OAI21X1 U572 ( .A(n764), .B(n784), .C(n144), .Y(dataOut[58]) );
  OAI21X1 U574 ( .A(n763), .B(n785), .C(n143), .Y(dataOut[57]) );
  OAI21X1 U576 ( .A(n764), .B(n786), .C(n142), .Y(dataOut[56]) );
  OAI21X1 U578 ( .A(n764), .B(n787), .C(n141), .Y(dataOut[55]) );
  OAI21X1 U580 ( .A(n762), .B(n788), .C(n634), .Y(dataOut[54]) );
  OAI21X1 U582 ( .A(n764), .B(n789), .C(n638), .Y(dataOut[53]) );
  OAI21X1 U584 ( .A(n764), .B(n790), .C(n646), .Y(dataOut[52]) );
  OAI21X1 U586 ( .A(n764), .B(n791), .C(n649), .Y(dataOut[51]) );
  OAI21X1 U588 ( .A(n765), .B(n792), .C(n642), .Y(dataOut[50]) );
  OAI21X1 U590 ( .A(n765), .B(n838), .C(n674), .Y(dataOut[4]) );
  OAI21X1 U592 ( .A(n764), .B(n793), .C(n657), .Y(dataOut[49]) );
  OAI21X1 U594 ( .A(n765), .B(n794), .C(n654), .Y(dataOut[48]) );
  OAI21X1 U596 ( .A(n765), .B(n795), .C(n666), .Y(dataOut[47]) );
  OAI21X1 U598 ( .A(n763), .B(n796), .C(n681), .Y(dataOut[46]) );
  OAI21X1 U600 ( .A(n766), .B(n797), .C(n662), .Y(dataOut[45]) );
  OAI21X1 U602 ( .A(n766), .B(n798), .C(n675), .Y(dataOut[44]) );
  OAI21X1 U604 ( .A(n764), .B(n799), .C(n140), .Y(dataOut[43]) );
  OAI21X1 U606 ( .A(n766), .B(n800), .C(n139), .Y(dataOut[42]) );
  OAI21X1 U608 ( .A(n766), .B(n801), .C(n138), .Y(dataOut[41]) );
  OAI21X1 U610 ( .A(n765), .B(n802), .C(n137), .Y(dataOut[40]) );
  OAI21X1 U612 ( .A(n766), .B(n839), .C(n682), .Y(dataOut[3]) );
  OAI21X1 U614 ( .A(n766), .B(n803), .C(n136), .Y(dataOut[39]) );
  OAI21X1 U616 ( .A(n764), .B(n804), .C(n635), .Y(dataOut[38]) );
  OAI21X1 U618 ( .A(n766), .B(n805), .C(n658), .Y(dataOut[37]) );
  OAI21X1 U620 ( .A(n767), .B(n806), .C(n639), .Y(dataOut[36]) );
  OAI21X1 U622 ( .A(n765), .B(n807), .C(n650), .Y(dataOut[35]) );
  OAI21X1 U624 ( .A(n767), .B(n808), .C(n643), .Y(dataOut[34]) );
  OAI21X1 U626 ( .A(n767), .B(n809), .C(n647), .Y(dataOut[33]) );
  OAI21X1 U628 ( .A(n766), .B(n810), .C(n667), .Y(dataOut[32]) );
  OAI21X1 U630 ( .A(n767), .B(n811), .C(n655), .Y(dataOut[31]) );
  OAI21X1 U632 ( .A(n767), .B(n812), .C(n663), .Y(dataOut[30]) );
  OAI21X1 U634 ( .A(n765), .B(n840), .C(n678), .Y(dataOut[2]) );
  OAI21X1 U636 ( .A(n766), .B(n813), .C(n135), .Y(dataOut[29]) );
  OAI21X1 U638 ( .A(n767), .B(n814), .C(n134), .Y(dataOut[28]) );
  OAI21X1 U640 ( .A(n767), .B(n815), .C(n133), .Y(dataOut[27]) );
  OAI21X1 U642 ( .A(n765), .B(n816), .C(n132), .Y(dataOut[26]) );
  OAI21X1 U644 ( .A(n766), .B(n817), .C(n131), .Y(dataOut[25]) );
  OAI21X1 U646 ( .A(n766), .B(n818), .C(n636), .Y(dataOut[24]) );
  OAI21X1 U648 ( .A(n765), .B(n819), .C(n640), .Y(dataOut[23]) );
  OAI21X1 U650 ( .A(n766), .B(n820), .C(n644), .Y(dataOut[22]) );
  OAI21X1 U652 ( .A(n765), .B(n821), .C(n648), .Y(dataOut[21]) );
  OAI21X1 U654 ( .A(n764), .B(n822), .C(n671), .Y(dataOut[20]) );
  OAI21X1 U656 ( .A(n765), .B(n841), .C(n683), .Y(dataOut[1]) );
  OAI21X1 U658 ( .A(n765), .B(n823), .C(n659), .Y(dataOut[19]) );
  OAI21X1 U660 ( .A(n763), .B(n824), .C(n651), .Y(dataOut[18]) );
  OAI21X1 U662 ( .A(n764), .B(n825), .C(n668), .Y(dataOut[17]) );
  OAI21X1 U664 ( .A(n764), .B(n826), .C(n676), .Y(dataOut[16]) );
  OAI21X1 U666 ( .A(n763), .B(n827), .C(n660), .Y(dataOut[15]) );
  OAI21X1 U668 ( .A(n763), .B(n828), .C(n664), .Y(dataOut[14]) );
  OAI21X1 U670 ( .A(n763), .B(n829), .C(n669), .Y(dataOut[13]) );
  OAI21X1 U672 ( .A(n762), .B(n830), .C(n652), .Y(dataOut[12]) );
  OAI21X1 U674 ( .A(n762), .B(n831), .C(n656), .Y(dataOut[11]) );
  OAI21X1 U676 ( .A(n762), .B(n832), .C(n672), .Y(dataOut[10]) );
  OAI21X1 U678 ( .A(n762), .B(n842), .C(n679), .Y(dataOut[0]) );
  OAI21X1 U681 ( .A(inputBufferRequest[0]), .B(n148), .C(n2), .Y(n1046) );
  AOI22X1 U682 ( .A(n687), .B(n1043), .C(n755), .D(n1042), .Y(n1044) );
  OAI21X1 U684 ( .A(inputBufferRequest[1]), .B(n148), .C(n1), .Y(n1041) );
  AOI22X1 U685 ( .A(n1043), .B(n776), .C(n1042), .D(n777), .Y(n1040) );
  DFFSR priorityRegOdd_reg ( .D(n911), .CLK(clk), .R(n907), .S(1'b1), .Q(
        priorityRegOdd) );
  DFFSR priorityRegEven_reg ( .D(n910), .CLK(clk), .R(n907), .S(1'b1), .Q(
        priorityRegEven) );
  DFFSR oddBufferFull_reg ( .D(n909), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBufferFull) );
  DFFSR evenBufferFull_reg ( .D(n908), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBufferFull) );
  DFFSR oddBuffer_reg_63_ ( .D(n975), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[63]) );
  DFFSR oddBuffer_reg_62_ ( .D(n974), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[62]) );
  DFFSR oddBuffer_reg_61_ ( .D(n973), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[61]) );
  DFFSR oddBuffer_reg_60_ ( .D(n972), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[60]) );
  DFFSR oddBuffer_reg_59_ ( .D(n971), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[59]) );
  DFFSR oddBuffer_reg_58_ ( .D(n970), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[58]) );
  DFFSR oddBuffer_reg_57_ ( .D(n969), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[57]) );
  DFFSR oddBuffer_reg_56_ ( .D(n968), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[56]) );
  DFFSR oddBuffer_reg_55_ ( .D(n967), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[55]) );
  DFFSR oddBuffer_reg_54_ ( .D(n966), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[54]) );
  DFFSR oddBuffer_reg_53_ ( .D(n965), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[53]) );
  DFFSR oddBuffer_reg_52_ ( .D(n964), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[52]) );
  DFFSR oddBuffer_reg_10_ ( .D(n922), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[10]) );
  DFFSR oddBuffer_reg_9_ ( .D(n921), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[9]) );
  DFFSR oddBuffer_reg_8_ ( .D(n920), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[8]) );
  DFFSR oddBuffer_reg_7_ ( .D(n919), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[7]) );
  DFFSR oddBuffer_reg_6_ ( .D(n918), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[6]) );
  DFFSR oddBuffer_reg_5_ ( .D(n917), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[5]) );
  DFFSR oddBuffer_reg_4_ ( .D(n916), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[4]) );
  DFFSR oddBuffer_reg_3_ ( .D(n915), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[3]) );
  DFFSR oddBuffer_reg_1_ ( .D(n913), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[1]) );
  DFFSR oddBuffer_reg_0_ ( .D(n912), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[0]) );
  DFFSR oddBuffer_reg_2_ ( .D(n914), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[2]) );
  DFFSR oddBuffer_reg_24_ ( .D(n936), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[24]) );
  DFFSR oddBuffer_reg_23_ ( .D(n935), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[23]) );
  DFFSR oddBuffer_reg_22_ ( .D(n934), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[22]) );
  DFFSR oddBuffer_reg_21_ ( .D(n933), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[21]) );
  DFFSR oddBuffer_reg_20_ ( .D(n932), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[20]) );
  DFFSR oddBuffer_reg_19_ ( .D(n931), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[19]) );
  DFFSR oddBuffer_reg_18_ ( .D(n930), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[18]) );
  DFFSR oddBuffer_reg_17_ ( .D(n929), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[17]) );
  DFFSR oddBuffer_reg_16_ ( .D(n928), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[16]) );
  DFFSR oddBuffer_reg_15_ ( .D(n927), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[15]) );
  DFFSR oddBuffer_reg_14_ ( .D(n926), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[14]) );
  DFFSR oddBuffer_reg_13_ ( .D(n925), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[13]) );
  DFFSR oddBuffer_reg_12_ ( .D(n924), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[12]) );
  DFFSR oddBuffer_reg_11_ ( .D(n923), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[11]) );
  DFFSR oddBuffer_reg_25_ ( .D(n937), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[25]) );
  DFFSR evenBuffer_reg_63_ ( .D(n1039), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[63]) );
  DFFSR evenBuffer_reg_62_ ( .D(n1038), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[62]) );
  DFFSR evenBuffer_reg_61_ ( .D(n1037), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[61]) );
  DFFSR evenBuffer_reg_60_ ( .D(n1036), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[60]) );
  DFFSR evenBuffer_reg_59_ ( .D(n1035), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[59]) );
  DFFSR evenBuffer_reg_58_ ( .D(n1034), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[58]) );
  DFFSR evenBuffer_reg_57_ ( .D(n1033), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[57]) );
  DFFSR evenBuffer_reg_56_ ( .D(n1032), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[56]) );
  DFFSR evenBuffer_reg_55_ ( .D(n1031), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[55]) );
  DFFSR evenBuffer_reg_54_ ( .D(n1030), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[54]) );
  DFFSR evenBuffer_reg_53_ ( .D(n1029), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[53]) );
  DFFSR evenBuffer_reg_52_ ( .D(n1028), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[52]) );
  DFFSR oddBuffer_reg_47_ ( .D(n959), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[47]) );
  DFFSR oddBuffer_reg_46_ ( .D(n958), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[46]) );
  DFFSR oddBuffer_reg_45_ ( .D(n957), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[45]) );
  DFFSR oddBuffer_reg_44_ ( .D(n956), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[44]) );
  DFFSR oddBuffer_reg_43_ ( .D(n955), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[43]) );
  DFFSR oddBuffer_reg_42_ ( .D(n954), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[42]) );
  DFFSR oddBuffer_reg_41_ ( .D(n953), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[41]) );
  DFFSR oddBuffer_reg_40_ ( .D(n952), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[40]) );
  DFFSR oddBuffer_reg_39_ ( .D(n951), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[39]) );
  DFFSR oddBuffer_reg_38_ ( .D(n950), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[38]) );
  DFFSR oddBuffer_reg_37_ ( .D(n949), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[37]) );
  DFFSR oddBuffer_reg_36_ ( .D(n948), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[36]) );
  DFFSR oddBuffer_reg_35_ ( .D(n947), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[35]) );
  DFFSR oddBuffer_reg_34_ ( .D(n946), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[34]) );
  DFFSR oddBuffer_reg_33_ ( .D(n945), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[33]) );
  DFFSR oddBuffer_reg_32_ ( .D(n944), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[32]) );
  DFFSR oddBuffer_reg_31_ ( .D(n943), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[31]) );
  DFFSR oddBuffer_reg_30_ ( .D(n942), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[30]) );
  DFFSR oddBuffer_reg_28_ ( .D(n940), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[28]) );
  DFFSR oddBuffer_reg_26_ ( .D(n938), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[26]) );
  DFFSR oddBuffer_reg_29_ ( .D(n941), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[29]) );
  DFFSR oddBuffer_reg_27_ ( .D(n939), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[27]) );
  DFFSR oddBuffer_reg_51_ ( .D(n963), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[51]) );
  DFFSR oddBuffer_reg_50_ ( .D(n962), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[50]) );
  DFFSR oddBuffer_reg_49_ ( .D(n961), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[49]) );
  DFFSR oddBuffer_reg_48_ ( .D(n960), .CLK(clk), .R(n907), .S(1'b1), .Q(
        oddBuffer[48]) );
  DFFSR evenBuffer_reg_10_ ( .D(n986), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[10]) );
  DFFSR evenBuffer_reg_9_ ( .D(n985), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[9]) );
  DFFSR evenBuffer_reg_8_ ( .D(n984), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[8]) );
  DFFSR evenBuffer_reg_7_ ( .D(n983), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[7]) );
  DFFSR evenBuffer_reg_6_ ( .D(n982), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[6]) );
  DFFSR evenBuffer_reg_5_ ( .D(n981), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[5]) );
  DFFSR evenBuffer_reg_4_ ( .D(n980), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[4]) );
  DFFSR evenBuffer_reg_3_ ( .D(n979), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[3]) );
  DFFSR evenBuffer_reg_2_ ( .D(n978), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[2]) );
  DFFSR evenBuffer_reg_1_ ( .D(n977), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[1]) );
  DFFSR evenBuffer_reg_0_ ( .D(n976), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[0]) );
  DFFSR evenBuffer_reg_25_ ( .D(n1001), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[25]) );
  DFFSR evenBuffer_reg_24_ ( .D(n1000), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[24]) );
  DFFSR evenBuffer_reg_23_ ( .D(n999), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[23]) );
  DFFSR evenBuffer_reg_22_ ( .D(n998), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[22]) );
  DFFSR evenBuffer_reg_21_ ( .D(n997), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[21]) );
  DFFSR evenBuffer_reg_20_ ( .D(n996), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[20]) );
  DFFSR evenBuffer_reg_19_ ( .D(n995), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[19]) );
  DFFSR evenBuffer_reg_18_ ( .D(n994), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[18]) );
  DFFSR evenBuffer_reg_17_ ( .D(n993), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[17]) );
  DFFSR evenBuffer_reg_16_ ( .D(n992), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[16]) );
  DFFSR evenBuffer_reg_15_ ( .D(n991), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[15]) );
  DFFSR evenBuffer_reg_14_ ( .D(n990), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[14]) );
  DFFSR evenBuffer_reg_13_ ( .D(n989), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[13]) );
  DFFSR evenBuffer_reg_12_ ( .D(n988), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[12]) );
  DFFSR evenBuffer_reg_11_ ( .D(n987), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[11]) );
  DFFSR evenBuffer_reg_51_ ( .D(n1027), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[51]) );
  DFFSR evenBuffer_reg_50_ ( .D(n1026), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[50]) );
  DFFSR evenBuffer_reg_49_ ( .D(n1025), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[49]) );
  DFFSR evenBuffer_reg_48_ ( .D(n1024), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[48]) );
  DFFSR evenBuffer_reg_47_ ( .D(n1023), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[47]) );
  DFFSR evenBuffer_reg_46_ ( .D(n1022), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[46]) );
  DFFSR evenBuffer_reg_45_ ( .D(n1021), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[45]) );
  DFFSR evenBuffer_reg_44_ ( .D(n1020), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[44]) );
  DFFSR evenBuffer_reg_43_ ( .D(n1019), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[43]) );
  DFFSR evenBuffer_reg_42_ ( .D(n1018), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[42]) );
  DFFSR evenBuffer_reg_41_ ( .D(n1017), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[41]) );
  DFFSR evenBuffer_reg_40_ ( .D(n1016), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[40]) );
  DFFSR evenBuffer_reg_39_ ( .D(n1015), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[39]) );
  DFFSR evenBuffer_reg_38_ ( .D(n1014), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[38]) );
  DFFSR evenBuffer_reg_37_ ( .D(n1013), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[37]) );
  DFFSR evenBuffer_reg_36_ ( .D(n1012), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[36]) );
  DFFSR evenBuffer_reg_35_ ( .D(n1011), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[35]) );
  DFFSR evenBuffer_reg_34_ ( .D(n1010), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[34]) );
  DFFSR evenBuffer_reg_33_ ( .D(n1009), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[33]) );
  DFFSR evenBuffer_reg_32_ ( .D(n1008), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[32]) );
  DFFSR evenBuffer_reg_31_ ( .D(n1007), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[31]) );
  DFFSR evenBuffer_reg_30_ ( .D(n1006), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[30]) );
  DFFSR evenBuffer_reg_29_ ( .D(n1005), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[29]) );
  DFFSR evenBuffer_reg_28_ ( .D(n1004), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[28]) );
  DFFSR evenBuffer_reg_27_ ( .D(n1003), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[27]) );
  DFFSR evenBuffer_reg_26_ ( .D(n1002), .CLK(clk), .R(n907), .S(1'b1), .Q(
        evenBuffer[26]) );
  AND2X1 U2 ( .A(n767), .B(n680), .Y(n1111) );
  AND2X1 U3 ( .A(inputBufferRequest[1]), .B(n1046), .Y(InputBufferGrant[1]) );
  AND2X1 U4 ( .A(inputBufferRequest[0]), .B(n1041), .Y(InputBufferGrant[0]) );
  OR2X1 U5 ( .A(n753), .B(n151), .Y(n1185) );
  OR2X1 U6 ( .A(n753), .B(n150), .Y(n1184) );
  OR2X1 U7 ( .A(n754), .B(n151), .Y(n1255) );
  OR2X1 U8 ( .A(n150), .B(n754), .Y(n1254) );
  BUFX2 U9 ( .A(n1040), .Y(n1) );
  BUFX2 U10 ( .A(n1044), .Y(n2) );
  BUFX2 U11 ( .A(n1121), .Y(n3) );
  BUFX2 U12 ( .A(n1122), .Y(n4) );
  BUFX2 U13 ( .A(n1123), .Y(n5) );
  BUFX2 U14 ( .A(n1124), .Y(n6) );
  BUFX2 U15 ( .A(n1125), .Y(n7) );
  BUFX2 U16 ( .A(n1126), .Y(n8) );
  BUFX2 U17 ( .A(n1127), .Y(n9) );
  BUFX2 U18 ( .A(n1128), .Y(n10) );
  BUFX2 U19 ( .A(n1129), .Y(n11) );
  BUFX2 U20 ( .A(n1130), .Y(n12) );
  BUFX2 U21 ( .A(n1131), .Y(n13) );
  BUFX2 U22 ( .A(n1132), .Y(n14) );
  BUFX2 U23 ( .A(n1133), .Y(n15) );
  BUFX2 U24 ( .A(n1134), .Y(n16) );
  BUFX2 U25 ( .A(n1135), .Y(n17) );
  BUFX2 U26 ( .A(n1136), .Y(n18) );
  BUFX2 U27 ( .A(n1137), .Y(n19) );
  BUFX2 U28 ( .A(n1138), .Y(n20) );
  BUFX2 U29 ( .A(n1139), .Y(n21) );
  BUFX2 U30 ( .A(n1140), .Y(n22) );
  BUFX2 U31 ( .A(n1141), .Y(n23) );
  BUFX2 U32 ( .A(n1142), .Y(n24) );
  BUFX2 U33 ( .A(n1143), .Y(n25) );
  BUFX2 U34 ( .A(n1144), .Y(n26) );
  BUFX2 U35 ( .A(n1145), .Y(n27) );
  BUFX2 U36 ( .A(n1146), .Y(n28) );
  BUFX2 U37 ( .A(n1147), .Y(n29) );
  BUFX2 U38 ( .A(n1148), .Y(n30) );
  BUFX2 U39 ( .A(n1149), .Y(n31) );
  BUFX2 U40 ( .A(n1150), .Y(n32) );
  BUFX2 U41 ( .A(n1151), .Y(n33) );
  BUFX2 U42 ( .A(n1152), .Y(n34) );
  BUFX2 U43 ( .A(n1153), .Y(n35) );
  BUFX2 U44 ( .A(n1154), .Y(n36) );
  BUFX2 U45 ( .A(n1155), .Y(n37) );
  BUFX2 U46 ( .A(n1156), .Y(n38) );
  BUFX2 U47 ( .A(n1157), .Y(n39) );
  BUFX2 U48 ( .A(n1158), .Y(n40) );
  BUFX2 U49 ( .A(n1159), .Y(n41) );
  BUFX2 U50 ( .A(n1160), .Y(n42) );
  BUFX2 U51 ( .A(n1161), .Y(n43) );
  BUFX2 U52 ( .A(n1162), .Y(n44) );
  BUFX2 U53 ( .A(n1163), .Y(n45) );
  BUFX2 U54 ( .A(n1164), .Y(n46) );
  BUFX2 U55 ( .A(n1165), .Y(n47) );
  BUFX2 U56 ( .A(n1166), .Y(n48) );
  BUFX2 U57 ( .A(n1167), .Y(n49) );
  BUFX2 U58 ( .A(n1168), .Y(n50) );
  BUFX2 U59 ( .A(n1169), .Y(n51) );
  BUFX2 U60 ( .A(n1170), .Y(n52) );
  BUFX2 U61 ( .A(n1171), .Y(n53) );
  BUFX2 U62 ( .A(n1172), .Y(n54) );
  BUFX2 U63 ( .A(n1173), .Y(n55) );
  BUFX2 U64 ( .A(n1174), .Y(n56) );
  BUFX2 U65 ( .A(n1175), .Y(n57) );
  BUFX2 U66 ( .A(n1176), .Y(n58) );
  BUFX2 U67 ( .A(n1177), .Y(n59) );
  BUFX2 U68 ( .A(n1178), .Y(n60) );
  BUFX2 U69 ( .A(n1179), .Y(n61) );
  BUFX2 U70 ( .A(n1180), .Y(n62) );
  BUFX2 U71 ( .A(n1181), .Y(n63) );
  BUFX2 U72 ( .A(n1182), .Y(n64) );
  BUFX2 U73 ( .A(n1183), .Y(n65) );
  BUFX2 U74 ( .A(n1186), .Y(n66) );
  BUFX2 U75 ( .A(n1191), .Y(n67) );
  BUFX2 U76 ( .A(n1192), .Y(n68) );
  BUFX2 U77 ( .A(n1193), .Y(n69) );
  BUFX2 U78 ( .A(n1194), .Y(n70) );
  BUFX2 U79 ( .A(n1195), .Y(n71) );
  BUFX2 U80 ( .A(n1196), .Y(n72) );
  BUFX2 U81 ( .A(n1197), .Y(n73) );
  BUFX2 U82 ( .A(n1198), .Y(n74) );
  BUFX2 U83 ( .A(n1199), .Y(n75) );
  BUFX2 U84 ( .A(n1200), .Y(n76) );
  BUFX2 U85 ( .A(n1201), .Y(n77) );
  BUFX2 U86 ( .A(n1202), .Y(n78) );
  BUFX2 U87 ( .A(n1203), .Y(n79) );
  BUFX2 U88 ( .A(n1204), .Y(n80) );
  BUFX2 U89 ( .A(n1205), .Y(n81) );
  BUFX2 U90 ( .A(n1206), .Y(n82) );
  BUFX2 U91 ( .A(n1207), .Y(n83) );
  BUFX2 U92 ( .A(n1208), .Y(n84) );
  BUFX2 U93 ( .A(n1209), .Y(n85) );
  BUFX2 U94 ( .A(n1210), .Y(n86) );
  BUFX2 U95 ( .A(n1211), .Y(n87) );
  BUFX2 U96 ( .A(n1212), .Y(n88) );
  BUFX2 U97 ( .A(n1213), .Y(n89) );
  BUFX2 U98 ( .A(n1214), .Y(n90) );
  BUFX2 U99 ( .A(n1215), .Y(n91) );
  BUFX2 U100 ( .A(n1216), .Y(n92) );
  BUFX2 U101 ( .A(n1217), .Y(n93) );
  BUFX2 U102 ( .A(n1218), .Y(n94) );
  BUFX2 U103 ( .A(n1219), .Y(n95) );
  BUFX2 U104 ( .A(n1220), .Y(n96) );
  BUFX2 U105 ( .A(n1221), .Y(n97) );
  BUFX2 U106 ( .A(n1222), .Y(n98) );
  BUFX2 U107 ( .A(n1223), .Y(n99) );
  BUFX2 U108 ( .A(n1224), .Y(n100) );
  BUFX2 U109 ( .A(n1225), .Y(n101) );
  BUFX2 U110 ( .A(n1226), .Y(n102) );
  BUFX2 U111 ( .A(n1227), .Y(n103) );
  BUFX2 U112 ( .A(n1228), .Y(n104) );
  BUFX2 U113 ( .A(n1229), .Y(n105) );
  BUFX2 U114 ( .A(n1230), .Y(n106) );
  BUFX2 U115 ( .A(n1231), .Y(n107) );
  BUFX2 U116 ( .A(n1232), .Y(n108) );
  BUFX2 U117 ( .A(n1233), .Y(n109) );
  BUFX2 U118 ( .A(n1234), .Y(n110) );
  BUFX2 U119 ( .A(n1235), .Y(n111) );
  BUFX2 U120 ( .A(n1236), .Y(n112) );
  BUFX2 U121 ( .A(n1237), .Y(n113) );
  BUFX2 U122 ( .A(n1238), .Y(n114) );
  BUFX2 U123 ( .A(n1239), .Y(n115) );
  BUFX2 U124 ( .A(n1240), .Y(n116) );
  BUFX2 U125 ( .A(n1241), .Y(n117) );
  BUFX2 U126 ( .A(n1242), .Y(n118) );
  BUFX2 U127 ( .A(n1243), .Y(n119) );
  BUFX2 U128 ( .A(n1244), .Y(n120) );
  BUFX2 U129 ( .A(n1245), .Y(n121) );
  BUFX2 U130 ( .A(n1246), .Y(n122) );
  BUFX2 U131 ( .A(n1247), .Y(n123) );
  BUFX2 U132 ( .A(n1248), .Y(n124) );
  BUFX2 U133 ( .A(n1249), .Y(n125) );
  BUFX2 U134 ( .A(n1250), .Y(n126) );
  BUFX2 U135 ( .A(n1251), .Y(n127) );
  BUFX2 U136 ( .A(n1252), .Y(n128) );
  BUFX2 U137 ( .A(n1253), .Y(n129) );
  BUFX2 U138 ( .A(n1256), .Y(n130) );
  AND2X1 U139 ( .A(n727), .B(n768), .Y(n1064) );
  INVX1 U140 ( .A(n1064), .Y(n131) );
  AND2X1 U141 ( .A(n726), .B(n768), .Y(n1065) );
  INVX1 U142 ( .A(n1065), .Y(n132) );
  AND2X1 U143 ( .A(n725), .B(n768), .Y(n1066) );
  INVX1 U144 ( .A(n1066), .Y(n133) );
  AND2X1 U145 ( .A(n724), .B(n768), .Y(n1067) );
  INVX1 U146 ( .A(n1067), .Y(n134) );
  AND2X1 U147 ( .A(n723), .B(n768), .Y(n1068) );
  INVX1 U148 ( .A(n1068), .Y(n135) );
  AND2X1 U149 ( .A(n713), .B(n769), .Y(n1079) );
  INVX1 U150 ( .A(n1079), .Y(n136) );
  AND2X1 U151 ( .A(n712), .B(n769), .Y(n1081) );
  INVX1 U152 ( .A(n1081), .Y(n137) );
  AND2X1 U153 ( .A(n711), .B(n769), .Y(n1082) );
  INVX1 U154 ( .A(n1082), .Y(n138) );
  AND2X1 U155 ( .A(n710), .B(n769), .Y(n1083) );
  INVX1 U156 ( .A(n1083), .Y(n139) );
  AND2X1 U157 ( .A(n709), .B(n769), .Y(n1084) );
  INVX1 U158 ( .A(n1084), .Y(n140) );
  AND2X1 U159 ( .A(n697), .B(n770), .Y(n1097) );
  INVX1 U160 ( .A(n1097), .Y(n141) );
  AND2X1 U161 ( .A(n696), .B(n770), .Y(n1098) );
  INVX1 U162 ( .A(n1098), .Y(n142) );
  AND2X1 U163 ( .A(n695), .B(n770), .Y(n1099) );
  INVX1 U164 ( .A(n1099), .Y(n143) );
  AND2X1 U165 ( .A(n694), .B(n770), .Y(n1100) );
  INVX1 U166 ( .A(n1100), .Y(n144) );
  AND2X1 U167 ( .A(n693), .B(n770), .Y(n1101) );
  INVX1 U168 ( .A(n1101), .Y(n145) );
  AND2X1 U169 ( .A(sendOut), .B(n771), .Y(n1113) );
  INVX1 U170 ( .A(n1113), .Y(n146) );
  AND2X1 U171 ( .A(n767), .B(n149), .Y(n1114) );
  INVX1 U172 ( .A(n1114), .Y(n147) );
  OR2X1 U173 ( .A(n1042), .B(n1043), .Y(n1045) );
  INVX1 U174 ( .A(n1045), .Y(n148) );
  AND2X1 U175 ( .A(n151), .B(n150), .Y(n1116) );
  INVX1 U176 ( .A(n1116), .Y(n149) );
  INVX1 U177 ( .A(InputBufferGrant[0]), .Y(n150) );
  INVX1 U178 ( .A(InputBufferGrant[1]), .Y(n151) );
  INVX8 U179 ( .A(reset), .Y(n907) );
  AND2X1 U601 ( .A(n698), .B(n770), .Y(n1096) );
  INVX1 U603 ( .A(n1096), .Y(n634) );
  AND2X1 U605 ( .A(n714), .B(n769), .Y(n1078) );
  INVX1 U607 ( .A(n1078), .Y(n635) );
  AND2X1 U609 ( .A(n728), .B(n768), .Y(n1063) );
  INVX1 U611 ( .A(n1063), .Y(n636) );
  AND2X1 U613 ( .A(n689), .B(n771), .Y(n1106) );
  INVX1 U615 ( .A(n1106), .Y(n637) );
  AND2X1 U617 ( .A(n699), .B(n770), .Y(n1095) );
  INVX1 U619 ( .A(n1095), .Y(n638) );
  AND2X1 U621 ( .A(n716), .B(n769), .Y(n1076) );
  INVX1 U623 ( .A(n1076), .Y(n639) );
  AND2X1 U625 ( .A(n729), .B(n768), .Y(n1062) );
  INVX1 U627 ( .A(n1062), .Y(n640) );
  AND2X1 U629 ( .A(n690), .B(n771), .Y(n1105) );
  INVX1 U631 ( .A(n1105), .Y(n641) );
  AND2X1 U633 ( .A(n702), .B(n770), .Y(n1092) );
  INVX1 U635 ( .A(n1092), .Y(n642) );
  AND2X1 U637 ( .A(n718), .B(n769), .Y(n1074) );
  INVX1 U639 ( .A(n1074), .Y(n643) );
  AND2X1 U641 ( .A(n730), .B(n768), .Y(n1061) );
  INVX1 U643 ( .A(n1061), .Y(n644) );
  AND2X1 U645 ( .A(n691), .B(n771), .Y(n1104) );
  INVX1 U647 ( .A(n1104), .Y(n645) );
  AND2X1 U649 ( .A(n700), .B(n770), .Y(n1094) );
  INVX1 U651 ( .A(n1094), .Y(n646) );
  AND2X1 U653 ( .A(n719), .B(n769), .Y(n1073) );
  INVX1 U655 ( .A(n1073), .Y(n647) );
  AND2X1 U657 ( .A(n731), .B(n768), .Y(n1060) );
  INVX1 U659 ( .A(n1060), .Y(n648) );
  AND2X1 U661 ( .A(n701), .B(n770), .Y(n1093) );
  INVX1 U663 ( .A(n1093), .Y(n649) );
  AND2X1 U665 ( .A(n717), .B(n769), .Y(n1075) );
  INVX1 U667 ( .A(n1075), .Y(n650) );
  AND2X1 U669 ( .A(n734), .B(n768), .Y(n1056) );
  INVX1 U671 ( .A(n1056), .Y(n651) );
  AND2X1 U673 ( .A(n740), .B(n767), .Y(n1050) );
  INVX1 U675 ( .A(n1050), .Y(n652) );
  AND2X1 U677 ( .A(n692), .B(n771), .Y(n1103) );
  INVX1 U679 ( .A(n1103), .Y(n653) );
  AND2X1 U680 ( .A(n704), .B(n770), .Y(n1089) );
  INVX1 U683 ( .A(n1089), .Y(n654) );
  AND2X1 U686 ( .A(n721), .B(n769), .Y(n1071) );
  INVX1 U687 ( .A(n1071), .Y(n655) );
  AND2X1 U688 ( .A(n741), .B(n768), .Y(n1049) );
  INVX1 U689 ( .A(n1049), .Y(n656) );
  AND2X1 U690 ( .A(n703), .B(n770), .Y(n1090) );
  INVX1 U691 ( .A(n1090), .Y(n657) );
  AND2X1 U692 ( .A(n715), .B(n769), .Y(n1077) );
  INVX1 U693 ( .A(n1077), .Y(n658) );
  AND2X1 U694 ( .A(n733), .B(n768), .Y(n1057) );
  INVX1 U695 ( .A(n1057), .Y(n659) );
  AND2X1 U696 ( .A(n737), .B(n767), .Y(n1053) );
  INVX1 U697 ( .A(n1053), .Y(n660) );
  AND2X1 U698 ( .A(n743), .B(n771), .Y(n1110) );
  INVX1 U699 ( .A(n1110), .Y(n661) );
  AND2X1 U700 ( .A(n707), .B(n770), .Y(n1086) );
  INVX1 U701 ( .A(n1086), .Y(n662) );
  AND2X1 U702 ( .A(n722), .B(n769), .Y(n1070) );
  INVX1 U703 ( .A(n1070), .Y(n663) );
  AND2X1 U704 ( .A(n738), .B(n768), .Y(n1052) );
  INVX1 U705 ( .A(n1052), .Y(n664) );
  AND2X1 U706 ( .A(n744), .B(n771), .Y(n1109) );
  INVX1 U707 ( .A(n1109), .Y(n665) );
  AND2X1 U708 ( .A(n705), .B(n770), .Y(n1088) );
  INVX1 U709 ( .A(n1088), .Y(n666) );
  AND2X1 U710 ( .A(n720), .B(n769), .Y(n1072) );
  INVX1 U711 ( .A(n1072), .Y(n667) );
  AND2X1 U712 ( .A(n735), .B(n768), .Y(n1055) );
  INVX1 U713 ( .A(n1055), .Y(n668) );
  AND2X1 U714 ( .A(n739), .B(n767), .Y(n1051) );
  INVX1 U715 ( .A(n1051), .Y(n669) );
  AND2X1 U716 ( .A(n745), .B(n771), .Y(n1108) );
  INVX1 U717 ( .A(n1108), .Y(n670) );
  AND2X1 U718 ( .A(n732), .B(n769), .Y(n1059) );
  INVX1 U719 ( .A(n1059), .Y(n671) );
  AND2X1 U720 ( .A(n742), .B(n768), .Y(n1048) );
  INVX1 U721 ( .A(n1048), .Y(n672) );
  AND2X1 U722 ( .A(n746), .B(n771), .Y(n1107) );
  INVX1 U723 ( .A(n1107), .Y(n673) );
  AND2X1 U724 ( .A(n748), .B(n770), .Y(n1091) );
  INVX1 U725 ( .A(n1091), .Y(n674) );
  AND2X1 U726 ( .A(n708), .B(n770), .Y(n1085) );
  INVX1 U727 ( .A(n1085), .Y(n675) );
  AND2X1 U728 ( .A(n736), .B(n767), .Y(n1054) );
  INVX1 U729 ( .A(n1054), .Y(n676) );
  AND2X1 U730 ( .A(n747), .B(n771), .Y(n1102) );
  INVX1 U731 ( .A(n1102), .Y(n677) );
  AND2X1 U732 ( .A(n750), .B(n768), .Y(n1069) );
  INVX1 U733 ( .A(n1069), .Y(n678) );
  AND2X1 U734 ( .A(n752), .B(n769), .Y(n1047) );
  INVX1 U735 ( .A(n1047), .Y(n679) );
  BUFX2 U736 ( .A(evenBufferFull), .Y(n680) );
  AND2X1 U737 ( .A(n706), .B(n770), .Y(n1087) );
  INVX1 U738 ( .A(n1087), .Y(n681) );
  AND2X1 U739 ( .A(n749), .B(n769), .Y(n1080) );
  INVX1 U740 ( .A(n1080), .Y(n682) );
  AND2X1 U741 ( .A(n751), .B(n768), .Y(n1058) );
  INVX1 U742 ( .A(n1058), .Y(n683) );
  AND2X1 U743 ( .A(n774), .B(n771), .Y(n1119) );
  INVX1 U744 ( .A(n1119), .Y(n684) );
  AND2X1 U745 ( .A(readyOut), .B(n1112), .Y(sendOut) );
  INVX1 U746 ( .A(sendOut), .Y(n685) );
  INVX1 U747 ( .A(n1111), .Y(n686) );
  BUFX2 U748 ( .A(priorityRegEven), .Y(n687) );
  AND2X1 U749 ( .A(n774), .B(n773), .Y(n1118) );
  INVX1 U750 ( .A(n1118), .Y(n688) );
  BUFX2 U751 ( .A(evenBuffer[63]), .Y(n689) );
  BUFX2 U752 ( .A(evenBuffer[62]), .Y(n690) );
  BUFX2 U753 ( .A(evenBuffer[61]), .Y(n691) );
  BUFX2 U754 ( .A(evenBuffer[60]), .Y(n692) );
  BUFX2 U755 ( .A(evenBuffer[59]), .Y(n693) );
  BUFX2 U756 ( .A(evenBuffer[58]), .Y(n694) );
  BUFX2 U757 ( .A(evenBuffer[57]), .Y(n695) );
  BUFX2 U758 ( .A(evenBuffer[56]), .Y(n696) );
  BUFX2 U759 ( .A(evenBuffer[55]), .Y(n697) );
  BUFX2 U760 ( .A(evenBuffer[54]), .Y(n698) );
  BUFX2 U761 ( .A(evenBuffer[53]), .Y(n699) );
  BUFX2 U762 ( .A(evenBuffer[52]), .Y(n700) );
  BUFX2 U763 ( .A(evenBuffer[51]), .Y(n701) );
  BUFX2 U764 ( .A(evenBuffer[50]), .Y(n702) );
  BUFX2 U765 ( .A(evenBuffer[49]), .Y(n703) );
  BUFX2 U766 ( .A(evenBuffer[48]), .Y(n704) );
  BUFX2 U767 ( .A(evenBuffer[47]), .Y(n705) );
  BUFX2 U768 ( .A(evenBuffer[46]), .Y(n706) );
  BUFX2 U769 ( .A(evenBuffer[45]), .Y(n707) );
  BUFX2 U770 ( .A(evenBuffer[44]), .Y(n708) );
  BUFX2 U771 ( .A(evenBuffer[43]), .Y(n709) );
  BUFX2 U772 ( .A(evenBuffer[42]), .Y(n710) );
  BUFX2 U773 ( .A(evenBuffer[41]), .Y(n711) );
  BUFX2 U774 ( .A(evenBuffer[40]), .Y(n712) );
  BUFX2 U775 ( .A(evenBuffer[39]), .Y(n713) );
  BUFX2 U776 ( .A(evenBuffer[38]), .Y(n714) );
  BUFX2 U777 ( .A(evenBuffer[37]), .Y(n715) );
  BUFX2 U778 ( .A(evenBuffer[36]), .Y(n716) );
  BUFX2 U779 ( .A(evenBuffer[35]), .Y(n717) );
  BUFX2 U780 ( .A(evenBuffer[34]), .Y(n718) );
  BUFX2 U781 ( .A(evenBuffer[33]), .Y(n719) );
  BUFX2 U782 ( .A(evenBuffer[32]), .Y(n720) );
  BUFX2 U783 ( .A(evenBuffer[31]), .Y(n721) );
  BUFX2 U784 ( .A(evenBuffer[30]), .Y(n722) );
  BUFX2 U785 ( .A(evenBuffer[29]), .Y(n723) );
  BUFX2 U786 ( .A(evenBuffer[28]), .Y(n724) );
  BUFX2 U787 ( .A(evenBuffer[27]), .Y(n725) );
  BUFX2 U788 ( .A(evenBuffer[26]), .Y(n726) );
  BUFX2 U789 ( .A(evenBuffer[25]), .Y(n727) );
  BUFX2 U790 ( .A(evenBuffer[24]), .Y(n728) );
  BUFX2 U791 ( .A(evenBuffer[23]), .Y(n729) );
  BUFX2 U792 ( .A(evenBuffer[22]), .Y(n730) );
  BUFX2 U793 ( .A(evenBuffer[21]), .Y(n731) );
  BUFX2 U794 ( .A(evenBuffer[20]), .Y(n732) );
  BUFX2 U795 ( .A(evenBuffer[19]), .Y(n733) );
  BUFX2 U796 ( .A(evenBuffer[18]), .Y(n734) );
  BUFX2 U797 ( .A(evenBuffer[17]), .Y(n735) );
  BUFX2 U798 ( .A(evenBuffer[16]), .Y(n736) );
  BUFX2 U799 ( .A(evenBuffer[15]), .Y(n737) );
  BUFX2 U800 ( .A(evenBuffer[14]), .Y(n738) );
  BUFX2 U801 ( .A(evenBuffer[13]), .Y(n739) );
  BUFX2 U802 ( .A(evenBuffer[12]), .Y(n740) );
  BUFX2 U803 ( .A(evenBuffer[11]), .Y(n741) );
  BUFX2 U804 ( .A(evenBuffer[10]), .Y(n742) );
  BUFX2 U805 ( .A(evenBuffer[9]), .Y(n743) );
  BUFX2 U806 ( .A(evenBuffer[8]), .Y(n744) );
  BUFX2 U807 ( .A(evenBuffer[7]), .Y(n745) );
  BUFX2 U808 ( .A(evenBuffer[6]), .Y(n746) );
  BUFX2 U809 ( .A(evenBuffer[5]), .Y(n747) );
  BUFX2 U810 ( .A(evenBuffer[4]), .Y(n748) );
  BUFX2 U811 ( .A(evenBuffer[3]), .Y(n749) );
  BUFX2 U812 ( .A(evenBuffer[2]), .Y(n750) );
  BUFX2 U813 ( .A(evenBuffer[1]), .Y(n751) );
  BUFX2 U814 ( .A(evenBuffer[0]), .Y(n752) );
  AND2X1 U815 ( .A(n767), .B(n1187), .Y(n1120) );
  INVX1 U816 ( .A(n1120), .Y(n753) );
  AND2X1 U817 ( .A(n1257), .B(n772), .Y(n1189) );
  INVX1 U818 ( .A(n1189), .Y(n754) );
  BUFX2 U819 ( .A(priorityRegOdd), .Y(n755) );
  INVX1 U820 ( .A(n773), .Y(n768) );
  INVX1 U821 ( .A(n773), .Y(n769) );
  INVX1 U822 ( .A(n773), .Y(n767) );
  INVX1 U823 ( .A(n772), .Y(n766) );
  INVX1 U824 ( .A(n772), .Y(n765) );
  INVX1 U825 ( .A(n773), .Y(n764) );
  INVX1 U826 ( .A(n773), .Y(n762) );
  INVX1 U827 ( .A(n773), .Y(n763) );
  INVX1 U828 ( .A(n772), .Y(n771) );
  INVX1 U829 ( .A(n760), .Y(n772) );
  INVX1 U830 ( .A(n760), .Y(n773) );
  INVX1 U831 ( .A(n1254), .Y(n758) );
  INVX1 U832 ( .A(n1185), .Y(n757) );
  INVX1 U833 ( .A(n761), .Y(n760) );
  INVX1 U834 ( .A(n1184), .Y(n756) );
  INVX1 U835 ( .A(n1255), .Y(n759) );
  INVX1 U836 ( .A(n773), .Y(n770) );
  INVX1 U837 ( .A(polarity), .Y(n761) );
  INVX1 U838 ( .A(n1117), .Y(n774) );
  AND2X1 U839 ( .A(n771), .B(n778), .Y(n1042) );
  AND2X1 U840 ( .A(n775), .B(n773), .Y(n1043) );
  INVX1 U841 ( .A(n755), .Y(n777) );
  INVX1 U842 ( .A(n741), .Y(n895) );
  INVX1 U843 ( .A(n740), .Y(n894) );
  INVX1 U844 ( .A(n739), .Y(n893) );
  INVX1 U845 ( .A(n738), .Y(n892) );
  INVX1 U846 ( .A(n737), .Y(n891) );
  INVX1 U847 ( .A(n736), .Y(n890) );
  INVX1 U848 ( .A(n735), .Y(n889) );
  INVX1 U849 ( .A(n734), .Y(n888) );
  INVX1 U850 ( .A(n733), .Y(n887) );
  INVX1 U851 ( .A(n732), .Y(n886) );
  INVX1 U852 ( .A(n731), .Y(n885) );
  INVX1 U853 ( .A(n730), .Y(n884) );
  INVX1 U854 ( .A(n729), .Y(n883) );
  INVX1 U855 ( .A(n728), .Y(n882) );
  INVX1 U856 ( .A(n727), .Y(n881) );
  INVX1 U857 ( .A(n726), .Y(n880) );
  INVX1 U858 ( .A(n725), .Y(n879) );
  INVX1 U859 ( .A(n724), .Y(n878) );
  INVX1 U860 ( .A(n723), .Y(n877) );
  INVX1 U861 ( .A(n722), .Y(n876) );
  INVX1 U862 ( .A(n721), .Y(n875) );
  INVX1 U863 ( .A(n720), .Y(n874) );
  INVX1 U864 ( .A(n719), .Y(n873) );
  INVX1 U865 ( .A(n718), .Y(n872) );
  INVX1 U866 ( .A(n717), .Y(n871) );
  INVX1 U867 ( .A(n716), .Y(n870) );
  INVX1 U868 ( .A(n715), .Y(n869) );
  INVX1 U869 ( .A(n714), .Y(n868) );
  INVX1 U870 ( .A(n713), .Y(n867) );
  INVX1 U871 ( .A(n712), .Y(n866) );
  INVX1 U872 ( .A(n711), .Y(n865) );
  INVX1 U873 ( .A(n710), .Y(n864) );
  INVX1 U874 ( .A(n709), .Y(n863) );
  INVX1 U875 ( .A(n708), .Y(n862) );
  INVX1 U876 ( .A(n707), .Y(n861) );
  INVX1 U877 ( .A(n706), .Y(n860) );
  INVX1 U878 ( .A(n705), .Y(n859) );
  INVX1 U879 ( .A(n704), .Y(n858) );
  INVX1 U880 ( .A(n703), .Y(n857) );
  INVX1 U881 ( .A(n702), .Y(n856) );
  INVX1 U882 ( .A(n701), .Y(n855) );
  INVX1 U883 ( .A(n700), .Y(n854) );
  INVX1 U884 ( .A(n699), .Y(n853) );
  INVX1 U885 ( .A(n698), .Y(n852) );
  INVX1 U886 ( .A(n697), .Y(n851) );
  INVX1 U887 ( .A(n696), .Y(n850) );
  INVX1 U888 ( .A(n695), .Y(n849) );
  INVX1 U889 ( .A(n694), .Y(n848) );
  INVX1 U890 ( .A(n693), .Y(n847) );
  INVX1 U891 ( .A(n692), .Y(n846) );
  INVX1 U892 ( .A(n691), .Y(n845) );
  INVX1 U893 ( .A(n690), .Y(n844) );
  INVX1 U894 ( .A(n752), .Y(n906) );
  INVX1 U895 ( .A(n751), .Y(n905) );
  INVX1 U896 ( .A(n750), .Y(n904) );
  INVX1 U897 ( .A(n749), .Y(n903) );
  INVX1 U898 ( .A(n748), .Y(n902) );
  INVX1 U899 ( .A(n747), .Y(n901) );
  INVX1 U900 ( .A(n746), .Y(n900) );
  INVX1 U901 ( .A(n745), .Y(n899) );
  INVX1 U902 ( .A(n744), .Y(n898) );
  INVX1 U903 ( .A(n743), .Y(n897) );
  INVX1 U904 ( .A(n742), .Y(n896) );
  INVX1 U905 ( .A(n689), .Y(n843) );
  INVX1 U906 ( .A(n687), .Y(n776) );
  INVX1 U907 ( .A(n680), .Y(n775) );
  INVX1 U908 ( .A(oddBufferFull), .Y(n778) );
  INVX1 U909 ( .A(oddBuffer[0]), .Y(n842) );
  INVX1 U910 ( .A(oddBuffer[1]), .Y(n841) );
  INVX1 U911 ( .A(oddBuffer[2]), .Y(n840) );
  INVX1 U912 ( .A(oddBuffer[3]), .Y(n839) );
  INVX1 U913 ( .A(oddBuffer[4]), .Y(n838) );
  INVX1 U914 ( .A(oddBuffer[5]), .Y(n837) );
  INVX1 U915 ( .A(oddBuffer[6]), .Y(n836) );
  INVX1 U916 ( .A(oddBuffer[7]), .Y(n835) );
  INVX1 U917 ( .A(oddBuffer[8]), .Y(n834) );
  INVX1 U918 ( .A(oddBuffer[9]), .Y(n833) );
  INVX1 U919 ( .A(oddBuffer[10]), .Y(n832) );
  INVX1 U920 ( .A(oddBuffer[11]), .Y(n831) );
  INVX1 U921 ( .A(oddBuffer[12]), .Y(n830) );
  INVX1 U922 ( .A(oddBuffer[13]), .Y(n829) );
  INVX1 U923 ( .A(oddBuffer[14]), .Y(n828) );
  INVX1 U924 ( .A(oddBuffer[15]), .Y(n827) );
  INVX1 U925 ( .A(oddBuffer[16]), .Y(n826) );
  INVX1 U926 ( .A(oddBuffer[17]), .Y(n825) );
  INVX1 U927 ( .A(oddBuffer[18]), .Y(n824) );
  INVX1 U928 ( .A(oddBuffer[19]), .Y(n823) );
  INVX1 U929 ( .A(oddBuffer[20]), .Y(n822) );
  INVX1 U930 ( .A(oddBuffer[21]), .Y(n821) );
  INVX1 U931 ( .A(oddBuffer[22]), .Y(n820) );
  INVX1 U932 ( .A(oddBuffer[23]), .Y(n819) );
  INVX1 U933 ( .A(oddBuffer[24]), .Y(n818) );
  INVX1 U934 ( .A(oddBuffer[25]), .Y(n817) );
  INVX1 U935 ( .A(oddBuffer[26]), .Y(n816) );
  INVX1 U936 ( .A(oddBuffer[27]), .Y(n815) );
  INVX1 U937 ( .A(oddBuffer[28]), .Y(n814) );
  INVX1 U938 ( .A(oddBuffer[29]), .Y(n813) );
  INVX1 U939 ( .A(oddBuffer[30]), .Y(n812) );
  INVX1 U940 ( .A(oddBuffer[31]), .Y(n811) );
  INVX1 U941 ( .A(oddBuffer[32]), .Y(n810) );
  INVX1 U942 ( .A(oddBuffer[33]), .Y(n809) );
  INVX1 U943 ( .A(oddBuffer[34]), .Y(n808) );
  INVX1 U944 ( .A(oddBuffer[35]), .Y(n807) );
  INVX1 U945 ( .A(oddBuffer[36]), .Y(n806) );
  INVX1 U946 ( .A(oddBuffer[37]), .Y(n805) );
  INVX1 U947 ( .A(oddBuffer[38]), .Y(n804) );
  INVX1 U948 ( .A(oddBuffer[39]), .Y(n803) );
  INVX1 U949 ( .A(oddBuffer[40]), .Y(n802) );
  INVX1 U950 ( .A(oddBuffer[41]), .Y(n801) );
  INVX1 U951 ( .A(oddBuffer[42]), .Y(n800) );
  INVX1 U952 ( .A(oddBuffer[43]), .Y(n799) );
  INVX1 U953 ( .A(oddBuffer[44]), .Y(n798) );
  INVX1 U954 ( .A(oddBuffer[45]), .Y(n797) );
  INVX1 U955 ( .A(oddBuffer[46]), .Y(n796) );
  INVX1 U956 ( .A(oddBuffer[47]), .Y(n795) );
  INVX1 U957 ( .A(oddBuffer[48]), .Y(n794) );
  INVX1 U958 ( .A(oddBuffer[49]), .Y(n793) );
  INVX1 U959 ( .A(oddBuffer[50]), .Y(n792) );
  INVX1 U960 ( .A(oddBuffer[51]), .Y(n791) );
  INVX1 U961 ( .A(oddBuffer[52]), .Y(n790) );
  INVX1 U962 ( .A(oddBuffer[53]), .Y(n789) );
  INVX1 U963 ( .A(oddBuffer[54]), .Y(n788) );
  INVX1 U964 ( .A(oddBuffer[55]), .Y(n787) );
  INVX1 U965 ( .A(oddBuffer[56]), .Y(n786) );
  INVX1 U966 ( .A(oddBuffer[57]), .Y(n785) );
  INVX1 U967 ( .A(oddBuffer[58]), .Y(n784) );
  INVX1 U968 ( .A(oddBuffer[59]), .Y(n783) );
  INVX1 U969 ( .A(oddBuffer[60]), .Y(n782) );
  INVX1 U970 ( .A(oddBuffer[61]), .Y(n781) );
  INVX1 U971 ( .A(oddBuffer[62]), .Y(n780) );
  INVX1 U972 ( .A(oddBuffer[63]), .Y(n779) );
endmodule


module gold_router ( clk, reset, polarity, cwsi, cwri, ccwsi, ccwri, pesi, 
        peri, cwdi, ccwdi, pedi, cwso, cwro, ccwso, ccwro, peso, pero, cwdo, 
        ccwdo, pedo );
  input [63:0] cwdi;
  input [63:0] ccwdi;
  input [63:0] pedi;
  output [63:0] cwdo;
  output [63:0] ccwdo;
  output [63:0] pedo;
  input clk, reset, cwsi, ccwsi, pesi, cwro, ccwro, pero;
  output polarity, cwri, ccwri, peri, cwso, ccwso, peso;
  wire   n7, n5, n6;
  wire   [63:0] inBufferOut0;
  wire   [1:0] request0;
  wire   [1:0] grant2;
  wire   [1:0] grant0;
  wire   [63:0] inBufferOut1;
  wire   [1:0] request1;
  wire   [1:0] grant1;
  wire   [63:0] inBufferOut2;
  wire   [1:0] request2;

  DFFSR polarity_reg ( .D(n5), .CLK(clk), .R(n6), .S(1'b1), .Q(n7) );
  inputBuffer_1 i0 ( .clk(clk), .reset(reset), .polarity(polarity), .sendIn(
        cwsi), .readyIn(cwri), .dataIn(cwdi), .dataOut(inBufferOut0), 
        .request(request0), .outputBufferGrant({grant2[0], grant0[0]}) );
  inputBuffer_0 i1 ( .clk(clk), .reset(reset), .polarity(polarity), .sendIn(
        ccwsi), .readyIn(ccwri), .dataIn(ccwdi), .dataOut(inBufferOut1), 
        .request(request1), .outputBufferGrant({grant2[1], grant1[0]}) );
  inputBuffer_PE1 i2 ( .clk(clk), .reset(reset), .polarity(polarity), .sendIn(
        pesi), .readyIn(peri), .dataIn(pedi), .dataOut(inBufferOut2), 
        .request(request2), .outputBufferGrant({grant1[1], grant0[1]}) );
  outputBuffer_2 o1 ( .clk(clk), .reset(reset), .polarity(polarity), 
        .inputBufferRequest({request2[0], request0[0]}), .dataIn0(inBufferOut0), .dataIn1(inBufferOut2), .sendOut(cwso), .readyOut(cwro), .dataOut(cwdo), 
        .InputBufferGrant(grant0) );
  outputBuffer_1 o2 ( .clk(clk), .reset(reset), .polarity(polarity), 
        .inputBufferRequest({request2[1], request1[0]}), .dataIn0(inBufferOut1), .dataIn1(inBufferOut2), .sendOut(ccwso), .readyOut(ccwro), .dataOut(ccwdo), 
        .InputBufferGrant(grant1) );
  outputBuffer_0 o3 ( .clk(clk), .reset(reset), .polarity(polarity), 
        .inputBufferRequest({request1[1], request0[1]}), .dataIn0(inBufferOut0), .dataIn1(inBufferOut1), .sendOut(peso), .readyOut(pero), .dataOut(pedo), 
        .InputBufferGrant(grant2) );
  INVX1 U6 ( .A(n5), .Y(polarity) );
  INVX1 U7 ( .A(n7), .Y(n5) );
  INVX1 U8 ( .A(reset), .Y(n6) );
endmodule



module program_counter_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  AND2X1 U1 ( .A(n2), .B(A[15]), .Y(n1) );
  AND2X1 U2 ( .A(n3), .B(A[14]), .Y(n2) );
  AND2X1 U3 ( .A(n4), .B(A[13]), .Y(n3) );
  AND2X1 U4 ( .A(n5), .B(A[12]), .Y(n4) );
  AND2X1 U5 ( .A(n6), .B(A[11]), .Y(n5) );
  AND2X1 U6 ( .A(n7), .B(A[10]), .Y(n6) );
  AND2X1 U7 ( .A(n22), .B(A[9]), .Y(n7) );
  INVX1 U8 ( .A(A[2]), .Y(SUM[2]) );
  AND2X1 U9 ( .A(n9), .B(A[29]), .Y(n8) );
  AND2X1 U10 ( .A(n10), .B(A[28]), .Y(n9) );
  AND2X1 U11 ( .A(n11), .B(A[27]), .Y(n10) );
  AND2X1 U12 ( .A(n12), .B(A[26]), .Y(n11) );
  AND2X1 U13 ( .A(n13), .B(A[25]), .Y(n12) );
  AND2X1 U14 ( .A(n14), .B(A[24]), .Y(n13) );
  AND2X1 U15 ( .A(n15), .B(A[23]), .Y(n14) );
  AND2X1 U16 ( .A(n16), .B(A[22]), .Y(n15) );
  AND2X1 U17 ( .A(n17), .B(A[21]), .Y(n16) );
  AND2X1 U18 ( .A(n18), .B(A[20]), .Y(n17) );
  AND2X1 U19 ( .A(n19), .B(A[19]), .Y(n18) );
  AND2X1 U20 ( .A(n20), .B(A[18]), .Y(n19) );
  AND2X1 U21 ( .A(n21), .B(A[17]), .Y(n20) );
  AND2X1 U22 ( .A(n1), .B(A[16]), .Y(n21) );
  AND2X1 U23 ( .A(n23), .B(A[8]), .Y(n22) );
  AND2X1 U24 ( .A(n24), .B(A[7]), .Y(n23) );
  AND2X1 U25 ( .A(n25), .B(A[6]), .Y(n24) );
  AND2X1 U26 ( .A(n26), .B(A[5]), .Y(n25) );
  AND2X1 U27 ( .A(n27), .B(A[4]), .Y(n26) );
  AND2X1 U28 ( .A(A[2]), .B(A[3]), .Y(n27) );
  AND2X1 U29 ( .A(n8), .B(A[30]), .Y(n28) );
  XOR2X1 U30 ( .A(A[31]), .B(n28), .Y(SUM[31]) );
  XOR2X1 U31 ( .A(n8), .B(A[30]), .Y(SUM[30]) );
  XOR2X1 U32 ( .A(n9), .B(A[29]), .Y(SUM[29]) );
  XOR2X1 U33 ( .A(n10), .B(A[28]), .Y(SUM[28]) );
  XOR2X1 U34 ( .A(n11), .B(A[27]), .Y(SUM[27]) );
  XOR2X1 U35 ( .A(n12), .B(A[26]), .Y(SUM[26]) );
  XOR2X1 U36 ( .A(n13), .B(A[25]), .Y(SUM[25]) );
  XOR2X1 U37 ( .A(n14), .B(A[24]), .Y(SUM[24]) );
  XOR2X1 U38 ( .A(n15), .B(A[23]), .Y(SUM[23]) );
  XOR2X1 U39 ( .A(n16), .B(A[22]), .Y(SUM[22]) );
  XOR2X1 U40 ( .A(n17), .B(A[21]), .Y(SUM[21]) );
  XOR2X1 U41 ( .A(n18), .B(A[20]), .Y(SUM[20]) );
  XOR2X1 U42 ( .A(n19), .B(A[19]), .Y(SUM[19]) );
  XOR2X1 U43 ( .A(n20), .B(A[18]), .Y(SUM[18]) );
  XOR2X1 U44 ( .A(n21), .B(A[17]), .Y(SUM[17]) );
  XOR2X1 U45 ( .A(n1), .B(A[16]), .Y(SUM[16]) );
  XOR2X1 U46 ( .A(n2), .B(A[15]), .Y(SUM[15]) );
  XOR2X1 U47 ( .A(n3), .B(A[14]), .Y(SUM[14]) );
  XOR2X1 U48 ( .A(n4), .B(A[13]), .Y(SUM[13]) );
  XOR2X1 U49 ( .A(n5), .B(A[12]), .Y(SUM[12]) );
  XOR2X1 U50 ( .A(n6), .B(A[11]), .Y(SUM[11]) );
  XOR2X1 U51 ( .A(n7), .B(A[10]), .Y(SUM[10]) );
  XOR2X1 U52 ( .A(n22), .B(A[9]), .Y(SUM[9]) );
  XOR2X1 U53 ( .A(n23), .B(A[8]), .Y(SUM[8]) );
  XOR2X1 U54 ( .A(n24), .B(A[7]), .Y(SUM[7]) );
  XOR2X1 U55 ( .A(n25), .B(A[6]), .Y(SUM[6]) );
  XOR2X1 U56 ( .A(n26), .B(A[5]), .Y(SUM[5]) );
  XOR2X1 U57 ( .A(n27), .B(A[4]), .Y(SUM[4]) );
  XOR2X1 U58 ( .A(A[2]), .B(A[3]), .Y(SUM[3]) );
endmodule


module program_counter ( clk, reset, stall, pc_load, data_in, data_out );
  input [0:15] data_in;
  output [0:31] data_out;
  input clk, reset, stall, pc_load;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n1, n2, n3, n4, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204;

  DFFPOSX1 data_out_reg_31_ ( .D(n37), .CLK(clk), .Q(data_out[31]) );
  DFFPOSX1 data_out_reg_30_ ( .D(n40), .CLK(clk), .Q(data_out[30]) );
  DFFPOSX1 data_out_reg_29_ ( .D(n2), .CLK(clk), .Q(data_out[29]) );
  DFFPOSX1 data_out_reg_28_ ( .D(n44), .CLK(clk), .Q(data_out[28]) );
  DFFPOSX1 data_out_reg_27_ ( .D(n48), .CLK(clk), .Q(data_out[27]) );
  DFFPOSX1 data_out_reg_26_ ( .D(n52), .CLK(clk), .Q(data_out[26]) );
  DFFPOSX1 data_out_reg_25_ ( .D(n56), .CLK(clk), .Q(data_out[25]) );
  DFFPOSX1 data_out_reg_24_ ( .D(n60), .CLK(clk), .Q(data_out[24]) );
  DFFPOSX1 data_out_reg_23_ ( .D(n64), .CLK(clk), .Q(data_out[23]) );
  DFFPOSX1 data_out_reg_22_ ( .D(n68), .CLK(clk), .Q(data_out[22]) );
  DFFPOSX1 data_out_reg_21_ ( .D(n73), .CLK(clk), .Q(data_out[21]) );
  DFFPOSX1 data_out_reg_20_ ( .D(n78), .CLK(clk), .Q(data_out[20]) );
  DFFPOSX1 data_out_reg_19_ ( .D(n83), .CLK(clk), .Q(data_out[19]) );
  DFFPOSX1 data_out_reg_18_ ( .D(n87), .CLK(clk), .Q(data_out[18]) );
  DFFPOSX1 data_out_reg_17_ ( .D(n91), .CLK(clk), .Q(data_out[17]) );
  DFFPOSX1 data_out_reg_16_ ( .D(n95), .CLK(clk), .Q(data_out[16]) );
  DFFPOSX1 data_out_reg_15_ ( .D(n204), .CLK(clk), .Q(data_out[15]) );
  DFFPOSX1 data_out_reg_14_ ( .D(n203), .CLK(clk), .Q(data_out[14]) );
  DFFPOSX1 data_out_reg_13_ ( .D(n202), .CLK(clk), .Q(data_out[13]) );
  DFFPOSX1 data_out_reg_12_ ( .D(n201), .CLK(clk), .Q(data_out[12]) );
  DFFPOSX1 data_out_reg_11_ ( .D(n200), .CLK(clk), .Q(data_out[11]) );
  DFFPOSX1 data_out_reg_10_ ( .D(n199), .CLK(clk), .Q(data_out[10]) );
  DFFPOSX1 data_out_reg_9_ ( .D(n198), .CLK(clk), .Q(data_out[9]) );
  DFFPOSX1 data_out_reg_8_ ( .D(n197), .CLK(clk), .Q(data_out[8]) );
  DFFPOSX1 data_out_reg_7_ ( .D(n196), .CLK(clk), .Q(data_out[7]) );
  DFFPOSX1 data_out_reg_6_ ( .D(n195), .CLK(clk), .Q(data_out[6]) );
  DFFPOSX1 data_out_reg_5_ ( .D(n194), .CLK(clk), .Q(data_out[5]) );
  DFFPOSX1 data_out_reg_4_ ( .D(n193), .CLK(clk), .Q(data_out[4]) );
  DFFPOSX1 data_out_reg_3_ ( .D(n192), .CLK(clk), .Q(data_out[3]) );
  DFFPOSX1 data_out_reg_2_ ( .D(n175), .CLK(clk), .Q(data_out[2]) );
  DFFPOSX1 data_out_reg_1_ ( .D(n174), .CLK(clk), .Q(data_out[1]) );
  DFFPOSX1 data_out_reg_0_ ( .D(n173), .CLK(clk), .Q(data_out[0]) );
  program_counter_DW01_add_0 add_384 ( .A(data_out), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM({n36, n35, n34, n33, 
        n32, n31, n30, n29, n28, n27, n26, n25, n24, n23, n22, n21, n20, n19, 
        n18, n17, n16, n15, n14, n13, n12, n11, n10, n9, n8, n7, n6, n5}), 
        .CO() );
  AND2X1 U3 ( .A(n96), .B(n97), .Y(n176) );
  AND2X1 U4 ( .A(n92), .B(n93), .Y(n177) );
  AND2X1 U6 ( .A(n88), .B(n89), .Y(n178) );
  AND2X1 U7 ( .A(n84), .B(n85), .Y(n179) );
  AND2X1 U8 ( .A(n79), .B(n80), .Y(n180) );
  AND2X1 U9 ( .A(n74), .B(n75), .Y(n181) );
  AND2X1 U10 ( .A(n69), .B(n70), .Y(n182) );
  AND2X1 U11 ( .A(n65), .B(n66), .Y(n183) );
  AND2X1 U12 ( .A(n61), .B(n62), .Y(n184) );
  AND2X1 U13 ( .A(n57), .B(n58), .Y(n185) );
  AND2X1 U14 ( .A(n53), .B(n54), .Y(n186) );
  AND2X1 U15 ( .A(n49), .B(n50), .Y(n187) );
  AND2X1 U16 ( .A(n45), .B(n46), .Y(n188) );
  AND2X1 U17 ( .A(n3), .B(n4), .Y(n189) );
  AND2X1 U18 ( .A(n41), .B(n42), .Y(n190) );
  AND2X1 U19 ( .A(n38), .B(n39), .Y(n191) );
  AND2X1 U20 ( .A(stall), .B(n135), .Y(n138) );
  INVX1 U21 ( .A(n138), .Y(n1) );
  INVX1 U22 ( .A(n189), .Y(n2) );
  BUFX2 U23 ( .A(n166), .Y(n3) );
  AND2X1 U24 ( .A(n7), .B(n170), .Y(n165) );
  INVX1 U25 ( .A(n165), .Y(n4) );
  INVX1 U26 ( .A(n191), .Y(n37) );
  BUFX2 U27 ( .A(n172), .Y(n38) );
  AND2X1 U28 ( .A(n5), .B(n170), .Y(n171) );
  INVX1 U29 ( .A(n171), .Y(n39) );
  INVX1 U30 ( .A(n190), .Y(n40) );
  BUFX2 U31 ( .A(n168), .Y(n41) );
  AND2X1 U32 ( .A(n6), .B(n170), .Y(n167) );
  INVX1 U33 ( .A(n167), .Y(n42) );
  AND2X1 U34 ( .A(n21), .B(n170), .Y(n133) );
  INVX1 U35 ( .A(n133), .Y(n43) );
  INVX1 U36 ( .A(n188), .Y(n44) );
  BUFX2 U37 ( .A(n164), .Y(n45) );
  AND2X1 U38 ( .A(n8), .B(n170), .Y(n163) );
  INVX1 U39 ( .A(n163), .Y(n46) );
  AND2X1 U40 ( .A(n22), .B(n170), .Y(n131) );
  INVX1 U41 ( .A(n131), .Y(n47) );
  INVX1 U42 ( .A(n187), .Y(n48) );
  BUFX2 U43 ( .A(n162), .Y(n49) );
  AND2X1 U44 ( .A(n9), .B(n170), .Y(n161) );
  INVX1 U45 ( .A(n161), .Y(n50) );
  AND2X1 U46 ( .A(n23), .B(n170), .Y(n129) );
  INVX1 U47 ( .A(n129), .Y(n51) );
  INVX1 U48 ( .A(n186), .Y(n52) );
  BUFX2 U49 ( .A(n160), .Y(n53) );
  AND2X1 U50 ( .A(n10), .B(n170), .Y(n159) );
  INVX1 U51 ( .A(n159), .Y(n54) );
  AND2X1 U52 ( .A(n24), .B(n170), .Y(n127) );
  INVX1 U53 ( .A(n127), .Y(n55) );
  INVX1 U54 ( .A(n185), .Y(n56) );
  BUFX2 U55 ( .A(n158), .Y(n57) );
  AND2X1 U56 ( .A(n11), .B(n170), .Y(n157) );
  INVX1 U57 ( .A(n157), .Y(n58) );
  AND2X1 U58 ( .A(n25), .B(n170), .Y(n125) );
  INVX1 U59 ( .A(n125), .Y(n59) );
  INVX1 U60 ( .A(n184), .Y(n60) );
  BUFX2 U61 ( .A(n156), .Y(n61) );
  AND2X1 U62 ( .A(n12), .B(n170), .Y(n155) );
  INVX1 U63 ( .A(n155), .Y(n62) );
  AND2X1 U64 ( .A(n26), .B(n170), .Y(n123) );
  INVX1 U65 ( .A(n123), .Y(n63) );
  INVX1 U66 ( .A(n183), .Y(n64) );
  BUFX2 U67 ( .A(n154), .Y(n65) );
  AND2X1 U68 ( .A(n13), .B(n170), .Y(n153) );
  INVX1 U69 ( .A(n153), .Y(n66) );
  AND2X1 U70 ( .A(n27), .B(n170), .Y(n121) );
  INVX1 U71 ( .A(n121), .Y(n67) );
  INVX1 U72 ( .A(n182), .Y(n68) );
  BUFX2 U73 ( .A(n152), .Y(n69) );
  AND2X1 U74 ( .A(n14), .B(n170), .Y(n151) );
  INVX1 U75 ( .A(n151), .Y(n70) );
  AND2X1 U76 ( .A(n28), .B(n170), .Y(n119) );
  INVX1 U77 ( .A(n119), .Y(n71) );
  AND2X1 U78 ( .A(n31), .B(n170), .Y(n113) );
  INVX1 U79 ( .A(n113), .Y(n72) );
  INVX1 U80 ( .A(n181), .Y(n73) );
  BUFX2 U81 ( .A(n150), .Y(n74) );
  AND2X1 U82 ( .A(n15), .B(n170), .Y(n149) );
  INVX1 U83 ( .A(n149), .Y(n75) );
  AND2X1 U84 ( .A(n29), .B(n170), .Y(n117) );
  INVX1 U85 ( .A(n117), .Y(n76) );
  AND2X1 U86 ( .A(n32), .B(n170), .Y(n111) );
  INVX1 U87 ( .A(n111), .Y(n77) );
  INVX1 U88 ( .A(n180), .Y(n78) );
  BUFX2 U89 ( .A(n148), .Y(n79) );
  AND2X1 U90 ( .A(n16), .B(n170), .Y(n147) );
  INVX1 U91 ( .A(n147), .Y(n80) );
  AND2X1 U92 ( .A(n30), .B(n170), .Y(n115) );
  INVX1 U93 ( .A(n115), .Y(n81) );
  AND2X1 U94 ( .A(n33), .B(n170), .Y(n109) );
  INVX1 U95 ( .A(n109), .Y(n82) );
  INVX1 U96 ( .A(n179), .Y(n83) );
  BUFX2 U97 ( .A(n146), .Y(n84) );
  AND2X1 U98 ( .A(n17), .B(n170), .Y(n145) );
  INVX1 U99 ( .A(n145), .Y(n85) );
  AND2X1 U100 ( .A(n34), .B(n170), .Y(n107) );
  INVX1 U101 ( .A(n107), .Y(n86) );
  INVX1 U102 ( .A(n178), .Y(n87) );
  BUFX2 U103 ( .A(n144), .Y(n88) );
  AND2X1 U104 ( .A(n18), .B(n170), .Y(n143) );
  INVX1 U105 ( .A(n143), .Y(n89) );
  AND2X1 U106 ( .A(n35), .B(n170), .Y(n104) );
  INVX1 U107 ( .A(n104), .Y(n90) );
  INVX1 U108 ( .A(n177), .Y(n91) );
  BUFX2 U109 ( .A(n142), .Y(n92) );
  AND2X1 U110 ( .A(n19), .B(n170), .Y(n141) );
  INVX1 U111 ( .A(n141), .Y(n93) );
  AND2X1 U112 ( .A(n36), .B(n170), .Y(n102) );
  INVX1 U113 ( .A(n102), .Y(n94) );
  INVX1 U114 ( .A(n176), .Y(n95) );
  BUFX2 U115 ( .A(n140), .Y(n96) );
  AND2X1 U116 ( .A(n20), .B(n170), .Y(n139) );
  INVX1 U117 ( .A(n139), .Y(n97) );
  BUFX2 U118 ( .A(n1), .Y(n99) );
  BUFX2 U119 ( .A(n1), .Y(n98) );
  INVX1 U120 ( .A(stall), .Y(n136) );
  INVX1 U121 ( .A(n137), .Y(n169) );
  INVX1 U122 ( .A(n101), .Y(n170) );
  INVX1 U123 ( .A(pc_load), .Y(n100) );
  INVX1 U124 ( .A(data_out[0]), .Y(n103) );
  INVX1 U125 ( .A(data_out[1]), .Y(n106) );
  INVX1 U126 ( .A(data_out[2]), .Y(n108) );
  INVX1 U127 ( .A(data_out[3]), .Y(n110) );
  INVX1 U128 ( .A(data_out[4]), .Y(n112) );
  INVX1 U129 ( .A(data_out[5]), .Y(n114) );
  INVX1 U130 ( .A(data_out[6]), .Y(n116) );
  INVX1 U131 ( .A(data_out[7]), .Y(n118) );
  INVX1 U132 ( .A(data_out[8]), .Y(n120) );
  INVX1 U133 ( .A(data_out[9]), .Y(n122) );
  INVX1 U134 ( .A(data_out[10]), .Y(n124) );
  INVX1 U135 ( .A(data_out[11]), .Y(n126) );
  INVX1 U136 ( .A(data_out[12]), .Y(n128) );
  INVX1 U137 ( .A(data_out[13]), .Y(n130) );
  INVX1 U138 ( .A(data_out[14]), .Y(n132) );
  INVX1 U139 ( .A(data_out[15]), .Y(n134) );
  INVX1 U140 ( .A(reset), .Y(n135) );
  NAND3X1 U141 ( .A(n135), .B(n136), .C(n100), .Y(n101) );
  OAI21X1 U142 ( .A(n98), .B(n103), .C(n94), .Y(n173) );
  OAI21X1 U143 ( .A(n98), .B(n106), .C(n90), .Y(n174) );
  OAI21X1 U144 ( .A(n98), .B(n108), .C(n86), .Y(n175) );
  OAI21X1 U145 ( .A(n98), .B(n110), .C(n82), .Y(n192) );
  OAI21X1 U146 ( .A(n98), .B(n112), .C(n77), .Y(n193) );
  OAI21X1 U147 ( .A(n98), .B(n114), .C(n72), .Y(n194) );
  OAI21X1 U148 ( .A(n99), .B(n116), .C(n81), .Y(n195) );
  OAI21X1 U149 ( .A(n99), .B(n118), .C(n76), .Y(n196) );
  OAI21X1 U150 ( .A(n99), .B(n120), .C(n71), .Y(n197) );
  OAI21X1 U151 ( .A(n99), .B(n122), .C(n67), .Y(n198) );
  OAI21X1 U152 ( .A(n99), .B(n124), .C(n63), .Y(n199) );
  OAI21X1 U153 ( .A(n99), .B(n126), .C(n59), .Y(n200) );
  OAI21X1 U154 ( .A(n99), .B(n128), .C(n55), .Y(n201) );
  OAI21X1 U155 ( .A(n99), .B(n130), .C(n51), .Y(n202) );
  OAI21X1 U156 ( .A(n99), .B(n132), .C(n47), .Y(n203) );
  OAI21X1 U157 ( .A(n99), .B(n134), .C(n43), .Y(n204) );
  NAND3X1 U158 ( .A(pc_load), .B(n136), .C(n135), .Y(n137) );
  AOI22X1 U159 ( .A(data_in[0]), .B(n169), .C(data_out[16]), .D(n138), .Y(n140) );
  AOI22X1 U160 ( .A(data_in[1]), .B(n169), .C(data_out[17]), .D(n138), .Y(n142) );
  AOI22X1 U161 ( .A(data_in[2]), .B(n169), .C(data_out[18]), .D(n138), .Y(n144) );
  AOI22X1 U162 ( .A(data_in[3]), .B(n169), .C(data_out[19]), .D(n138), .Y(n146) );
  AOI22X1 U163 ( .A(data_in[4]), .B(n169), .C(data_out[20]), .D(n138), .Y(n148) );
  AOI22X1 U164 ( .A(data_in[5]), .B(n169), .C(data_out[21]), .D(n138), .Y(n150) );
  AOI22X1 U165 ( .A(data_in[6]), .B(n169), .C(data_out[22]), .D(n138), .Y(n152) );
  AOI22X1 U166 ( .A(data_in[7]), .B(n169), .C(data_out[23]), .D(n138), .Y(n154) );
  AOI22X1 U167 ( .A(data_in[8]), .B(n169), .C(data_out[24]), .D(n138), .Y(n156) );
  AOI22X1 U168 ( .A(data_in[9]), .B(n169), .C(data_out[25]), .D(n138), .Y(n158) );
  AOI22X1 U169 ( .A(data_in[10]), .B(n169), .C(data_out[26]), .D(n138), .Y(
        n160) );
  AOI22X1 U170 ( .A(data_in[11]), .B(n169), .C(data_out[27]), .D(n138), .Y(
        n162) );
  AOI22X1 U171 ( .A(data_in[12]), .B(n169), .C(data_out[28]), .D(n138), .Y(
        n164) );
  AOI22X1 U172 ( .A(data_in[13]), .B(n169), .C(data_out[29]), .D(n138), .Y(
        n166) );
  AOI22X1 U173 ( .A(data_in[14]), .B(n169), .C(data_out[30]), .D(n138), .Y(
        n168) );
  AOI22X1 U174 ( .A(data_in[15]), .B(n169), .C(data_out[31]), .D(n138), .Y(
        n172) );
endmodule


module register_file ( clk, reset, write_en, read1_addr, read2_addr, 
        write_addr, Din, Dout1, Dout2, PPP );
  input [0:4] read1_addr;
  input [0:4] read2_addr;
  input [0:4] write_addr;
  input [0:63] Din;
  output [0:63] Dout1;
  output [0:63] Dout2;
  input [0:2] PPP;
  input clk, reset, write_en;
  wire   n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n2517, n2584, n2651,
         n2718, n2785, n2852, n2919, n2986, n4508, n4576, n4577, n4578, n4579,
         n4580, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n120, n121, n122, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229;
  wire   [2047:0] ram;
  wire   [0:63] current_ram;

  DFFPOSX1 ram_reg_0__0_ ( .D(n6716), .CLK(clk), .Q(ram[2047]) );
  DFFPOSX1 ram_reg_0__1_ ( .D(n6715), .CLK(clk), .Q(ram[2046]) );
  DFFPOSX1 ram_reg_0__2_ ( .D(n6714), .CLK(clk), .Q(ram[2045]) );
  DFFPOSX1 ram_reg_0__3_ ( .D(n6713), .CLK(clk), .Q(ram[2044]) );
  DFFPOSX1 ram_reg_0__4_ ( .D(n6712), .CLK(clk), .Q(ram[2043]) );
  DFFPOSX1 ram_reg_0__5_ ( .D(n6711), .CLK(clk), .Q(ram[2042]) );
  DFFPOSX1 ram_reg_0__6_ ( .D(n6710), .CLK(clk), .Q(ram[2041]) );
  DFFPOSX1 ram_reg_0__7_ ( .D(n6709), .CLK(clk), .Q(ram[2040]) );
  DFFPOSX1 ram_reg_0__8_ ( .D(n6708), .CLK(clk), .Q(ram[2039]) );
  DFFPOSX1 ram_reg_0__9_ ( .D(n6707), .CLK(clk), .Q(ram[2038]) );
  DFFPOSX1 ram_reg_0__10_ ( .D(n6706), .CLK(clk), .Q(ram[2037]) );
  DFFPOSX1 ram_reg_0__11_ ( .D(n6705), .CLK(clk), .Q(ram[2036]) );
  DFFPOSX1 ram_reg_0__12_ ( .D(n6704), .CLK(clk), .Q(ram[2035]) );
  DFFPOSX1 ram_reg_0__13_ ( .D(n6703), .CLK(clk), .Q(ram[2034]) );
  DFFPOSX1 ram_reg_0__14_ ( .D(n6702), .CLK(clk), .Q(ram[2033]) );
  DFFPOSX1 ram_reg_0__15_ ( .D(n6701), .CLK(clk), .Q(ram[2032]) );
  DFFPOSX1 ram_reg_0__16_ ( .D(n6700), .CLK(clk), .Q(ram[2031]) );
  DFFPOSX1 ram_reg_0__17_ ( .D(n6699), .CLK(clk), .Q(ram[2030]) );
  DFFPOSX1 ram_reg_0__18_ ( .D(n6698), .CLK(clk), .Q(ram[2029]) );
  DFFPOSX1 ram_reg_0__19_ ( .D(n6697), .CLK(clk), .Q(ram[2028]) );
  DFFPOSX1 ram_reg_0__20_ ( .D(n6696), .CLK(clk), .Q(ram[2027]) );
  DFFPOSX1 ram_reg_0__21_ ( .D(n6695), .CLK(clk), .Q(ram[2026]) );
  DFFPOSX1 ram_reg_0__22_ ( .D(n6694), .CLK(clk), .Q(ram[2025]) );
  DFFPOSX1 ram_reg_0__23_ ( .D(n6693), .CLK(clk), .Q(ram[2024]) );
  DFFPOSX1 ram_reg_0__24_ ( .D(n6692), .CLK(clk), .Q(ram[2023]) );
  DFFPOSX1 ram_reg_0__25_ ( .D(n6691), .CLK(clk), .Q(ram[2022]) );
  DFFPOSX1 ram_reg_0__26_ ( .D(n6690), .CLK(clk), .Q(ram[2021]) );
  DFFPOSX1 ram_reg_0__27_ ( .D(n6689), .CLK(clk), .Q(ram[2020]) );
  DFFPOSX1 ram_reg_0__28_ ( .D(n6688), .CLK(clk), .Q(ram[2019]) );
  DFFPOSX1 ram_reg_0__29_ ( .D(n6687), .CLK(clk), .Q(ram[2018]) );
  DFFPOSX1 ram_reg_0__30_ ( .D(n6686), .CLK(clk), .Q(ram[2017]) );
  DFFPOSX1 ram_reg_0__31_ ( .D(n6685), .CLK(clk), .Q(ram[2016]) );
  DFFPOSX1 ram_reg_0__32_ ( .D(n6684), .CLK(clk), .Q(ram[2015]) );
  DFFPOSX1 ram_reg_0__33_ ( .D(n6683), .CLK(clk), .Q(ram[2014]) );
  DFFPOSX1 ram_reg_0__34_ ( .D(n6682), .CLK(clk), .Q(ram[2013]) );
  DFFPOSX1 ram_reg_0__35_ ( .D(n6681), .CLK(clk), .Q(ram[2012]) );
  DFFPOSX1 ram_reg_0__36_ ( .D(n6680), .CLK(clk), .Q(ram[2011]) );
  DFFPOSX1 ram_reg_0__37_ ( .D(n6679), .CLK(clk), .Q(ram[2010]) );
  DFFPOSX1 ram_reg_0__38_ ( .D(n6678), .CLK(clk), .Q(ram[2009]) );
  DFFPOSX1 ram_reg_0__39_ ( .D(n6677), .CLK(clk), .Q(ram[2008]) );
  DFFPOSX1 ram_reg_0__40_ ( .D(n6676), .CLK(clk), .Q(ram[2007]) );
  DFFPOSX1 ram_reg_0__41_ ( .D(n6675), .CLK(clk), .Q(ram[2006]) );
  DFFPOSX1 ram_reg_0__42_ ( .D(n6674), .CLK(clk), .Q(ram[2005]) );
  DFFPOSX1 ram_reg_0__43_ ( .D(n6673), .CLK(clk), .Q(ram[2004]) );
  DFFPOSX1 ram_reg_0__44_ ( .D(n6672), .CLK(clk), .Q(ram[2003]) );
  DFFPOSX1 ram_reg_0__45_ ( .D(n6671), .CLK(clk), .Q(ram[2002]) );
  DFFPOSX1 ram_reg_0__46_ ( .D(n6670), .CLK(clk), .Q(ram[2001]) );
  DFFPOSX1 ram_reg_0__47_ ( .D(n6669), .CLK(clk), .Q(ram[2000]) );
  DFFPOSX1 ram_reg_0__48_ ( .D(n6668), .CLK(clk), .Q(ram[1999]) );
  DFFPOSX1 ram_reg_0__49_ ( .D(n6667), .CLK(clk), .Q(ram[1998]) );
  DFFPOSX1 ram_reg_0__50_ ( .D(n6666), .CLK(clk), .Q(ram[1997]) );
  DFFPOSX1 ram_reg_0__51_ ( .D(n6665), .CLK(clk), .Q(ram[1996]) );
  DFFPOSX1 ram_reg_0__52_ ( .D(n6664), .CLK(clk), .Q(ram[1995]) );
  DFFPOSX1 ram_reg_0__53_ ( .D(n6663), .CLK(clk), .Q(ram[1994]) );
  DFFPOSX1 ram_reg_0__54_ ( .D(n6662), .CLK(clk), .Q(ram[1993]) );
  DFFPOSX1 ram_reg_0__55_ ( .D(n6661), .CLK(clk), .Q(ram[1992]) );
  DFFPOSX1 ram_reg_0__56_ ( .D(n6660), .CLK(clk), .Q(ram[1991]) );
  DFFPOSX1 ram_reg_0__57_ ( .D(n6659), .CLK(clk), .Q(ram[1990]) );
  DFFPOSX1 ram_reg_0__58_ ( .D(n6658), .CLK(clk), .Q(ram[1989]) );
  DFFPOSX1 ram_reg_0__59_ ( .D(n6657), .CLK(clk), .Q(ram[1988]) );
  DFFPOSX1 ram_reg_0__60_ ( .D(n6656), .CLK(clk), .Q(ram[1987]) );
  DFFPOSX1 ram_reg_0__61_ ( .D(n6655), .CLK(clk), .Q(ram[1986]) );
  DFFPOSX1 ram_reg_0__62_ ( .D(n6654), .CLK(clk), .Q(ram[1985]) );
  DFFPOSX1 ram_reg_0__63_ ( .D(n6653), .CLK(clk), .Q(ram[1984]) );
  DFFPOSX1 ram_reg_1__0_ ( .D(n6652), .CLK(clk), .Q(ram[1983]) );
  DFFPOSX1 ram_reg_1__1_ ( .D(n6651), .CLK(clk), .Q(ram[1982]) );
  DFFPOSX1 ram_reg_1__2_ ( .D(n6650), .CLK(clk), .Q(ram[1981]) );
  DFFPOSX1 ram_reg_1__3_ ( .D(n6649), .CLK(clk), .Q(ram[1980]) );
  DFFPOSX1 ram_reg_1__4_ ( .D(n6648), .CLK(clk), .Q(ram[1979]) );
  DFFPOSX1 ram_reg_1__5_ ( .D(n6647), .CLK(clk), .Q(ram[1978]) );
  DFFPOSX1 ram_reg_1__6_ ( .D(n6646), .CLK(clk), .Q(ram[1977]) );
  DFFPOSX1 ram_reg_1__7_ ( .D(n6645), .CLK(clk), .Q(ram[1976]) );
  DFFPOSX1 ram_reg_1__8_ ( .D(n6644), .CLK(clk), .Q(ram[1975]) );
  DFFPOSX1 ram_reg_1__9_ ( .D(n6643), .CLK(clk), .Q(ram[1974]) );
  DFFPOSX1 ram_reg_1__10_ ( .D(n6642), .CLK(clk), .Q(ram[1973]) );
  DFFPOSX1 ram_reg_1__11_ ( .D(n6641), .CLK(clk), .Q(ram[1972]) );
  DFFPOSX1 ram_reg_1__12_ ( .D(n6640), .CLK(clk), .Q(ram[1971]) );
  DFFPOSX1 ram_reg_1__13_ ( .D(n6639), .CLK(clk), .Q(ram[1970]) );
  DFFPOSX1 ram_reg_1__14_ ( .D(n6638), .CLK(clk), .Q(ram[1969]) );
  DFFPOSX1 ram_reg_1__15_ ( .D(n6637), .CLK(clk), .Q(ram[1968]) );
  DFFPOSX1 ram_reg_1__16_ ( .D(n6636), .CLK(clk), .Q(ram[1967]) );
  DFFPOSX1 ram_reg_1__17_ ( .D(n6635), .CLK(clk), .Q(ram[1966]) );
  DFFPOSX1 ram_reg_1__18_ ( .D(n6634), .CLK(clk), .Q(ram[1965]) );
  DFFPOSX1 ram_reg_1__19_ ( .D(n6633), .CLK(clk), .Q(ram[1964]) );
  DFFPOSX1 ram_reg_1__20_ ( .D(n6632), .CLK(clk), .Q(ram[1963]) );
  DFFPOSX1 ram_reg_1__21_ ( .D(n6631), .CLK(clk), .Q(ram[1962]) );
  DFFPOSX1 ram_reg_1__22_ ( .D(n6630), .CLK(clk), .Q(ram[1961]) );
  DFFPOSX1 ram_reg_1__23_ ( .D(n6629), .CLK(clk), .Q(ram[1960]) );
  DFFPOSX1 ram_reg_1__24_ ( .D(n6628), .CLK(clk), .Q(ram[1959]) );
  DFFPOSX1 ram_reg_1__25_ ( .D(n6627), .CLK(clk), .Q(ram[1958]) );
  DFFPOSX1 ram_reg_1__26_ ( .D(n6626), .CLK(clk), .Q(ram[1957]) );
  DFFPOSX1 ram_reg_1__27_ ( .D(n6625), .CLK(clk), .Q(ram[1956]) );
  DFFPOSX1 ram_reg_1__28_ ( .D(n6624), .CLK(clk), .Q(ram[1955]) );
  DFFPOSX1 ram_reg_1__29_ ( .D(n6623), .CLK(clk), .Q(ram[1954]) );
  DFFPOSX1 ram_reg_1__30_ ( .D(n6622), .CLK(clk), .Q(ram[1953]) );
  DFFPOSX1 ram_reg_1__31_ ( .D(n6621), .CLK(clk), .Q(ram[1952]) );
  DFFPOSX1 ram_reg_1__32_ ( .D(n6620), .CLK(clk), .Q(ram[1951]) );
  DFFPOSX1 ram_reg_1__33_ ( .D(n6619), .CLK(clk), .Q(ram[1950]) );
  DFFPOSX1 ram_reg_1__34_ ( .D(n6618), .CLK(clk), .Q(ram[1949]) );
  DFFPOSX1 ram_reg_1__35_ ( .D(n6617), .CLK(clk), .Q(ram[1948]) );
  DFFPOSX1 ram_reg_1__36_ ( .D(n6616), .CLK(clk), .Q(ram[1947]) );
  DFFPOSX1 ram_reg_1__37_ ( .D(n6615), .CLK(clk), .Q(ram[1946]) );
  DFFPOSX1 ram_reg_1__38_ ( .D(n6614), .CLK(clk), .Q(ram[1945]) );
  DFFPOSX1 ram_reg_1__39_ ( .D(n6613), .CLK(clk), .Q(ram[1944]) );
  DFFPOSX1 ram_reg_1__40_ ( .D(n6612), .CLK(clk), .Q(ram[1943]) );
  DFFPOSX1 ram_reg_1__41_ ( .D(n6611), .CLK(clk), .Q(ram[1942]) );
  DFFPOSX1 ram_reg_1__42_ ( .D(n6610), .CLK(clk), .Q(ram[1941]) );
  DFFPOSX1 ram_reg_1__43_ ( .D(n6609), .CLK(clk), .Q(ram[1940]) );
  DFFPOSX1 ram_reg_1__44_ ( .D(n6608), .CLK(clk), .Q(ram[1939]) );
  DFFPOSX1 ram_reg_1__45_ ( .D(n6607), .CLK(clk), .Q(ram[1938]) );
  DFFPOSX1 ram_reg_1__46_ ( .D(n6606), .CLK(clk), .Q(ram[1937]) );
  DFFPOSX1 ram_reg_1__47_ ( .D(n6605), .CLK(clk), .Q(ram[1936]) );
  DFFPOSX1 ram_reg_1__48_ ( .D(n6604), .CLK(clk), .Q(ram[1935]) );
  DFFPOSX1 ram_reg_1__49_ ( .D(n6603), .CLK(clk), .Q(ram[1934]) );
  DFFPOSX1 ram_reg_1__50_ ( .D(n6602), .CLK(clk), .Q(ram[1933]) );
  DFFPOSX1 ram_reg_1__51_ ( .D(n6601), .CLK(clk), .Q(ram[1932]) );
  DFFPOSX1 ram_reg_1__52_ ( .D(n6600), .CLK(clk), .Q(ram[1931]) );
  DFFPOSX1 ram_reg_1__53_ ( .D(n6599), .CLK(clk), .Q(ram[1930]) );
  DFFPOSX1 ram_reg_1__54_ ( .D(n6598), .CLK(clk), .Q(ram[1929]) );
  DFFPOSX1 ram_reg_1__55_ ( .D(n6597), .CLK(clk), .Q(ram[1928]) );
  DFFPOSX1 ram_reg_1__56_ ( .D(n6596), .CLK(clk), .Q(ram[1927]) );
  DFFPOSX1 ram_reg_1__57_ ( .D(n6595), .CLK(clk), .Q(ram[1926]) );
  DFFPOSX1 ram_reg_1__58_ ( .D(n6594), .CLK(clk), .Q(ram[1925]) );
  DFFPOSX1 ram_reg_1__59_ ( .D(n6593), .CLK(clk), .Q(ram[1924]) );
  DFFPOSX1 ram_reg_1__60_ ( .D(n6592), .CLK(clk), .Q(ram[1923]) );
  DFFPOSX1 ram_reg_1__61_ ( .D(n6591), .CLK(clk), .Q(ram[1922]) );
  DFFPOSX1 ram_reg_1__62_ ( .D(n6590), .CLK(clk), .Q(ram[1921]) );
  DFFPOSX1 ram_reg_1__63_ ( .D(n6589), .CLK(clk), .Q(ram[1920]) );
  DFFPOSX1 ram_reg_2__0_ ( .D(n6588), .CLK(clk), .Q(ram[1919]) );
  DFFPOSX1 ram_reg_2__1_ ( .D(n6587), .CLK(clk), .Q(ram[1918]) );
  DFFPOSX1 ram_reg_2__2_ ( .D(n6586), .CLK(clk), .Q(ram[1917]) );
  DFFPOSX1 ram_reg_2__3_ ( .D(n6585), .CLK(clk), .Q(ram[1916]) );
  DFFPOSX1 ram_reg_2__4_ ( .D(n6584), .CLK(clk), .Q(ram[1915]) );
  DFFPOSX1 ram_reg_2__5_ ( .D(n6583), .CLK(clk), .Q(ram[1914]) );
  DFFPOSX1 ram_reg_2__6_ ( .D(n6582), .CLK(clk), .Q(ram[1913]) );
  DFFPOSX1 ram_reg_2__7_ ( .D(n6581), .CLK(clk), .Q(ram[1912]) );
  DFFPOSX1 ram_reg_2__8_ ( .D(n6580), .CLK(clk), .Q(ram[1911]) );
  DFFPOSX1 ram_reg_2__9_ ( .D(n6579), .CLK(clk), .Q(ram[1910]) );
  DFFPOSX1 ram_reg_2__10_ ( .D(n6578), .CLK(clk), .Q(ram[1909]) );
  DFFPOSX1 ram_reg_2__11_ ( .D(n6577), .CLK(clk), .Q(ram[1908]) );
  DFFPOSX1 ram_reg_2__12_ ( .D(n6576), .CLK(clk), .Q(ram[1907]) );
  DFFPOSX1 ram_reg_2__13_ ( .D(n6575), .CLK(clk), .Q(ram[1906]) );
  DFFPOSX1 ram_reg_2__14_ ( .D(n6574), .CLK(clk), .Q(ram[1905]) );
  DFFPOSX1 ram_reg_2__15_ ( .D(n6573), .CLK(clk), .Q(ram[1904]) );
  DFFPOSX1 ram_reg_2__16_ ( .D(n6572), .CLK(clk), .Q(ram[1903]) );
  DFFPOSX1 ram_reg_2__17_ ( .D(n6571), .CLK(clk), .Q(ram[1902]) );
  DFFPOSX1 ram_reg_2__18_ ( .D(n6570), .CLK(clk), .Q(ram[1901]) );
  DFFPOSX1 ram_reg_2__19_ ( .D(n6569), .CLK(clk), .Q(ram[1900]) );
  DFFPOSX1 ram_reg_2__20_ ( .D(n6568), .CLK(clk), .Q(ram[1899]) );
  DFFPOSX1 ram_reg_2__21_ ( .D(n6567), .CLK(clk), .Q(ram[1898]) );
  DFFPOSX1 ram_reg_2__22_ ( .D(n6566), .CLK(clk), .Q(ram[1897]) );
  DFFPOSX1 ram_reg_2__23_ ( .D(n6565), .CLK(clk), .Q(ram[1896]) );
  DFFPOSX1 ram_reg_2__24_ ( .D(n6564), .CLK(clk), .Q(ram[1895]) );
  DFFPOSX1 ram_reg_2__25_ ( .D(n6563), .CLK(clk), .Q(ram[1894]) );
  DFFPOSX1 ram_reg_2__26_ ( .D(n6562), .CLK(clk), .Q(ram[1893]) );
  DFFPOSX1 ram_reg_2__27_ ( .D(n6561), .CLK(clk), .Q(ram[1892]) );
  DFFPOSX1 ram_reg_2__28_ ( .D(n6560), .CLK(clk), .Q(ram[1891]) );
  DFFPOSX1 ram_reg_2__29_ ( .D(n6559), .CLK(clk), .Q(ram[1890]) );
  DFFPOSX1 ram_reg_2__30_ ( .D(n6558), .CLK(clk), .Q(ram[1889]) );
  DFFPOSX1 ram_reg_2__31_ ( .D(n6557), .CLK(clk), .Q(ram[1888]) );
  DFFPOSX1 ram_reg_2__32_ ( .D(n6556), .CLK(clk), .Q(ram[1887]) );
  DFFPOSX1 ram_reg_2__33_ ( .D(n6555), .CLK(clk), .Q(ram[1886]) );
  DFFPOSX1 ram_reg_2__34_ ( .D(n6554), .CLK(clk), .Q(ram[1885]) );
  DFFPOSX1 ram_reg_2__35_ ( .D(n6553), .CLK(clk), .Q(ram[1884]) );
  DFFPOSX1 ram_reg_2__36_ ( .D(n6552), .CLK(clk), .Q(ram[1883]) );
  DFFPOSX1 ram_reg_2__37_ ( .D(n6551), .CLK(clk), .Q(ram[1882]) );
  DFFPOSX1 ram_reg_2__38_ ( .D(n6550), .CLK(clk), .Q(ram[1881]) );
  DFFPOSX1 ram_reg_2__39_ ( .D(n6549), .CLK(clk), .Q(ram[1880]) );
  DFFPOSX1 ram_reg_2__40_ ( .D(n6548), .CLK(clk), .Q(ram[1879]) );
  DFFPOSX1 ram_reg_2__41_ ( .D(n6547), .CLK(clk), .Q(ram[1878]) );
  DFFPOSX1 ram_reg_2__42_ ( .D(n6546), .CLK(clk), .Q(ram[1877]) );
  DFFPOSX1 ram_reg_2__43_ ( .D(n6545), .CLK(clk), .Q(ram[1876]) );
  DFFPOSX1 ram_reg_2__44_ ( .D(n6544), .CLK(clk), .Q(ram[1875]) );
  DFFPOSX1 ram_reg_2__45_ ( .D(n6543), .CLK(clk), .Q(ram[1874]) );
  DFFPOSX1 ram_reg_2__46_ ( .D(n6542), .CLK(clk), .Q(ram[1873]) );
  DFFPOSX1 ram_reg_2__47_ ( .D(n6541), .CLK(clk), .Q(ram[1872]) );
  DFFPOSX1 ram_reg_2__48_ ( .D(n6540), .CLK(clk), .Q(ram[1871]) );
  DFFPOSX1 ram_reg_2__49_ ( .D(n6539), .CLK(clk), .Q(ram[1870]) );
  DFFPOSX1 ram_reg_2__50_ ( .D(n6538), .CLK(clk), .Q(ram[1869]) );
  DFFPOSX1 ram_reg_2__51_ ( .D(n6537), .CLK(clk), .Q(ram[1868]) );
  DFFPOSX1 ram_reg_2__52_ ( .D(n6536), .CLK(clk), .Q(ram[1867]) );
  DFFPOSX1 ram_reg_2__53_ ( .D(n6535), .CLK(clk), .Q(ram[1866]) );
  DFFPOSX1 ram_reg_2__54_ ( .D(n6534), .CLK(clk), .Q(ram[1865]) );
  DFFPOSX1 ram_reg_2__55_ ( .D(n6533), .CLK(clk), .Q(ram[1864]) );
  DFFPOSX1 ram_reg_2__56_ ( .D(n6532), .CLK(clk), .Q(ram[1863]) );
  DFFPOSX1 ram_reg_2__57_ ( .D(n6531), .CLK(clk), .Q(ram[1862]) );
  DFFPOSX1 ram_reg_2__58_ ( .D(n6530), .CLK(clk), .Q(ram[1861]) );
  DFFPOSX1 ram_reg_2__59_ ( .D(n6529), .CLK(clk), .Q(ram[1860]) );
  DFFPOSX1 ram_reg_2__60_ ( .D(n6528), .CLK(clk), .Q(ram[1859]) );
  DFFPOSX1 ram_reg_2__61_ ( .D(n6527), .CLK(clk), .Q(ram[1858]) );
  DFFPOSX1 ram_reg_2__62_ ( .D(n6526), .CLK(clk), .Q(ram[1857]) );
  DFFPOSX1 ram_reg_2__63_ ( .D(n6525), .CLK(clk), .Q(ram[1856]) );
  DFFPOSX1 ram_reg_3__0_ ( .D(n6524), .CLK(clk), .Q(ram[1855]) );
  DFFPOSX1 ram_reg_3__1_ ( .D(n6523), .CLK(clk), .Q(ram[1854]) );
  DFFPOSX1 ram_reg_3__2_ ( .D(n6522), .CLK(clk), .Q(ram[1853]) );
  DFFPOSX1 ram_reg_3__3_ ( .D(n6521), .CLK(clk), .Q(ram[1852]) );
  DFFPOSX1 ram_reg_3__4_ ( .D(n6520), .CLK(clk), .Q(ram[1851]) );
  DFFPOSX1 ram_reg_3__5_ ( .D(n6519), .CLK(clk), .Q(ram[1850]) );
  DFFPOSX1 ram_reg_3__6_ ( .D(n6518), .CLK(clk), .Q(ram[1849]) );
  DFFPOSX1 ram_reg_3__7_ ( .D(n6517), .CLK(clk), .Q(ram[1848]) );
  DFFPOSX1 ram_reg_3__8_ ( .D(n6516), .CLK(clk), .Q(ram[1847]) );
  DFFPOSX1 ram_reg_3__9_ ( .D(n6515), .CLK(clk), .Q(ram[1846]) );
  DFFPOSX1 ram_reg_3__10_ ( .D(n6514), .CLK(clk), .Q(ram[1845]) );
  DFFPOSX1 ram_reg_3__11_ ( .D(n6513), .CLK(clk), .Q(ram[1844]) );
  DFFPOSX1 ram_reg_3__12_ ( .D(n6512), .CLK(clk), .Q(ram[1843]) );
  DFFPOSX1 ram_reg_3__13_ ( .D(n6511), .CLK(clk), .Q(ram[1842]) );
  DFFPOSX1 ram_reg_3__14_ ( .D(n6510), .CLK(clk), .Q(ram[1841]) );
  DFFPOSX1 ram_reg_3__15_ ( .D(n6509), .CLK(clk), .Q(ram[1840]) );
  DFFPOSX1 ram_reg_3__16_ ( .D(n6508), .CLK(clk), .Q(ram[1839]) );
  DFFPOSX1 ram_reg_3__17_ ( .D(n6507), .CLK(clk), .Q(ram[1838]) );
  DFFPOSX1 ram_reg_3__18_ ( .D(n6506), .CLK(clk), .Q(ram[1837]) );
  DFFPOSX1 ram_reg_3__19_ ( .D(n6505), .CLK(clk), .Q(ram[1836]) );
  DFFPOSX1 ram_reg_3__20_ ( .D(n6504), .CLK(clk), .Q(ram[1835]) );
  DFFPOSX1 ram_reg_3__21_ ( .D(n6503), .CLK(clk), .Q(ram[1834]) );
  DFFPOSX1 ram_reg_3__22_ ( .D(n6502), .CLK(clk), .Q(ram[1833]) );
  DFFPOSX1 ram_reg_3__23_ ( .D(n6501), .CLK(clk), .Q(ram[1832]) );
  DFFPOSX1 ram_reg_3__24_ ( .D(n6500), .CLK(clk), .Q(ram[1831]) );
  DFFPOSX1 ram_reg_3__25_ ( .D(n6499), .CLK(clk), .Q(ram[1830]) );
  DFFPOSX1 ram_reg_3__26_ ( .D(n6498), .CLK(clk), .Q(ram[1829]) );
  DFFPOSX1 ram_reg_3__27_ ( .D(n6497), .CLK(clk), .Q(ram[1828]) );
  DFFPOSX1 ram_reg_3__28_ ( .D(n6496), .CLK(clk), .Q(ram[1827]) );
  DFFPOSX1 ram_reg_3__29_ ( .D(n6495), .CLK(clk), .Q(ram[1826]) );
  DFFPOSX1 ram_reg_3__30_ ( .D(n6494), .CLK(clk), .Q(ram[1825]) );
  DFFPOSX1 ram_reg_3__31_ ( .D(n6493), .CLK(clk), .Q(ram[1824]) );
  DFFPOSX1 ram_reg_3__32_ ( .D(n6492), .CLK(clk), .Q(ram[1823]) );
  DFFPOSX1 ram_reg_3__33_ ( .D(n6491), .CLK(clk), .Q(ram[1822]) );
  DFFPOSX1 ram_reg_3__34_ ( .D(n6490), .CLK(clk), .Q(ram[1821]) );
  DFFPOSX1 ram_reg_3__35_ ( .D(n6489), .CLK(clk), .Q(ram[1820]) );
  DFFPOSX1 ram_reg_3__36_ ( .D(n6488), .CLK(clk), .Q(ram[1819]) );
  DFFPOSX1 ram_reg_3__37_ ( .D(n6487), .CLK(clk), .Q(ram[1818]) );
  DFFPOSX1 ram_reg_3__38_ ( .D(n6486), .CLK(clk), .Q(ram[1817]) );
  DFFPOSX1 ram_reg_3__39_ ( .D(n6485), .CLK(clk), .Q(ram[1816]) );
  DFFPOSX1 ram_reg_3__40_ ( .D(n6484), .CLK(clk), .Q(ram[1815]) );
  DFFPOSX1 ram_reg_3__41_ ( .D(n6483), .CLK(clk), .Q(ram[1814]) );
  DFFPOSX1 ram_reg_3__42_ ( .D(n6482), .CLK(clk), .Q(ram[1813]) );
  DFFPOSX1 ram_reg_3__43_ ( .D(n6481), .CLK(clk), .Q(ram[1812]) );
  DFFPOSX1 ram_reg_3__44_ ( .D(n6480), .CLK(clk), .Q(ram[1811]) );
  DFFPOSX1 ram_reg_3__45_ ( .D(n6479), .CLK(clk), .Q(ram[1810]) );
  DFFPOSX1 ram_reg_3__46_ ( .D(n6478), .CLK(clk), .Q(ram[1809]) );
  DFFPOSX1 ram_reg_3__47_ ( .D(n6477), .CLK(clk), .Q(ram[1808]) );
  DFFPOSX1 ram_reg_3__48_ ( .D(n6476), .CLK(clk), .Q(ram[1807]) );
  DFFPOSX1 ram_reg_3__49_ ( .D(n6475), .CLK(clk), .Q(ram[1806]) );
  DFFPOSX1 ram_reg_3__50_ ( .D(n6474), .CLK(clk), .Q(ram[1805]) );
  DFFPOSX1 ram_reg_3__51_ ( .D(n6473), .CLK(clk), .Q(ram[1804]) );
  DFFPOSX1 ram_reg_3__52_ ( .D(n6472), .CLK(clk), .Q(ram[1803]) );
  DFFPOSX1 ram_reg_3__53_ ( .D(n6471), .CLK(clk), .Q(ram[1802]) );
  DFFPOSX1 ram_reg_3__54_ ( .D(n6470), .CLK(clk), .Q(ram[1801]) );
  DFFPOSX1 ram_reg_3__55_ ( .D(n6469), .CLK(clk), .Q(ram[1800]) );
  DFFPOSX1 ram_reg_3__56_ ( .D(n6468), .CLK(clk), .Q(ram[1799]) );
  DFFPOSX1 ram_reg_3__57_ ( .D(n6467), .CLK(clk), .Q(ram[1798]) );
  DFFPOSX1 ram_reg_3__58_ ( .D(n6466), .CLK(clk), .Q(ram[1797]) );
  DFFPOSX1 ram_reg_3__59_ ( .D(n6465), .CLK(clk), .Q(ram[1796]) );
  DFFPOSX1 ram_reg_3__60_ ( .D(n6464), .CLK(clk), .Q(ram[1795]) );
  DFFPOSX1 ram_reg_3__61_ ( .D(n6463), .CLK(clk), .Q(ram[1794]) );
  DFFPOSX1 ram_reg_3__62_ ( .D(n6462), .CLK(clk), .Q(ram[1793]) );
  DFFPOSX1 ram_reg_3__63_ ( .D(n6461), .CLK(clk), .Q(ram[1792]) );
  DFFPOSX1 ram_reg_4__0_ ( .D(n6460), .CLK(clk), .Q(ram[1791]) );
  DFFPOSX1 ram_reg_4__1_ ( .D(n6459), .CLK(clk), .Q(ram[1790]) );
  DFFPOSX1 ram_reg_4__2_ ( .D(n6458), .CLK(clk), .Q(ram[1789]) );
  DFFPOSX1 ram_reg_4__3_ ( .D(n6457), .CLK(clk), .Q(ram[1788]) );
  DFFPOSX1 ram_reg_4__4_ ( .D(n6456), .CLK(clk), .Q(ram[1787]) );
  DFFPOSX1 ram_reg_4__5_ ( .D(n6455), .CLK(clk), .Q(ram[1786]) );
  DFFPOSX1 ram_reg_4__6_ ( .D(n6454), .CLK(clk), .Q(ram[1785]) );
  DFFPOSX1 ram_reg_4__7_ ( .D(n6453), .CLK(clk), .Q(ram[1784]) );
  DFFPOSX1 ram_reg_4__8_ ( .D(n6452), .CLK(clk), .Q(ram[1783]) );
  DFFPOSX1 ram_reg_4__9_ ( .D(n6451), .CLK(clk), .Q(ram[1782]) );
  DFFPOSX1 ram_reg_4__10_ ( .D(n6450), .CLK(clk), .Q(ram[1781]) );
  DFFPOSX1 ram_reg_4__11_ ( .D(n6449), .CLK(clk), .Q(ram[1780]) );
  DFFPOSX1 ram_reg_4__12_ ( .D(n6448), .CLK(clk), .Q(ram[1779]) );
  DFFPOSX1 ram_reg_4__13_ ( .D(n6447), .CLK(clk), .Q(ram[1778]) );
  DFFPOSX1 ram_reg_4__14_ ( .D(n6446), .CLK(clk), .Q(ram[1777]) );
  DFFPOSX1 ram_reg_4__15_ ( .D(n6445), .CLK(clk), .Q(ram[1776]) );
  DFFPOSX1 ram_reg_4__16_ ( .D(n6444), .CLK(clk), .Q(ram[1775]) );
  DFFPOSX1 ram_reg_4__17_ ( .D(n6443), .CLK(clk), .Q(ram[1774]) );
  DFFPOSX1 ram_reg_4__18_ ( .D(n6442), .CLK(clk), .Q(ram[1773]) );
  DFFPOSX1 ram_reg_4__19_ ( .D(n6441), .CLK(clk), .Q(ram[1772]) );
  DFFPOSX1 ram_reg_4__20_ ( .D(n6440), .CLK(clk), .Q(ram[1771]) );
  DFFPOSX1 ram_reg_4__21_ ( .D(n6439), .CLK(clk), .Q(ram[1770]) );
  DFFPOSX1 ram_reg_4__22_ ( .D(n6438), .CLK(clk), .Q(ram[1769]) );
  DFFPOSX1 ram_reg_4__23_ ( .D(n6437), .CLK(clk), .Q(ram[1768]) );
  DFFPOSX1 ram_reg_4__24_ ( .D(n6436), .CLK(clk), .Q(ram[1767]) );
  DFFPOSX1 ram_reg_4__25_ ( .D(n6435), .CLK(clk), .Q(ram[1766]) );
  DFFPOSX1 ram_reg_4__26_ ( .D(n6434), .CLK(clk), .Q(ram[1765]) );
  DFFPOSX1 ram_reg_4__27_ ( .D(n6433), .CLK(clk), .Q(ram[1764]) );
  DFFPOSX1 ram_reg_4__28_ ( .D(n6432), .CLK(clk), .Q(ram[1763]) );
  DFFPOSX1 ram_reg_4__29_ ( .D(n6431), .CLK(clk), .Q(ram[1762]) );
  DFFPOSX1 ram_reg_4__30_ ( .D(n6430), .CLK(clk), .Q(ram[1761]) );
  DFFPOSX1 ram_reg_4__31_ ( .D(n6429), .CLK(clk), .Q(ram[1760]) );
  DFFPOSX1 ram_reg_4__32_ ( .D(n6428), .CLK(clk), .Q(ram[1759]) );
  DFFPOSX1 ram_reg_4__33_ ( .D(n6427), .CLK(clk), .Q(ram[1758]) );
  DFFPOSX1 ram_reg_4__34_ ( .D(n6426), .CLK(clk), .Q(ram[1757]) );
  DFFPOSX1 ram_reg_4__35_ ( .D(n6425), .CLK(clk), .Q(ram[1756]) );
  DFFPOSX1 ram_reg_4__36_ ( .D(n6424), .CLK(clk), .Q(ram[1755]) );
  DFFPOSX1 ram_reg_4__37_ ( .D(n6423), .CLK(clk), .Q(ram[1754]) );
  DFFPOSX1 ram_reg_4__38_ ( .D(n6422), .CLK(clk), .Q(ram[1753]) );
  DFFPOSX1 ram_reg_4__39_ ( .D(n6421), .CLK(clk), .Q(ram[1752]) );
  DFFPOSX1 ram_reg_4__40_ ( .D(n6420), .CLK(clk), .Q(ram[1751]) );
  DFFPOSX1 ram_reg_4__41_ ( .D(n6419), .CLK(clk), .Q(ram[1750]) );
  DFFPOSX1 ram_reg_4__42_ ( .D(n6418), .CLK(clk), .Q(ram[1749]) );
  DFFPOSX1 ram_reg_4__43_ ( .D(n6417), .CLK(clk), .Q(ram[1748]) );
  DFFPOSX1 ram_reg_4__44_ ( .D(n6416), .CLK(clk), .Q(ram[1747]) );
  DFFPOSX1 ram_reg_4__45_ ( .D(n6415), .CLK(clk), .Q(ram[1746]) );
  DFFPOSX1 ram_reg_4__46_ ( .D(n6414), .CLK(clk), .Q(ram[1745]) );
  DFFPOSX1 ram_reg_4__47_ ( .D(n6413), .CLK(clk), .Q(ram[1744]) );
  DFFPOSX1 ram_reg_4__48_ ( .D(n6412), .CLK(clk), .Q(ram[1743]) );
  DFFPOSX1 ram_reg_4__49_ ( .D(n6411), .CLK(clk), .Q(ram[1742]) );
  DFFPOSX1 ram_reg_4__50_ ( .D(n6410), .CLK(clk), .Q(ram[1741]) );
  DFFPOSX1 ram_reg_4__51_ ( .D(n6409), .CLK(clk), .Q(ram[1740]) );
  DFFPOSX1 ram_reg_4__52_ ( .D(n6408), .CLK(clk), .Q(ram[1739]) );
  DFFPOSX1 ram_reg_4__53_ ( .D(n6407), .CLK(clk), .Q(ram[1738]) );
  DFFPOSX1 ram_reg_4__54_ ( .D(n6406), .CLK(clk), .Q(ram[1737]) );
  DFFPOSX1 ram_reg_4__55_ ( .D(n6405), .CLK(clk), .Q(ram[1736]) );
  DFFPOSX1 ram_reg_4__56_ ( .D(n6404), .CLK(clk), .Q(ram[1735]) );
  DFFPOSX1 ram_reg_4__57_ ( .D(n6403), .CLK(clk), .Q(ram[1734]) );
  DFFPOSX1 ram_reg_4__58_ ( .D(n6402), .CLK(clk), .Q(ram[1733]) );
  DFFPOSX1 ram_reg_4__59_ ( .D(n6401), .CLK(clk), .Q(ram[1732]) );
  DFFPOSX1 ram_reg_4__60_ ( .D(n6400), .CLK(clk), .Q(ram[1731]) );
  DFFPOSX1 ram_reg_4__61_ ( .D(n6399), .CLK(clk), .Q(ram[1730]) );
  DFFPOSX1 ram_reg_4__62_ ( .D(n6398), .CLK(clk), .Q(ram[1729]) );
  DFFPOSX1 ram_reg_4__63_ ( .D(n6397), .CLK(clk), .Q(ram[1728]) );
  DFFPOSX1 ram_reg_5__0_ ( .D(n6396), .CLK(clk), .Q(ram[1727]) );
  DFFPOSX1 ram_reg_5__1_ ( .D(n6395), .CLK(clk), .Q(ram[1726]) );
  DFFPOSX1 ram_reg_5__2_ ( .D(n6394), .CLK(clk), .Q(ram[1725]) );
  DFFPOSX1 ram_reg_5__3_ ( .D(n6393), .CLK(clk), .Q(ram[1724]) );
  DFFPOSX1 ram_reg_5__4_ ( .D(n6392), .CLK(clk), .Q(ram[1723]) );
  DFFPOSX1 ram_reg_5__5_ ( .D(n6391), .CLK(clk), .Q(ram[1722]) );
  DFFPOSX1 ram_reg_5__6_ ( .D(n6390), .CLK(clk), .Q(ram[1721]) );
  DFFPOSX1 ram_reg_5__7_ ( .D(n6389), .CLK(clk), .Q(ram[1720]) );
  DFFPOSX1 ram_reg_5__8_ ( .D(n6388), .CLK(clk), .Q(ram[1719]) );
  DFFPOSX1 ram_reg_5__9_ ( .D(n6387), .CLK(clk), .Q(ram[1718]) );
  DFFPOSX1 ram_reg_5__10_ ( .D(n6386), .CLK(clk), .Q(ram[1717]) );
  DFFPOSX1 ram_reg_5__11_ ( .D(n6385), .CLK(clk), .Q(ram[1716]) );
  DFFPOSX1 ram_reg_5__12_ ( .D(n6384), .CLK(clk), .Q(ram[1715]) );
  DFFPOSX1 ram_reg_5__13_ ( .D(n6383), .CLK(clk), .Q(ram[1714]) );
  DFFPOSX1 ram_reg_5__14_ ( .D(n6382), .CLK(clk), .Q(ram[1713]) );
  DFFPOSX1 ram_reg_5__15_ ( .D(n6381), .CLK(clk), .Q(ram[1712]) );
  DFFPOSX1 ram_reg_5__16_ ( .D(n6380), .CLK(clk), .Q(ram[1711]) );
  DFFPOSX1 ram_reg_5__17_ ( .D(n6379), .CLK(clk), .Q(ram[1710]) );
  DFFPOSX1 ram_reg_5__18_ ( .D(n6378), .CLK(clk), .Q(ram[1709]) );
  DFFPOSX1 ram_reg_5__19_ ( .D(n6377), .CLK(clk), .Q(ram[1708]) );
  DFFPOSX1 ram_reg_5__20_ ( .D(n6376), .CLK(clk), .Q(ram[1707]) );
  DFFPOSX1 ram_reg_5__21_ ( .D(n6375), .CLK(clk), .Q(ram[1706]) );
  DFFPOSX1 ram_reg_5__22_ ( .D(n6374), .CLK(clk), .Q(ram[1705]) );
  DFFPOSX1 ram_reg_5__23_ ( .D(n6373), .CLK(clk), .Q(ram[1704]) );
  DFFPOSX1 ram_reg_5__24_ ( .D(n6372), .CLK(clk), .Q(ram[1703]) );
  DFFPOSX1 ram_reg_5__25_ ( .D(n6371), .CLK(clk), .Q(ram[1702]) );
  DFFPOSX1 ram_reg_5__26_ ( .D(n6370), .CLK(clk), .Q(ram[1701]) );
  DFFPOSX1 ram_reg_5__27_ ( .D(n6369), .CLK(clk), .Q(ram[1700]) );
  DFFPOSX1 ram_reg_5__28_ ( .D(n6368), .CLK(clk), .Q(ram[1699]) );
  DFFPOSX1 ram_reg_5__29_ ( .D(n6367), .CLK(clk), .Q(ram[1698]) );
  DFFPOSX1 ram_reg_5__30_ ( .D(n6366), .CLK(clk), .Q(ram[1697]) );
  DFFPOSX1 ram_reg_5__31_ ( .D(n6365), .CLK(clk), .Q(ram[1696]) );
  DFFPOSX1 ram_reg_5__32_ ( .D(n6364), .CLK(clk), .Q(ram[1695]) );
  DFFPOSX1 ram_reg_5__33_ ( .D(n6363), .CLK(clk), .Q(ram[1694]) );
  DFFPOSX1 ram_reg_5__34_ ( .D(n6362), .CLK(clk), .Q(ram[1693]) );
  DFFPOSX1 ram_reg_5__35_ ( .D(n6361), .CLK(clk), .Q(ram[1692]) );
  DFFPOSX1 ram_reg_5__36_ ( .D(n6360), .CLK(clk), .Q(ram[1691]) );
  DFFPOSX1 ram_reg_5__37_ ( .D(n6359), .CLK(clk), .Q(ram[1690]) );
  DFFPOSX1 ram_reg_5__38_ ( .D(n6358), .CLK(clk), .Q(ram[1689]) );
  DFFPOSX1 ram_reg_5__39_ ( .D(n6357), .CLK(clk), .Q(ram[1688]) );
  DFFPOSX1 ram_reg_5__40_ ( .D(n6356), .CLK(clk), .Q(ram[1687]) );
  DFFPOSX1 ram_reg_5__41_ ( .D(n6355), .CLK(clk), .Q(ram[1686]) );
  DFFPOSX1 ram_reg_5__42_ ( .D(n6354), .CLK(clk), .Q(ram[1685]) );
  DFFPOSX1 ram_reg_5__43_ ( .D(n6353), .CLK(clk), .Q(ram[1684]) );
  DFFPOSX1 ram_reg_5__44_ ( .D(n6352), .CLK(clk), .Q(ram[1683]) );
  DFFPOSX1 ram_reg_5__45_ ( .D(n6351), .CLK(clk), .Q(ram[1682]) );
  DFFPOSX1 ram_reg_5__46_ ( .D(n6350), .CLK(clk), .Q(ram[1681]) );
  DFFPOSX1 ram_reg_5__47_ ( .D(n6349), .CLK(clk), .Q(ram[1680]) );
  DFFPOSX1 ram_reg_5__48_ ( .D(n6348), .CLK(clk), .Q(ram[1679]) );
  DFFPOSX1 ram_reg_5__49_ ( .D(n6347), .CLK(clk), .Q(ram[1678]) );
  DFFPOSX1 ram_reg_5__50_ ( .D(n6346), .CLK(clk), .Q(ram[1677]) );
  DFFPOSX1 ram_reg_5__51_ ( .D(n6345), .CLK(clk), .Q(ram[1676]) );
  DFFPOSX1 ram_reg_5__52_ ( .D(n6344), .CLK(clk), .Q(ram[1675]) );
  DFFPOSX1 ram_reg_5__53_ ( .D(n6343), .CLK(clk), .Q(ram[1674]) );
  DFFPOSX1 ram_reg_5__54_ ( .D(n6342), .CLK(clk), .Q(ram[1673]) );
  DFFPOSX1 ram_reg_5__55_ ( .D(n6341), .CLK(clk), .Q(ram[1672]) );
  DFFPOSX1 ram_reg_5__56_ ( .D(n6340), .CLK(clk), .Q(ram[1671]) );
  DFFPOSX1 ram_reg_5__57_ ( .D(n6339), .CLK(clk), .Q(ram[1670]) );
  DFFPOSX1 ram_reg_5__58_ ( .D(n6338), .CLK(clk), .Q(ram[1669]) );
  DFFPOSX1 ram_reg_5__59_ ( .D(n6337), .CLK(clk), .Q(ram[1668]) );
  DFFPOSX1 ram_reg_5__60_ ( .D(n6336), .CLK(clk), .Q(ram[1667]) );
  DFFPOSX1 ram_reg_5__61_ ( .D(n6335), .CLK(clk), .Q(ram[1666]) );
  DFFPOSX1 ram_reg_5__62_ ( .D(n6334), .CLK(clk), .Q(ram[1665]) );
  DFFPOSX1 ram_reg_5__63_ ( .D(n6333), .CLK(clk), .Q(ram[1664]) );
  DFFPOSX1 ram_reg_6__0_ ( .D(n6332), .CLK(clk), .Q(ram[1663]) );
  DFFPOSX1 ram_reg_6__1_ ( .D(n6331), .CLK(clk), .Q(ram[1662]) );
  DFFPOSX1 ram_reg_6__2_ ( .D(n6330), .CLK(clk), .Q(ram[1661]) );
  DFFPOSX1 ram_reg_6__3_ ( .D(n6329), .CLK(clk), .Q(ram[1660]) );
  DFFPOSX1 ram_reg_6__4_ ( .D(n6328), .CLK(clk), .Q(ram[1659]) );
  DFFPOSX1 ram_reg_6__5_ ( .D(n6327), .CLK(clk), .Q(ram[1658]) );
  DFFPOSX1 ram_reg_6__6_ ( .D(n6326), .CLK(clk), .Q(ram[1657]) );
  DFFPOSX1 ram_reg_6__7_ ( .D(n6325), .CLK(clk), .Q(ram[1656]) );
  DFFPOSX1 ram_reg_6__8_ ( .D(n6324), .CLK(clk), .Q(ram[1655]) );
  DFFPOSX1 ram_reg_6__9_ ( .D(n6323), .CLK(clk), .Q(ram[1654]) );
  DFFPOSX1 ram_reg_6__10_ ( .D(n6322), .CLK(clk), .Q(ram[1653]) );
  DFFPOSX1 ram_reg_6__11_ ( .D(n6321), .CLK(clk), .Q(ram[1652]) );
  DFFPOSX1 ram_reg_6__12_ ( .D(n6320), .CLK(clk), .Q(ram[1651]) );
  DFFPOSX1 ram_reg_6__13_ ( .D(n6319), .CLK(clk), .Q(ram[1650]) );
  DFFPOSX1 ram_reg_6__14_ ( .D(n6318), .CLK(clk), .Q(ram[1649]) );
  DFFPOSX1 ram_reg_6__15_ ( .D(n6317), .CLK(clk), .Q(ram[1648]) );
  DFFPOSX1 ram_reg_6__16_ ( .D(n6316), .CLK(clk), .Q(ram[1647]) );
  DFFPOSX1 ram_reg_6__17_ ( .D(n6315), .CLK(clk), .Q(ram[1646]) );
  DFFPOSX1 ram_reg_6__18_ ( .D(n6314), .CLK(clk), .Q(ram[1645]) );
  DFFPOSX1 ram_reg_6__19_ ( .D(n6313), .CLK(clk), .Q(ram[1644]) );
  DFFPOSX1 ram_reg_6__20_ ( .D(n6312), .CLK(clk), .Q(ram[1643]) );
  DFFPOSX1 ram_reg_6__21_ ( .D(n6311), .CLK(clk), .Q(ram[1642]) );
  DFFPOSX1 ram_reg_6__22_ ( .D(n6310), .CLK(clk), .Q(ram[1641]) );
  DFFPOSX1 ram_reg_6__23_ ( .D(n6309), .CLK(clk), .Q(ram[1640]) );
  DFFPOSX1 ram_reg_6__24_ ( .D(n6308), .CLK(clk), .Q(ram[1639]) );
  DFFPOSX1 ram_reg_6__25_ ( .D(n6307), .CLK(clk), .Q(ram[1638]) );
  DFFPOSX1 ram_reg_6__26_ ( .D(n6306), .CLK(clk), .Q(ram[1637]) );
  DFFPOSX1 ram_reg_6__27_ ( .D(n6305), .CLK(clk), .Q(ram[1636]) );
  DFFPOSX1 ram_reg_6__28_ ( .D(n6304), .CLK(clk), .Q(ram[1635]) );
  DFFPOSX1 ram_reg_6__29_ ( .D(n6303), .CLK(clk), .Q(ram[1634]) );
  DFFPOSX1 ram_reg_6__30_ ( .D(n6302), .CLK(clk), .Q(ram[1633]) );
  DFFPOSX1 ram_reg_6__31_ ( .D(n6301), .CLK(clk), .Q(ram[1632]) );
  DFFPOSX1 ram_reg_6__32_ ( .D(n6300), .CLK(clk), .Q(ram[1631]) );
  DFFPOSX1 ram_reg_6__33_ ( .D(n6299), .CLK(clk), .Q(ram[1630]) );
  DFFPOSX1 ram_reg_6__34_ ( .D(n6298), .CLK(clk), .Q(ram[1629]) );
  DFFPOSX1 ram_reg_6__35_ ( .D(n6297), .CLK(clk), .Q(ram[1628]) );
  DFFPOSX1 ram_reg_6__36_ ( .D(n6296), .CLK(clk), .Q(ram[1627]) );
  DFFPOSX1 ram_reg_6__37_ ( .D(n6295), .CLK(clk), .Q(ram[1626]) );
  DFFPOSX1 ram_reg_6__38_ ( .D(n6294), .CLK(clk), .Q(ram[1625]) );
  DFFPOSX1 ram_reg_6__39_ ( .D(n6293), .CLK(clk), .Q(ram[1624]) );
  DFFPOSX1 ram_reg_6__40_ ( .D(n6292), .CLK(clk), .Q(ram[1623]) );
  DFFPOSX1 ram_reg_6__41_ ( .D(n6291), .CLK(clk), .Q(ram[1622]) );
  DFFPOSX1 ram_reg_6__42_ ( .D(n6290), .CLK(clk), .Q(ram[1621]) );
  DFFPOSX1 ram_reg_6__43_ ( .D(n6289), .CLK(clk), .Q(ram[1620]) );
  DFFPOSX1 ram_reg_6__44_ ( .D(n6288), .CLK(clk), .Q(ram[1619]) );
  DFFPOSX1 ram_reg_6__45_ ( .D(n6287), .CLK(clk), .Q(ram[1618]) );
  DFFPOSX1 ram_reg_6__46_ ( .D(n6286), .CLK(clk), .Q(ram[1617]) );
  DFFPOSX1 ram_reg_6__47_ ( .D(n6285), .CLK(clk), .Q(ram[1616]) );
  DFFPOSX1 ram_reg_6__48_ ( .D(n6284), .CLK(clk), .Q(ram[1615]) );
  DFFPOSX1 ram_reg_6__49_ ( .D(n6283), .CLK(clk), .Q(ram[1614]) );
  DFFPOSX1 ram_reg_6__50_ ( .D(n6282), .CLK(clk), .Q(ram[1613]) );
  DFFPOSX1 ram_reg_6__51_ ( .D(n6281), .CLK(clk), .Q(ram[1612]) );
  DFFPOSX1 ram_reg_6__52_ ( .D(n6280), .CLK(clk), .Q(ram[1611]) );
  DFFPOSX1 ram_reg_6__53_ ( .D(n6279), .CLK(clk), .Q(ram[1610]) );
  DFFPOSX1 ram_reg_6__54_ ( .D(n6278), .CLK(clk), .Q(ram[1609]) );
  DFFPOSX1 ram_reg_6__55_ ( .D(n6277), .CLK(clk), .Q(ram[1608]) );
  DFFPOSX1 ram_reg_6__56_ ( .D(n6276), .CLK(clk), .Q(ram[1607]) );
  DFFPOSX1 ram_reg_6__57_ ( .D(n6275), .CLK(clk), .Q(ram[1606]) );
  DFFPOSX1 ram_reg_6__58_ ( .D(n6274), .CLK(clk), .Q(ram[1605]) );
  DFFPOSX1 ram_reg_6__59_ ( .D(n6273), .CLK(clk), .Q(ram[1604]) );
  DFFPOSX1 ram_reg_6__60_ ( .D(n6272), .CLK(clk), .Q(ram[1603]) );
  DFFPOSX1 ram_reg_6__61_ ( .D(n6271), .CLK(clk), .Q(ram[1602]) );
  DFFPOSX1 ram_reg_6__62_ ( .D(n6270), .CLK(clk), .Q(ram[1601]) );
  DFFPOSX1 ram_reg_6__63_ ( .D(n6269), .CLK(clk), .Q(ram[1600]) );
  DFFPOSX1 ram_reg_7__0_ ( .D(n6268), .CLK(clk), .Q(ram[1599]) );
  DFFPOSX1 ram_reg_7__1_ ( .D(n6267), .CLK(clk), .Q(ram[1598]) );
  DFFPOSX1 ram_reg_7__2_ ( .D(n6266), .CLK(clk), .Q(ram[1597]) );
  DFFPOSX1 ram_reg_7__3_ ( .D(n6265), .CLK(clk), .Q(ram[1596]) );
  DFFPOSX1 ram_reg_7__4_ ( .D(n6264), .CLK(clk), .Q(ram[1595]) );
  DFFPOSX1 ram_reg_7__5_ ( .D(n6263), .CLK(clk), .Q(ram[1594]) );
  DFFPOSX1 ram_reg_7__6_ ( .D(n6262), .CLK(clk), .Q(ram[1593]) );
  DFFPOSX1 ram_reg_7__7_ ( .D(n6261), .CLK(clk), .Q(ram[1592]) );
  DFFPOSX1 ram_reg_7__8_ ( .D(n6260), .CLK(clk), .Q(ram[1591]) );
  DFFPOSX1 ram_reg_7__9_ ( .D(n6259), .CLK(clk), .Q(ram[1590]) );
  DFFPOSX1 ram_reg_7__10_ ( .D(n6258), .CLK(clk), .Q(ram[1589]) );
  DFFPOSX1 ram_reg_7__11_ ( .D(n6257), .CLK(clk), .Q(ram[1588]) );
  DFFPOSX1 ram_reg_7__12_ ( .D(n6256), .CLK(clk), .Q(ram[1587]) );
  DFFPOSX1 ram_reg_7__13_ ( .D(n6255), .CLK(clk), .Q(ram[1586]) );
  DFFPOSX1 ram_reg_7__14_ ( .D(n6254), .CLK(clk), .Q(ram[1585]) );
  DFFPOSX1 ram_reg_7__15_ ( .D(n6253), .CLK(clk), .Q(ram[1584]) );
  DFFPOSX1 ram_reg_7__16_ ( .D(n6252), .CLK(clk), .Q(ram[1583]) );
  DFFPOSX1 ram_reg_7__17_ ( .D(n6251), .CLK(clk), .Q(ram[1582]) );
  DFFPOSX1 ram_reg_7__18_ ( .D(n6250), .CLK(clk), .Q(ram[1581]) );
  DFFPOSX1 ram_reg_7__19_ ( .D(n6249), .CLK(clk), .Q(ram[1580]) );
  DFFPOSX1 ram_reg_7__20_ ( .D(n6248), .CLK(clk), .Q(ram[1579]) );
  DFFPOSX1 ram_reg_7__21_ ( .D(n6247), .CLK(clk), .Q(ram[1578]) );
  DFFPOSX1 ram_reg_7__22_ ( .D(n6246), .CLK(clk), .Q(ram[1577]) );
  DFFPOSX1 ram_reg_7__23_ ( .D(n6245), .CLK(clk), .Q(ram[1576]) );
  DFFPOSX1 ram_reg_7__24_ ( .D(n6244), .CLK(clk), .Q(ram[1575]) );
  DFFPOSX1 ram_reg_7__25_ ( .D(n6243), .CLK(clk), .Q(ram[1574]) );
  DFFPOSX1 ram_reg_7__26_ ( .D(n6242), .CLK(clk), .Q(ram[1573]) );
  DFFPOSX1 ram_reg_7__27_ ( .D(n6241), .CLK(clk), .Q(ram[1572]) );
  DFFPOSX1 ram_reg_7__28_ ( .D(n6240), .CLK(clk), .Q(ram[1571]) );
  DFFPOSX1 ram_reg_7__29_ ( .D(n6239), .CLK(clk), .Q(ram[1570]) );
  DFFPOSX1 ram_reg_7__30_ ( .D(n6238), .CLK(clk), .Q(ram[1569]) );
  DFFPOSX1 ram_reg_7__31_ ( .D(n6237), .CLK(clk), .Q(ram[1568]) );
  DFFPOSX1 ram_reg_7__32_ ( .D(n6236), .CLK(clk), .Q(ram[1567]) );
  DFFPOSX1 ram_reg_7__33_ ( .D(n6235), .CLK(clk), .Q(ram[1566]) );
  DFFPOSX1 ram_reg_7__34_ ( .D(n6234), .CLK(clk), .Q(ram[1565]) );
  DFFPOSX1 ram_reg_7__35_ ( .D(n6233), .CLK(clk), .Q(ram[1564]) );
  DFFPOSX1 ram_reg_7__36_ ( .D(n6232), .CLK(clk), .Q(ram[1563]) );
  DFFPOSX1 ram_reg_7__37_ ( .D(n6231), .CLK(clk), .Q(ram[1562]) );
  DFFPOSX1 ram_reg_7__38_ ( .D(n6230), .CLK(clk), .Q(ram[1561]) );
  DFFPOSX1 ram_reg_7__39_ ( .D(n6229), .CLK(clk), .Q(ram[1560]) );
  DFFPOSX1 ram_reg_7__40_ ( .D(n6228), .CLK(clk), .Q(ram[1559]) );
  DFFPOSX1 ram_reg_7__41_ ( .D(n6227), .CLK(clk), .Q(ram[1558]) );
  DFFPOSX1 ram_reg_7__42_ ( .D(n6226), .CLK(clk), .Q(ram[1557]) );
  DFFPOSX1 ram_reg_7__43_ ( .D(n6225), .CLK(clk), .Q(ram[1556]) );
  DFFPOSX1 ram_reg_7__44_ ( .D(n6224), .CLK(clk), .Q(ram[1555]) );
  DFFPOSX1 ram_reg_7__45_ ( .D(n6223), .CLK(clk), .Q(ram[1554]) );
  DFFPOSX1 ram_reg_7__46_ ( .D(n6222), .CLK(clk), .Q(ram[1553]) );
  DFFPOSX1 ram_reg_7__47_ ( .D(n6221), .CLK(clk), .Q(ram[1552]) );
  DFFPOSX1 ram_reg_7__48_ ( .D(n6220), .CLK(clk), .Q(ram[1551]) );
  DFFPOSX1 ram_reg_7__49_ ( .D(n6219), .CLK(clk), .Q(ram[1550]) );
  DFFPOSX1 ram_reg_7__50_ ( .D(n6218), .CLK(clk), .Q(ram[1549]) );
  DFFPOSX1 ram_reg_7__51_ ( .D(n6217), .CLK(clk), .Q(ram[1548]) );
  DFFPOSX1 ram_reg_7__52_ ( .D(n6216), .CLK(clk), .Q(ram[1547]) );
  DFFPOSX1 ram_reg_7__53_ ( .D(n6215), .CLK(clk), .Q(ram[1546]) );
  DFFPOSX1 ram_reg_7__54_ ( .D(n6214), .CLK(clk), .Q(ram[1545]) );
  DFFPOSX1 ram_reg_7__55_ ( .D(n6213), .CLK(clk), .Q(ram[1544]) );
  DFFPOSX1 ram_reg_7__56_ ( .D(n6212), .CLK(clk), .Q(ram[1543]) );
  DFFPOSX1 ram_reg_7__57_ ( .D(n6211), .CLK(clk), .Q(ram[1542]) );
  DFFPOSX1 ram_reg_7__58_ ( .D(n6210), .CLK(clk), .Q(ram[1541]) );
  DFFPOSX1 ram_reg_7__59_ ( .D(n6209), .CLK(clk), .Q(ram[1540]) );
  DFFPOSX1 ram_reg_7__60_ ( .D(n6208), .CLK(clk), .Q(ram[1539]) );
  DFFPOSX1 ram_reg_7__61_ ( .D(n6207), .CLK(clk), .Q(ram[1538]) );
  DFFPOSX1 ram_reg_7__62_ ( .D(n6206), .CLK(clk), .Q(ram[1537]) );
  DFFPOSX1 ram_reg_7__63_ ( .D(n6205), .CLK(clk), .Q(ram[1536]) );
  DFFPOSX1 ram_reg_8__0_ ( .D(n6204), .CLK(clk), .Q(ram[1535]) );
  DFFPOSX1 ram_reg_8__1_ ( .D(n6203), .CLK(clk), .Q(ram[1534]) );
  DFFPOSX1 ram_reg_8__2_ ( .D(n6202), .CLK(clk), .Q(ram[1533]) );
  DFFPOSX1 ram_reg_8__3_ ( .D(n6201), .CLK(clk), .Q(ram[1532]) );
  DFFPOSX1 ram_reg_8__4_ ( .D(n6200), .CLK(clk), .Q(ram[1531]) );
  DFFPOSX1 ram_reg_8__5_ ( .D(n6199), .CLK(clk), .Q(ram[1530]) );
  DFFPOSX1 ram_reg_8__6_ ( .D(n6198), .CLK(clk), .Q(ram[1529]) );
  DFFPOSX1 ram_reg_8__7_ ( .D(n6197), .CLK(clk), .Q(ram[1528]) );
  DFFPOSX1 ram_reg_8__8_ ( .D(n6196), .CLK(clk), .Q(ram[1527]) );
  DFFPOSX1 ram_reg_8__9_ ( .D(n6195), .CLK(clk), .Q(ram[1526]) );
  DFFPOSX1 ram_reg_8__10_ ( .D(n6194), .CLK(clk), .Q(ram[1525]) );
  DFFPOSX1 ram_reg_8__11_ ( .D(n6193), .CLK(clk), .Q(ram[1524]) );
  DFFPOSX1 ram_reg_8__12_ ( .D(n6192), .CLK(clk), .Q(ram[1523]) );
  DFFPOSX1 ram_reg_8__13_ ( .D(n6191), .CLK(clk), .Q(ram[1522]) );
  DFFPOSX1 ram_reg_8__14_ ( .D(n6190), .CLK(clk), .Q(ram[1521]) );
  DFFPOSX1 ram_reg_8__15_ ( .D(n6189), .CLK(clk), .Q(ram[1520]) );
  DFFPOSX1 ram_reg_8__16_ ( .D(n6188), .CLK(clk), .Q(ram[1519]) );
  DFFPOSX1 ram_reg_8__17_ ( .D(n6187), .CLK(clk), .Q(ram[1518]) );
  DFFPOSX1 ram_reg_8__18_ ( .D(n6186), .CLK(clk), .Q(ram[1517]) );
  DFFPOSX1 ram_reg_8__19_ ( .D(n6185), .CLK(clk), .Q(ram[1516]) );
  DFFPOSX1 ram_reg_8__20_ ( .D(n6184), .CLK(clk), .Q(ram[1515]) );
  DFFPOSX1 ram_reg_8__21_ ( .D(n6183), .CLK(clk), .Q(ram[1514]) );
  DFFPOSX1 ram_reg_8__22_ ( .D(n6182), .CLK(clk), .Q(ram[1513]) );
  DFFPOSX1 ram_reg_8__23_ ( .D(n6181), .CLK(clk), .Q(ram[1512]) );
  DFFPOSX1 ram_reg_8__24_ ( .D(n6180), .CLK(clk), .Q(ram[1511]) );
  DFFPOSX1 ram_reg_8__25_ ( .D(n6179), .CLK(clk), .Q(ram[1510]) );
  DFFPOSX1 ram_reg_8__26_ ( .D(n6178), .CLK(clk), .Q(ram[1509]) );
  DFFPOSX1 ram_reg_8__27_ ( .D(n6177), .CLK(clk), .Q(ram[1508]) );
  DFFPOSX1 ram_reg_8__28_ ( .D(n6176), .CLK(clk), .Q(ram[1507]) );
  DFFPOSX1 ram_reg_8__29_ ( .D(n6175), .CLK(clk), .Q(ram[1506]) );
  DFFPOSX1 ram_reg_8__30_ ( .D(n6174), .CLK(clk), .Q(ram[1505]) );
  DFFPOSX1 ram_reg_8__31_ ( .D(n6173), .CLK(clk), .Q(ram[1504]) );
  DFFPOSX1 ram_reg_8__32_ ( .D(n6172), .CLK(clk), .Q(ram[1503]) );
  DFFPOSX1 ram_reg_8__33_ ( .D(n6171), .CLK(clk), .Q(ram[1502]) );
  DFFPOSX1 ram_reg_8__34_ ( .D(n6170), .CLK(clk), .Q(ram[1501]) );
  DFFPOSX1 ram_reg_8__35_ ( .D(n6169), .CLK(clk), .Q(ram[1500]) );
  DFFPOSX1 ram_reg_8__36_ ( .D(n6168), .CLK(clk), .Q(ram[1499]) );
  DFFPOSX1 ram_reg_8__37_ ( .D(n6167), .CLK(clk), .Q(ram[1498]) );
  DFFPOSX1 ram_reg_8__38_ ( .D(n6166), .CLK(clk), .Q(ram[1497]) );
  DFFPOSX1 ram_reg_8__39_ ( .D(n6165), .CLK(clk), .Q(ram[1496]) );
  DFFPOSX1 ram_reg_8__40_ ( .D(n6164), .CLK(clk), .Q(ram[1495]) );
  DFFPOSX1 ram_reg_8__41_ ( .D(n6163), .CLK(clk), .Q(ram[1494]) );
  DFFPOSX1 ram_reg_8__42_ ( .D(n6162), .CLK(clk), .Q(ram[1493]) );
  DFFPOSX1 ram_reg_8__43_ ( .D(n6161), .CLK(clk), .Q(ram[1492]) );
  DFFPOSX1 ram_reg_8__44_ ( .D(n6160), .CLK(clk), .Q(ram[1491]) );
  DFFPOSX1 ram_reg_8__45_ ( .D(n6159), .CLK(clk), .Q(ram[1490]) );
  DFFPOSX1 ram_reg_8__46_ ( .D(n6158), .CLK(clk), .Q(ram[1489]) );
  DFFPOSX1 ram_reg_8__47_ ( .D(n6157), .CLK(clk), .Q(ram[1488]) );
  DFFPOSX1 ram_reg_8__48_ ( .D(n6156), .CLK(clk), .Q(ram[1487]) );
  DFFPOSX1 ram_reg_8__49_ ( .D(n6155), .CLK(clk), .Q(ram[1486]) );
  DFFPOSX1 ram_reg_8__50_ ( .D(n6154), .CLK(clk), .Q(ram[1485]) );
  DFFPOSX1 ram_reg_8__51_ ( .D(n6153), .CLK(clk), .Q(ram[1484]) );
  DFFPOSX1 ram_reg_8__52_ ( .D(n6152), .CLK(clk), .Q(ram[1483]) );
  DFFPOSX1 ram_reg_8__53_ ( .D(n6151), .CLK(clk), .Q(ram[1482]) );
  DFFPOSX1 ram_reg_8__54_ ( .D(n6150), .CLK(clk), .Q(ram[1481]) );
  DFFPOSX1 ram_reg_8__55_ ( .D(n6149), .CLK(clk), .Q(ram[1480]) );
  DFFPOSX1 ram_reg_8__56_ ( .D(n6148), .CLK(clk), .Q(ram[1479]) );
  DFFPOSX1 ram_reg_8__57_ ( .D(n6147), .CLK(clk), .Q(ram[1478]) );
  DFFPOSX1 ram_reg_8__58_ ( .D(n6146), .CLK(clk), .Q(ram[1477]) );
  DFFPOSX1 ram_reg_8__59_ ( .D(n6145), .CLK(clk), .Q(ram[1476]) );
  DFFPOSX1 ram_reg_8__60_ ( .D(n6144), .CLK(clk), .Q(ram[1475]) );
  DFFPOSX1 ram_reg_8__61_ ( .D(n6143), .CLK(clk), .Q(ram[1474]) );
  DFFPOSX1 ram_reg_8__62_ ( .D(n6142), .CLK(clk), .Q(ram[1473]) );
  DFFPOSX1 ram_reg_8__63_ ( .D(n6141), .CLK(clk), .Q(ram[1472]) );
  DFFPOSX1 ram_reg_9__0_ ( .D(n6140), .CLK(clk), .Q(ram[1471]) );
  DFFPOSX1 ram_reg_9__1_ ( .D(n6139), .CLK(clk), .Q(ram[1470]) );
  DFFPOSX1 ram_reg_9__2_ ( .D(n6138), .CLK(clk), .Q(ram[1469]) );
  DFFPOSX1 ram_reg_9__3_ ( .D(n6137), .CLK(clk), .Q(ram[1468]) );
  DFFPOSX1 ram_reg_9__4_ ( .D(n6136), .CLK(clk), .Q(ram[1467]) );
  DFFPOSX1 ram_reg_9__5_ ( .D(n6135), .CLK(clk), .Q(ram[1466]) );
  DFFPOSX1 ram_reg_9__6_ ( .D(n6134), .CLK(clk), .Q(ram[1465]) );
  DFFPOSX1 ram_reg_9__7_ ( .D(n6133), .CLK(clk), .Q(ram[1464]) );
  DFFPOSX1 ram_reg_9__8_ ( .D(n6132), .CLK(clk), .Q(ram[1463]) );
  DFFPOSX1 ram_reg_9__9_ ( .D(n6131), .CLK(clk), .Q(ram[1462]) );
  DFFPOSX1 ram_reg_9__10_ ( .D(n6130), .CLK(clk), .Q(ram[1461]) );
  DFFPOSX1 ram_reg_9__11_ ( .D(n6129), .CLK(clk), .Q(ram[1460]) );
  DFFPOSX1 ram_reg_9__12_ ( .D(n6128), .CLK(clk), .Q(ram[1459]) );
  DFFPOSX1 ram_reg_9__13_ ( .D(n6127), .CLK(clk), .Q(ram[1458]) );
  DFFPOSX1 ram_reg_9__14_ ( .D(n6126), .CLK(clk), .Q(ram[1457]) );
  DFFPOSX1 ram_reg_9__15_ ( .D(n6125), .CLK(clk), .Q(ram[1456]) );
  DFFPOSX1 ram_reg_9__16_ ( .D(n6124), .CLK(clk), .Q(ram[1455]) );
  DFFPOSX1 ram_reg_9__17_ ( .D(n6123), .CLK(clk), .Q(ram[1454]) );
  DFFPOSX1 ram_reg_9__18_ ( .D(n6122), .CLK(clk), .Q(ram[1453]) );
  DFFPOSX1 ram_reg_9__19_ ( .D(n6121), .CLK(clk), .Q(ram[1452]) );
  DFFPOSX1 ram_reg_9__20_ ( .D(n6120), .CLK(clk), .Q(ram[1451]) );
  DFFPOSX1 ram_reg_9__21_ ( .D(n6119), .CLK(clk), .Q(ram[1450]) );
  DFFPOSX1 ram_reg_9__22_ ( .D(n6118), .CLK(clk), .Q(ram[1449]) );
  DFFPOSX1 ram_reg_9__23_ ( .D(n6117), .CLK(clk), .Q(ram[1448]) );
  DFFPOSX1 ram_reg_9__24_ ( .D(n6116), .CLK(clk), .Q(ram[1447]) );
  DFFPOSX1 ram_reg_9__25_ ( .D(n6115), .CLK(clk), .Q(ram[1446]) );
  DFFPOSX1 ram_reg_9__26_ ( .D(n6114), .CLK(clk), .Q(ram[1445]) );
  DFFPOSX1 ram_reg_9__27_ ( .D(n6113), .CLK(clk), .Q(ram[1444]) );
  DFFPOSX1 ram_reg_9__28_ ( .D(n6112), .CLK(clk), .Q(ram[1443]) );
  DFFPOSX1 ram_reg_9__29_ ( .D(n6111), .CLK(clk), .Q(ram[1442]) );
  DFFPOSX1 ram_reg_9__30_ ( .D(n6110), .CLK(clk), .Q(ram[1441]) );
  DFFPOSX1 ram_reg_9__31_ ( .D(n6109), .CLK(clk), .Q(ram[1440]) );
  DFFPOSX1 ram_reg_9__32_ ( .D(n6108), .CLK(clk), .Q(ram[1439]) );
  DFFPOSX1 ram_reg_9__33_ ( .D(n6107), .CLK(clk), .Q(ram[1438]) );
  DFFPOSX1 ram_reg_9__34_ ( .D(n6106), .CLK(clk), .Q(ram[1437]) );
  DFFPOSX1 ram_reg_9__35_ ( .D(n6105), .CLK(clk), .Q(ram[1436]) );
  DFFPOSX1 ram_reg_9__36_ ( .D(n6104), .CLK(clk), .Q(ram[1435]) );
  DFFPOSX1 ram_reg_9__37_ ( .D(n6103), .CLK(clk), .Q(ram[1434]) );
  DFFPOSX1 ram_reg_9__38_ ( .D(n6102), .CLK(clk), .Q(ram[1433]) );
  DFFPOSX1 ram_reg_9__39_ ( .D(n6101), .CLK(clk), .Q(ram[1432]) );
  DFFPOSX1 ram_reg_9__40_ ( .D(n6100), .CLK(clk), .Q(ram[1431]) );
  DFFPOSX1 ram_reg_9__41_ ( .D(n6099), .CLK(clk), .Q(ram[1430]) );
  DFFPOSX1 ram_reg_9__42_ ( .D(n6098), .CLK(clk), .Q(ram[1429]) );
  DFFPOSX1 ram_reg_9__43_ ( .D(n6097), .CLK(clk), .Q(ram[1428]) );
  DFFPOSX1 ram_reg_9__44_ ( .D(n6096), .CLK(clk), .Q(ram[1427]) );
  DFFPOSX1 ram_reg_9__45_ ( .D(n6095), .CLK(clk), .Q(ram[1426]) );
  DFFPOSX1 ram_reg_9__46_ ( .D(n6094), .CLK(clk), .Q(ram[1425]) );
  DFFPOSX1 ram_reg_9__47_ ( .D(n6093), .CLK(clk), .Q(ram[1424]) );
  DFFPOSX1 ram_reg_9__48_ ( .D(n6092), .CLK(clk), .Q(ram[1423]) );
  DFFPOSX1 ram_reg_9__49_ ( .D(n6091), .CLK(clk), .Q(ram[1422]) );
  DFFPOSX1 ram_reg_9__50_ ( .D(n6090), .CLK(clk), .Q(ram[1421]) );
  DFFPOSX1 ram_reg_9__51_ ( .D(n6089), .CLK(clk), .Q(ram[1420]) );
  DFFPOSX1 ram_reg_9__52_ ( .D(n6088), .CLK(clk), .Q(ram[1419]) );
  DFFPOSX1 ram_reg_9__53_ ( .D(n6087), .CLK(clk), .Q(ram[1418]) );
  DFFPOSX1 ram_reg_9__54_ ( .D(n6086), .CLK(clk), .Q(ram[1417]) );
  DFFPOSX1 ram_reg_9__55_ ( .D(n6085), .CLK(clk), .Q(ram[1416]) );
  DFFPOSX1 ram_reg_9__56_ ( .D(n6084), .CLK(clk), .Q(ram[1415]) );
  DFFPOSX1 ram_reg_9__57_ ( .D(n6083), .CLK(clk), .Q(ram[1414]) );
  DFFPOSX1 ram_reg_9__58_ ( .D(n6082), .CLK(clk), .Q(ram[1413]) );
  DFFPOSX1 ram_reg_9__59_ ( .D(n6081), .CLK(clk), .Q(ram[1412]) );
  DFFPOSX1 ram_reg_9__60_ ( .D(n6080), .CLK(clk), .Q(ram[1411]) );
  DFFPOSX1 ram_reg_9__61_ ( .D(n6079), .CLK(clk), .Q(ram[1410]) );
  DFFPOSX1 ram_reg_9__62_ ( .D(n6078), .CLK(clk), .Q(ram[1409]) );
  DFFPOSX1 ram_reg_9__63_ ( .D(n6077), .CLK(clk), .Q(ram[1408]) );
  DFFPOSX1 ram_reg_10__0_ ( .D(n6076), .CLK(clk), .Q(ram[1407]) );
  DFFPOSX1 ram_reg_10__1_ ( .D(n6075), .CLK(clk), .Q(ram[1406]) );
  DFFPOSX1 ram_reg_10__2_ ( .D(n6074), .CLK(clk), .Q(ram[1405]) );
  DFFPOSX1 ram_reg_10__3_ ( .D(n6073), .CLK(clk), .Q(ram[1404]) );
  DFFPOSX1 ram_reg_10__4_ ( .D(n6072), .CLK(clk), .Q(ram[1403]) );
  DFFPOSX1 ram_reg_10__5_ ( .D(n6071), .CLK(clk), .Q(ram[1402]) );
  DFFPOSX1 ram_reg_10__6_ ( .D(n6070), .CLK(clk), .Q(ram[1401]) );
  DFFPOSX1 ram_reg_10__7_ ( .D(n6069), .CLK(clk), .Q(ram[1400]) );
  DFFPOSX1 ram_reg_10__8_ ( .D(n6068), .CLK(clk), .Q(ram[1399]) );
  DFFPOSX1 ram_reg_10__9_ ( .D(n6067), .CLK(clk), .Q(ram[1398]) );
  DFFPOSX1 ram_reg_10__10_ ( .D(n6066), .CLK(clk), .Q(ram[1397]) );
  DFFPOSX1 ram_reg_10__11_ ( .D(n6065), .CLK(clk), .Q(ram[1396]) );
  DFFPOSX1 ram_reg_10__12_ ( .D(n6064), .CLK(clk), .Q(ram[1395]) );
  DFFPOSX1 ram_reg_10__13_ ( .D(n6063), .CLK(clk), .Q(ram[1394]) );
  DFFPOSX1 ram_reg_10__14_ ( .D(n6062), .CLK(clk), .Q(ram[1393]) );
  DFFPOSX1 ram_reg_10__15_ ( .D(n6061), .CLK(clk), .Q(ram[1392]) );
  DFFPOSX1 ram_reg_10__16_ ( .D(n6060), .CLK(clk), .Q(ram[1391]) );
  DFFPOSX1 ram_reg_10__17_ ( .D(n6059), .CLK(clk), .Q(ram[1390]) );
  DFFPOSX1 ram_reg_10__18_ ( .D(n6058), .CLK(clk), .Q(ram[1389]) );
  DFFPOSX1 ram_reg_10__19_ ( .D(n6057), .CLK(clk), .Q(ram[1388]) );
  DFFPOSX1 ram_reg_10__20_ ( .D(n6056), .CLK(clk), .Q(ram[1387]) );
  DFFPOSX1 ram_reg_10__21_ ( .D(n6055), .CLK(clk), .Q(ram[1386]) );
  DFFPOSX1 ram_reg_10__22_ ( .D(n6054), .CLK(clk), .Q(ram[1385]) );
  DFFPOSX1 ram_reg_10__23_ ( .D(n6053), .CLK(clk), .Q(ram[1384]) );
  DFFPOSX1 ram_reg_10__24_ ( .D(n6052), .CLK(clk), .Q(ram[1383]) );
  DFFPOSX1 ram_reg_10__25_ ( .D(n6051), .CLK(clk), .Q(ram[1382]) );
  DFFPOSX1 ram_reg_10__26_ ( .D(n6050), .CLK(clk), .Q(ram[1381]) );
  DFFPOSX1 ram_reg_10__27_ ( .D(n6049), .CLK(clk), .Q(ram[1380]) );
  DFFPOSX1 ram_reg_10__28_ ( .D(n6048), .CLK(clk), .Q(ram[1379]) );
  DFFPOSX1 ram_reg_10__29_ ( .D(n6047), .CLK(clk), .Q(ram[1378]) );
  DFFPOSX1 ram_reg_10__30_ ( .D(n6046), .CLK(clk), .Q(ram[1377]) );
  DFFPOSX1 ram_reg_10__31_ ( .D(n6045), .CLK(clk), .Q(ram[1376]) );
  DFFPOSX1 ram_reg_10__32_ ( .D(n6044), .CLK(clk), .Q(ram[1375]) );
  DFFPOSX1 ram_reg_10__33_ ( .D(n6043), .CLK(clk), .Q(ram[1374]) );
  DFFPOSX1 ram_reg_10__34_ ( .D(n6042), .CLK(clk), .Q(ram[1373]) );
  DFFPOSX1 ram_reg_10__35_ ( .D(n6041), .CLK(clk), .Q(ram[1372]) );
  DFFPOSX1 ram_reg_10__36_ ( .D(n6040), .CLK(clk), .Q(ram[1371]) );
  DFFPOSX1 ram_reg_10__37_ ( .D(n6039), .CLK(clk), .Q(ram[1370]) );
  DFFPOSX1 ram_reg_10__38_ ( .D(n6038), .CLK(clk), .Q(ram[1369]) );
  DFFPOSX1 ram_reg_10__39_ ( .D(n6037), .CLK(clk), .Q(ram[1368]) );
  DFFPOSX1 ram_reg_10__40_ ( .D(n6036), .CLK(clk), .Q(ram[1367]) );
  DFFPOSX1 ram_reg_10__41_ ( .D(n6035), .CLK(clk), .Q(ram[1366]) );
  DFFPOSX1 ram_reg_10__42_ ( .D(n6034), .CLK(clk), .Q(ram[1365]) );
  DFFPOSX1 ram_reg_10__43_ ( .D(n6033), .CLK(clk), .Q(ram[1364]) );
  DFFPOSX1 ram_reg_10__44_ ( .D(n6032), .CLK(clk), .Q(ram[1363]) );
  DFFPOSX1 ram_reg_10__45_ ( .D(n6031), .CLK(clk), .Q(ram[1362]) );
  DFFPOSX1 ram_reg_10__46_ ( .D(n6030), .CLK(clk), .Q(ram[1361]) );
  DFFPOSX1 ram_reg_10__47_ ( .D(n6029), .CLK(clk), .Q(ram[1360]) );
  DFFPOSX1 ram_reg_10__48_ ( .D(n6028), .CLK(clk), .Q(ram[1359]) );
  DFFPOSX1 ram_reg_10__49_ ( .D(n6027), .CLK(clk), .Q(ram[1358]) );
  DFFPOSX1 ram_reg_10__50_ ( .D(n6026), .CLK(clk), .Q(ram[1357]) );
  DFFPOSX1 ram_reg_10__51_ ( .D(n6025), .CLK(clk), .Q(ram[1356]) );
  DFFPOSX1 ram_reg_10__52_ ( .D(n6024), .CLK(clk), .Q(ram[1355]) );
  DFFPOSX1 ram_reg_10__53_ ( .D(n6023), .CLK(clk), .Q(ram[1354]) );
  DFFPOSX1 ram_reg_10__54_ ( .D(n6022), .CLK(clk), .Q(ram[1353]) );
  DFFPOSX1 ram_reg_10__55_ ( .D(n6021), .CLK(clk), .Q(ram[1352]) );
  DFFPOSX1 ram_reg_10__56_ ( .D(n6020), .CLK(clk), .Q(ram[1351]) );
  DFFPOSX1 ram_reg_10__57_ ( .D(n6019), .CLK(clk), .Q(ram[1350]) );
  DFFPOSX1 ram_reg_10__58_ ( .D(n6018), .CLK(clk), .Q(ram[1349]) );
  DFFPOSX1 ram_reg_10__59_ ( .D(n6017), .CLK(clk), .Q(ram[1348]) );
  DFFPOSX1 ram_reg_10__60_ ( .D(n6016), .CLK(clk), .Q(ram[1347]) );
  DFFPOSX1 ram_reg_10__61_ ( .D(n6015), .CLK(clk), .Q(ram[1346]) );
  DFFPOSX1 ram_reg_10__62_ ( .D(n6014), .CLK(clk), .Q(ram[1345]) );
  DFFPOSX1 ram_reg_10__63_ ( .D(n6013), .CLK(clk), .Q(ram[1344]) );
  DFFPOSX1 ram_reg_11__0_ ( .D(n6012), .CLK(clk), .Q(ram[1343]) );
  DFFPOSX1 ram_reg_11__1_ ( .D(n6011), .CLK(clk), .Q(ram[1342]) );
  DFFPOSX1 ram_reg_11__2_ ( .D(n6010), .CLK(clk), .Q(ram[1341]) );
  DFFPOSX1 ram_reg_11__3_ ( .D(n6009), .CLK(clk), .Q(ram[1340]) );
  DFFPOSX1 ram_reg_11__4_ ( .D(n6008), .CLK(clk), .Q(ram[1339]) );
  DFFPOSX1 ram_reg_11__5_ ( .D(n6007), .CLK(clk), .Q(ram[1338]) );
  DFFPOSX1 ram_reg_11__6_ ( .D(n6006), .CLK(clk), .Q(ram[1337]) );
  DFFPOSX1 ram_reg_11__7_ ( .D(n6005), .CLK(clk), .Q(ram[1336]) );
  DFFPOSX1 ram_reg_11__8_ ( .D(n6004), .CLK(clk), .Q(ram[1335]) );
  DFFPOSX1 ram_reg_11__9_ ( .D(n6003), .CLK(clk), .Q(ram[1334]) );
  DFFPOSX1 ram_reg_11__10_ ( .D(n6002), .CLK(clk), .Q(ram[1333]) );
  DFFPOSX1 ram_reg_11__11_ ( .D(n6001), .CLK(clk), .Q(ram[1332]) );
  DFFPOSX1 ram_reg_11__12_ ( .D(n6000), .CLK(clk), .Q(ram[1331]) );
  DFFPOSX1 ram_reg_11__13_ ( .D(n5999), .CLK(clk), .Q(ram[1330]) );
  DFFPOSX1 ram_reg_11__14_ ( .D(n5998), .CLK(clk), .Q(ram[1329]) );
  DFFPOSX1 ram_reg_11__15_ ( .D(n5997), .CLK(clk), .Q(ram[1328]) );
  DFFPOSX1 ram_reg_11__16_ ( .D(n5996), .CLK(clk), .Q(ram[1327]) );
  DFFPOSX1 ram_reg_11__17_ ( .D(n5995), .CLK(clk), .Q(ram[1326]) );
  DFFPOSX1 ram_reg_11__18_ ( .D(n5994), .CLK(clk), .Q(ram[1325]) );
  DFFPOSX1 ram_reg_11__19_ ( .D(n5993), .CLK(clk), .Q(ram[1324]) );
  DFFPOSX1 ram_reg_11__20_ ( .D(n5992), .CLK(clk), .Q(ram[1323]) );
  DFFPOSX1 ram_reg_11__21_ ( .D(n5991), .CLK(clk), .Q(ram[1322]) );
  DFFPOSX1 ram_reg_11__22_ ( .D(n5990), .CLK(clk), .Q(ram[1321]) );
  DFFPOSX1 ram_reg_11__23_ ( .D(n5989), .CLK(clk), .Q(ram[1320]) );
  DFFPOSX1 ram_reg_11__24_ ( .D(n5988), .CLK(clk), .Q(ram[1319]) );
  DFFPOSX1 ram_reg_11__25_ ( .D(n5987), .CLK(clk), .Q(ram[1318]) );
  DFFPOSX1 ram_reg_11__26_ ( .D(n5986), .CLK(clk), .Q(ram[1317]) );
  DFFPOSX1 ram_reg_11__27_ ( .D(n5985), .CLK(clk), .Q(ram[1316]) );
  DFFPOSX1 ram_reg_11__28_ ( .D(n5984), .CLK(clk), .Q(ram[1315]) );
  DFFPOSX1 ram_reg_11__29_ ( .D(n5983), .CLK(clk), .Q(ram[1314]) );
  DFFPOSX1 ram_reg_11__30_ ( .D(n5982), .CLK(clk), .Q(ram[1313]) );
  DFFPOSX1 ram_reg_11__31_ ( .D(n5981), .CLK(clk), .Q(ram[1312]) );
  DFFPOSX1 ram_reg_11__32_ ( .D(n5980), .CLK(clk), .Q(ram[1311]) );
  DFFPOSX1 ram_reg_11__33_ ( .D(n5979), .CLK(clk), .Q(ram[1310]) );
  DFFPOSX1 ram_reg_11__34_ ( .D(n5978), .CLK(clk), .Q(ram[1309]) );
  DFFPOSX1 ram_reg_11__35_ ( .D(n5977), .CLK(clk), .Q(ram[1308]) );
  DFFPOSX1 ram_reg_11__36_ ( .D(n5976), .CLK(clk), .Q(ram[1307]) );
  DFFPOSX1 ram_reg_11__37_ ( .D(n5975), .CLK(clk), .Q(ram[1306]) );
  DFFPOSX1 ram_reg_11__38_ ( .D(n5974), .CLK(clk), .Q(ram[1305]) );
  DFFPOSX1 ram_reg_11__39_ ( .D(n5973), .CLK(clk), .Q(ram[1304]) );
  DFFPOSX1 ram_reg_11__40_ ( .D(n5972), .CLK(clk), .Q(ram[1303]) );
  DFFPOSX1 ram_reg_11__41_ ( .D(n5971), .CLK(clk), .Q(ram[1302]) );
  DFFPOSX1 ram_reg_11__42_ ( .D(n5970), .CLK(clk), .Q(ram[1301]) );
  DFFPOSX1 ram_reg_11__43_ ( .D(n5969), .CLK(clk), .Q(ram[1300]) );
  DFFPOSX1 ram_reg_11__44_ ( .D(n5968), .CLK(clk), .Q(ram[1299]) );
  DFFPOSX1 ram_reg_11__45_ ( .D(n5967), .CLK(clk), .Q(ram[1298]) );
  DFFPOSX1 ram_reg_11__46_ ( .D(n5966), .CLK(clk), .Q(ram[1297]) );
  DFFPOSX1 ram_reg_11__47_ ( .D(n5965), .CLK(clk), .Q(ram[1296]) );
  DFFPOSX1 ram_reg_11__48_ ( .D(n5964), .CLK(clk), .Q(ram[1295]) );
  DFFPOSX1 ram_reg_11__49_ ( .D(n5963), .CLK(clk), .Q(ram[1294]) );
  DFFPOSX1 ram_reg_11__50_ ( .D(n5962), .CLK(clk), .Q(ram[1293]) );
  DFFPOSX1 ram_reg_11__51_ ( .D(n5961), .CLK(clk), .Q(ram[1292]) );
  DFFPOSX1 ram_reg_11__52_ ( .D(n5960), .CLK(clk), .Q(ram[1291]) );
  DFFPOSX1 ram_reg_11__53_ ( .D(n5959), .CLK(clk), .Q(ram[1290]) );
  DFFPOSX1 ram_reg_11__54_ ( .D(n5958), .CLK(clk), .Q(ram[1289]) );
  DFFPOSX1 ram_reg_11__55_ ( .D(n5957), .CLK(clk), .Q(ram[1288]) );
  DFFPOSX1 ram_reg_11__56_ ( .D(n5956), .CLK(clk), .Q(ram[1287]) );
  DFFPOSX1 ram_reg_11__57_ ( .D(n5955), .CLK(clk), .Q(ram[1286]) );
  DFFPOSX1 ram_reg_11__58_ ( .D(n5954), .CLK(clk), .Q(ram[1285]) );
  DFFPOSX1 ram_reg_11__59_ ( .D(n5953), .CLK(clk), .Q(ram[1284]) );
  DFFPOSX1 ram_reg_11__60_ ( .D(n5952), .CLK(clk), .Q(ram[1283]) );
  DFFPOSX1 ram_reg_11__61_ ( .D(n5951), .CLK(clk), .Q(ram[1282]) );
  DFFPOSX1 ram_reg_11__62_ ( .D(n5950), .CLK(clk), .Q(ram[1281]) );
  DFFPOSX1 ram_reg_11__63_ ( .D(n5949), .CLK(clk), .Q(ram[1280]) );
  DFFPOSX1 ram_reg_12__0_ ( .D(n5948), .CLK(clk), .Q(ram[1279]) );
  DFFPOSX1 ram_reg_12__1_ ( .D(n5947), .CLK(clk), .Q(ram[1278]) );
  DFFPOSX1 ram_reg_12__2_ ( .D(n5946), .CLK(clk), .Q(ram[1277]) );
  DFFPOSX1 ram_reg_12__3_ ( .D(n5945), .CLK(clk), .Q(ram[1276]) );
  DFFPOSX1 ram_reg_12__4_ ( .D(n5944), .CLK(clk), .Q(ram[1275]) );
  DFFPOSX1 ram_reg_12__5_ ( .D(n5943), .CLK(clk), .Q(ram[1274]) );
  DFFPOSX1 ram_reg_12__6_ ( .D(n5942), .CLK(clk), .Q(ram[1273]) );
  DFFPOSX1 ram_reg_12__7_ ( .D(n5941), .CLK(clk), .Q(ram[1272]) );
  DFFPOSX1 ram_reg_12__8_ ( .D(n5940), .CLK(clk), .Q(ram[1271]) );
  DFFPOSX1 ram_reg_12__9_ ( .D(n5939), .CLK(clk), .Q(ram[1270]) );
  DFFPOSX1 ram_reg_12__10_ ( .D(n5938), .CLK(clk), .Q(ram[1269]) );
  DFFPOSX1 ram_reg_12__11_ ( .D(n5937), .CLK(clk), .Q(ram[1268]) );
  DFFPOSX1 ram_reg_12__12_ ( .D(n5936), .CLK(clk), .Q(ram[1267]) );
  DFFPOSX1 ram_reg_12__13_ ( .D(n5935), .CLK(clk), .Q(ram[1266]) );
  DFFPOSX1 ram_reg_12__14_ ( .D(n5934), .CLK(clk), .Q(ram[1265]) );
  DFFPOSX1 ram_reg_12__15_ ( .D(n5933), .CLK(clk), .Q(ram[1264]) );
  DFFPOSX1 ram_reg_12__16_ ( .D(n5932), .CLK(clk), .Q(ram[1263]) );
  DFFPOSX1 ram_reg_12__17_ ( .D(n5931), .CLK(clk), .Q(ram[1262]) );
  DFFPOSX1 ram_reg_12__18_ ( .D(n5930), .CLK(clk), .Q(ram[1261]) );
  DFFPOSX1 ram_reg_12__19_ ( .D(n5929), .CLK(clk), .Q(ram[1260]) );
  DFFPOSX1 ram_reg_12__20_ ( .D(n5928), .CLK(clk), .Q(ram[1259]) );
  DFFPOSX1 ram_reg_12__21_ ( .D(n5927), .CLK(clk), .Q(ram[1258]) );
  DFFPOSX1 ram_reg_12__22_ ( .D(n5926), .CLK(clk), .Q(ram[1257]) );
  DFFPOSX1 ram_reg_12__23_ ( .D(n5925), .CLK(clk), .Q(ram[1256]) );
  DFFPOSX1 ram_reg_12__24_ ( .D(n5924), .CLK(clk), .Q(ram[1255]) );
  DFFPOSX1 ram_reg_12__25_ ( .D(n5923), .CLK(clk), .Q(ram[1254]) );
  DFFPOSX1 ram_reg_12__26_ ( .D(n5922), .CLK(clk), .Q(ram[1253]) );
  DFFPOSX1 ram_reg_12__27_ ( .D(n5921), .CLK(clk), .Q(ram[1252]) );
  DFFPOSX1 ram_reg_12__28_ ( .D(n5920), .CLK(clk), .Q(ram[1251]) );
  DFFPOSX1 ram_reg_12__29_ ( .D(n5919), .CLK(clk), .Q(ram[1250]) );
  DFFPOSX1 ram_reg_12__30_ ( .D(n5918), .CLK(clk), .Q(ram[1249]) );
  DFFPOSX1 ram_reg_12__31_ ( .D(n5917), .CLK(clk), .Q(ram[1248]) );
  DFFPOSX1 ram_reg_12__32_ ( .D(n5916), .CLK(clk), .Q(ram[1247]) );
  DFFPOSX1 ram_reg_12__33_ ( .D(n5915), .CLK(clk), .Q(ram[1246]) );
  DFFPOSX1 ram_reg_12__34_ ( .D(n5914), .CLK(clk), .Q(ram[1245]) );
  DFFPOSX1 ram_reg_12__35_ ( .D(n5913), .CLK(clk), .Q(ram[1244]) );
  DFFPOSX1 ram_reg_12__36_ ( .D(n5912), .CLK(clk), .Q(ram[1243]) );
  DFFPOSX1 ram_reg_12__37_ ( .D(n5911), .CLK(clk), .Q(ram[1242]) );
  DFFPOSX1 ram_reg_12__38_ ( .D(n5910), .CLK(clk), .Q(ram[1241]) );
  DFFPOSX1 ram_reg_12__39_ ( .D(n5909), .CLK(clk), .Q(ram[1240]) );
  DFFPOSX1 ram_reg_12__40_ ( .D(n5908), .CLK(clk), .Q(ram[1239]) );
  DFFPOSX1 ram_reg_12__41_ ( .D(n5907), .CLK(clk), .Q(ram[1238]) );
  DFFPOSX1 ram_reg_12__42_ ( .D(n5906), .CLK(clk), .Q(ram[1237]) );
  DFFPOSX1 ram_reg_12__43_ ( .D(n5905), .CLK(clk), .Q(ram[1236]) );
  DFFPOSX1 ram_reg_12__44_ ( .D(n5904), .CLK(clk), .Q(ram[1235]) );
  DFFPOSX1 ram_reg_12__45_ ( .D(n5903), .CLK(clk), .Q(ram[1234]) );
  DFFPOSX1 ram_reg_12__46_ ( .D(n5902), .CLK(clk), .Q(ram[1233]) );
  DFFPOSX1 ram_reg_12__47_ ( .D(n5901), .CLK(clk), .Q(ram[1232]) );
  DFFPOSX1 ram_reg_12__48_ ( .D(n5900), .CLK(clk), .Q(ram[1231]) );
  DFFPOSX1 ram_reg_12__49_ ( .D(n5899), .CLK(clk), .Q(ram[1230]) );
  DFFPOSX1 ram_reg_12__50_ ( .D(n5898), .CLK(clk), .Q(ram[1229]) );
  DFFPOSX1 ram_reg_12__51_ ( .D(n5897), .CLK(clk), .Q(ram[1228]) );
  DFFPOSX1 ram_reg_12__52_ ( .D(n5896), .CLK(clk), .Q(ram[1227]) );
  DFFPOSX1 ram_reg_12__53_ ( .D(n5895), .CLK(clk), .Q(ram[1226]) );
  DFFPOSX1 ram_reg_12__54_ ( .D(n5894), .CLK(clk), .Q(ram[1225]) );
  DFFPOSX1 ram_reg_12__55_ ( .D(n5893), .CLK(clk), .Q(ram[1224]) );
  DFFPOSX1 ram_reg_12__56_ ( .D(n5892), .CLK(clk), .Q(ram[1223]) );
  DFFPOSX1 ram_reg_12__57_ ( .D(n5891), .CLK(clk), .Q(ram[1222]) );
  DFFPOSX1 ram_reg_12__58_ ( .D(n5890), .CLK(clk), .Q(ram[1221]) );
  DFFPOSX1 ram_reg_12__59_ ( .D(n5889), .CLK(clk), .Q(ram[1220]) );
  DFFPOSX1 ram_reg_12__60_ ( .D(n5888), .CLK(clk), .Q(ram[1219]) );
  DFFPOSX1 ram_reg_12__61_ ( .D(n5887), .CLK(clk), .Q(ram[1218]) );
  DFFPOSX1 ram_reg_12__62_ ( .D(n5886), .CLK(clk), .Q(ram[1217]) );
  DFFPOSX1 ram_reg_12__63_ ( .D(n5885), .CLK(clk), .Q(ram[1216]) );
  DFFPOSX1 ram_reg_13__0_ ( .D(n5884), .CLK(clk), .Q(ram[1215]) );
  DFFPOSX1 ram_reg_13__1_ ( .D(n5883), .CLK(clk), .Q(ram[1214]) );
  DFFPOSX1 ram_reg_13__2_ ( .D(n5882), .CLK(clk), .Q(ram[1213]) );
  DFFPOSX1 ram_reg_13__3_ ( .D(n5881), .CLK(clk), .Q(ram[1212]) );
  DFFPOSX1 ram_reg_13__4_ ( .D(n5880), .CLK(clk), .Q(ram[1211]) );
  DFFPOSX1 ram_reg_13__5_ ( .D(n5879), .CLK(clk), .Q(ram[1210]) );
  DFFPOSX1 ram_reg_13__6_ ( .D(n5878), .CLK(clk), .Q(ram[1209]) );
  DFFPOSX1 ram_reg_13__7_ ( .D(n5877), .CLK(clk), .Q(ram[1208]) );
  DFFPOSX1 ram_reg_13__8_ ( .D(n5876), .CLK(clk), .Q(ram[1207]) );
  DFFPOSX1 ram_reg_13__9_ ( .D(n5875), .CLK(clk), .Q(ram[1206]) );
  DFFPOSX1 ram_reg_13__10_ ( .D(n5874), .CLK(clk), .Q(ram[1205]) );
  DFFPOSX1 ram_reg_13__11_ ( .D(n5873), .CLK(clk), .Q(ram[1204]) );
  DFFPOSX1 ram_reg_13__12_ ( .D(n5872), .CLK(clk), .Q(ram[1203]) );
  DFFPOSX1 ram_reg_13__13_ ( .D(n5871), .CLK(clk), .Q(ram[1202]) );
  DFFPOSX1 ram_reg_13__14_ ( .D(n5870), .CLK(clk), .Q(ram[1201]) );
  DFFPOSX1 ram_reg_13__15_ ( .D(n5869), .CLK(clk), .Q(ram[1200]) );
  DFFPOSX1 ram_reg_13__16_ ( .D(n5868), .CLK(clk), .Q(ram[1199]) );
  DFFPOSX1 ram_reg_13__17_ ( .D(n5867), .CLK(clk), .Q(ram[1198]) );
  DFFPOSX1 ram_reg_13__18_ ( .D(n5866), .CLK(clk), .Q(ram[1197]) );
  DFFPOSX1 ram_reg_13__19_ ( .D(n5865), .CLK(clk), .Q(ram[1196]) );
  DFFPOSX1 ram_reg_13__20_ ( .D(n5864), .CLK(clk), .Q(ram[1195]) );
  DFFPOSX1 ram_reg_13__21_ ( .D(n5863), .CLK(clk), .Q(ram[1194]) );
  DFFPOSX1 ram_reg_13__22_ ( .D(n5862), .CLK(clk), .Q(ram[1193]) );
  DFFPOSX1 ram_reg_13__23_ ( .D(n5861), .CLK(clk), .Q(ram[1192]) );
  DFFPOSX1 ram_reg_13__24_ ( .D(n5860), .CLK(clk), .Q(ram[1191]) );
  DFFPOSX1 ram_reg_13__25_ ( .D(n5859), .CLK(clk), .Q(ram[1190]) );
  DFFPOSX1 ram_reg_13__26_ ( .D(n5858), .CLK(clk), .Q(ram[1189]) );
  DFFPOSX1 ram_reg_13__27_ ( .D(n5857), .CLK(clk), .Q(ram[1188]) );
  DFFPOSX1 ram_reg_13__28_ ( .D(n5856), .CLK(clk), .Q(ram[1187]) );
  DFFPOSX1 ram_reg_13__29_ ( .D(n5855), .CLK(clk), .Q(ram[1186]) );
  DFFPOSX1 ram_reg_13__30_ ( .D(n5854), .CLK(clk), .Q(ram[1185]) );
  DFFPOSX1 ram_reg_13__31_ ( .D(n5853), .CLK(clk), .Q(ram[1184]) );
  DFFPOSX1 ram_reg_13__32_ ( .D(n5852), .CLK(clk), .Q(ram[1183]) );
  DFFPOSX1 ram_reg_13__33_ ( .D(n5851), .CLK(clk), .Q(ram[1182]) );
  DFFPOSX1 ram_reg_13__34_ ( .D(n5850), .CLK(clk), .Q(ram[1181]) );
  DFFPOSX1 ram_reg_13__35_ ( .D(n5849), .CLK(clk), .Q(ram[1180]) );
  DFFPOSX1 ram_reg_13__36_ ( .D(n5848), .CLK(clk), .Q(ram[1179]) );
  DFFPOSX1 ram_reg_13__37_ ( .D(n5847), .CLK(clk), .Q(ram[1178]) );
  DFFPOSX1 ram_reg_13__38_ ( .D(n5846), .CLK(clk), .Q(ram[1177]) );
  DFFPOSX1 ram_reg_13__39_ ( .D(n5845), .CLK(clk), .Q(ram[1176]) );
  DFFPOSX1 ram_reg_13__40_ ( .D(n5844), .CLK(clk), .Q(ram[1175]) );
  DFFPOSX1 ram_reg_13__41_ ( .D(n5843), .CLK(clk), .Q(ram[1174]) );
  DFFPOSX1 ram_reg_13__42_ ( .D(n5842), .CLK(clk), .Q(ram[1173]) );
  DFFPOSX1 ram_reg_13__43_ ( .D(n5841), .CLK(clk), .Q(ram[1172]) );
  DFFPOSX1 ram_reg_13__44_ ( .D(n5840), .CLK(clk), .Q(ram[1171]) );
  DFFPOSX1 ram_reg_13__45_ ( .D(n5839), .CLK(clk), .Q(ram[1170]) );
  DFFPOSX1 ram_reg_13__46_ ( .D(n5838), .CLK(clk), .Q(ram[1169]) );
  DFFPOSX1 ram_reg_13__47_ ( .D(n5837), .CLK(clk), .Q(ram[1168]) );
  DFFPOSX1 ram_reg_13__48_ ( .D(n5836), .CLK(clk), .Q(ram[1167]) );
  DFFPOSX1 ram_reg_13__49_ ( .D(n5835), .CLK(clk), .Q(ram[1166]) );
  DFFPOSX1 ram_reg_13__50_ ( .D(n5834), .CLK(clk), .Q(ram[1165]) );
  DFFPOSX1 ram_reg_13__51_ ( .D(n5833), .CLK(clk), .Q(ram[1164]) );
  DFFPOSX1 ram_reg_13__52_ ( .D(n5832), .CLK(clk), .Q(ram[1163]) );
  DFFPOSX1 ram_reg_13__53_ ( .D(n5831), .CLK(clk), .Q(ram[1162]) );
  DFFPOSX1 ram_reg_13__54_ ( .D(n5830), .CLK(clk), .Q(ram[1161]) );
  DFFPOSX1 ram_reg_13__55_ ( .D(n5829), .CLK(clk), .Q(ram[1160]) );
  DFFPOSX1 ram_reg_13__56_ ( .D(n5828), .CLK(clk), .Q(ram[1159]) );
  DFFPOSX1 ram_reg_13__57_ ( .D(n5827), .CLK(clk), .Q(ram[1158]) );
  DFFPOSX1 ram_reg_13__58_ ( .D(n5826), .CLK(clk), .Q(ram[1157]) );
  DFFPOSX1 ram_reg_13__59_ ( .D(n5825), .CLK(clk), .Q(ram[1156]) );
  DFFPOSX1 ram_reg_13__60_ ( .D(n5824), .CLK(clk), .Q(ram[1155]) );
  DFFPOSX1 ram_reg_13__61_ ( .D(n5823), .CLK(clk), .Q(ram[1154]) );
  DFFPOSX1 ram_reg_13__62_ ( .D(n5822), .CLK(clk), .Q(ram[1153]) );
  DFFPOSX1 ram_reg_13__63_ ( .D(n5821), .CLK(clk), .Q(ram[1152]) );
  DFFPOSX1 ram_reg_14__0_ ( .D(n5820), .CLK(clk), .Q(ram[1151]) );
  DFFPOSX1 ram_reg_14__1_ ( .D(n5819), .CLK(clk), .Q(ram[1150]) );
  DFFPOSX1 ram_reg_14__2_ ( .D(n5818), .CLK(clk), .Q(ram[1149]) );
  DFFPOSX1 ram_reg_14__3_ ( .D(n5817), .CLK(clk), .Q(ram[1148]) );
  DFFPOSX1 ram_reg_14__4_ ( .D(n5816), .CLK(clk), .Q(ram[1147]) );
  DFFPOSX1 ram_reg_14__5_ ( .D(n5815), .CLK(clk), .Q(ram[1146]) );
  DFFPOSX1 ram_reg_14__6_ ( .D(n5814), .CLK(clk), .Q(ram[1145]) );
  DFFPOSX1 ram_reg_14__7_ ( .D(n5813), .CLK(clk), .Q(ram[1144]) );
  DFFPOSX1 ram_reg_14__8_ ( .D(n5812), .CLK(clk), .Q(ram[1143]) );
  DFFPOSX1 ram_reg_14__9_ ( .D(n5811), .CLK(clk), .Q(ram[1142]) );
  DFFPOSX1 ram_reg_14__10_ ( .D(n5810), .CLK(clk), .Q(ram[1141]) );
  DFFPOSX1 ram_reg_14__11_ ( .D(n5809), .CLK(clk), .Q(ram[1140]) );
  DFFPOSX1 ram_reg_14__12_ ( .D(n5808), .CLK(clk), .Q(ram[1139]) );
  DFFPOSX1 ram_reg_14__13_ ( .D(n5807), .CLK(clk), .Q(ram[1138]) );
  DFFPOSX1 ram_reg_14__14_ ( .D(n5806), .CLK(clk), .Q(ram[1137]) );
  DFFPOSX1 ram_reg_14__15_ ( .D(n5805), .CLK(clk), .Q(ram[1136]) );
  DFFPOSX1 ram_reg_14__16_ ( .D(n5804), .CLK(clk), .Q(ram[1135]) );
  DFFPOSX1 ram_reg_14__17_ ( .D(n5803), .CLK(clk), .Q(ram[1134]) );
  DFFPOSX1 ram_reg_14__18_ ( .D(n5802), .CLK(clk), .Q(ram[1133]) );
  DFFPOSX1 ram_reg_14__19_ ( .D(n5801), .CLK(clk), .Q(ram[1132]) );
  DFFPOSX1 ram_reg_14__20_ ( .D(n5800), .CLK(clk), .Q(ram[1131]) );
  DFFPOSX1 ram_reg_14__21_ ( .D(n5799), .CLK(clk), .Q(ram[1130]) );
  DFFPOSX1 ram_reg_14__22_ ( .D(n5798), .CLK(clk), .Q(ram[1129]) );
  DFFPOSX1 ram_reg_14__23_ ( .D(n5797), .CLK(clk), .Q(ram[1128]) );
  DFFPOSX1 ram_reg_14__24_ ( .D(n5796), .CLK(clk), .Q(ram[1127]) );
  DFFPOSX1 ram_reg_14__25_ ( .D(n5795), .CLK(clk), .Q(ram[1126]) );
  DFFPOSX1 ram_reg_14__26_ ( .D(n5794), .CLK(clk), .Q(ram[1125]) );
  DFFPOSX1 ram_reg_14__27_ ( .D(n5793), .CLK(clk), .Q(ram[1124]) );
  DFFPOSX1 ram_reg_14__28_ ( .D(n5792), .CLK(clk), .Q(ram[1123]) );
  DFFPOSX1 ram_reg_14__29_ ( .D(n5791), .CLK(clk), .Q(ram[1122]) );
  DFFPOSX1 ram_reg_14__30_ ( .D(n5790), .CLK(clk), .Q(ram[1121]) );
  DFFPOSX1 ram_reg_14__31_ ( .D(n5789), .CLK(clk), .Q(ram[1120]) );
  DFFPOSX1 ram_reg_14__32_ ( .D(n5788), .CLK(clk), .Q(ram[1119]) );
  DFFPOSX1 ram_reg_14__33_ ( .D(n5787), .CLK(clk), .Q(ram[1118]) );
  DFFPOSX1 ram_reg_14__34_ ( .D(n5786), .CLK(clk), .Q(ram[1117]) );
  DFFPOSX1 ram_reg_14__35_ ( .D(n5785), .CLK(clk), .Q(ram[1116]) );
  DFFPOSX1 ram_reg_14__36_ ( .D(n5784), .CLK(clk), .Q(ram[1115]) );
  DFFPOSX1 ram_reg_14__37_ ( .D(n5783), .CLK(clk), .Q(ram[1114]) );
  DFFPOSX1 ram_reg_14__38_ ( .D(n5782), .CLK(clk), .Q(ram[1113]) );
  DFFPOSX1 ram_reg_14__39_ ( .D(n5781), .CLK(clk), .Q(ram[1112]) );
  DFFPOSX1 ram_reg_14__40_ ( .D(n5780), .CLK(clk), .Q(ram[1111]) );
  DFFPOSX1 ram_reg_14__41_ ( .D(n5779), .CLK(clk), .Q(ram[1110]) );
  DFFPOSX1 ram_reg_14__42_ ( .D(n5778), .CLK(clk), .Q(ram[1109]) );
  DFFPOSX1 ram_reg_14__43_ ( .D(n5777), .CLK(clk), .Q(ram[1108]) );
  DFFPOSX1 ram_reg_14__44_ ( .D(n5776), .CLK(clk), .Q(ram[1107]) );
  DFFPOSX1 ram_reg_14__45_ ( .D(n5775), .CLK(clk), .Q(ram[1106]) );
  DFFPOSX1 ram_reg_14__46_ ( .D(n5774), .CLK(clk), .Q(ram[1105]) );
  DFFPOSX1 ram_reg_14__47_ ( .D(n5773), .CLK(clk), .Q(ram[1104]) );
  DFFPOSX1 ram_reg_14__48_ ( .D(n5772), .CLK(clk), .Q(ram[1103]) );
  DFFPOSX1 ram_reg_14__49_ ( .D(n5771), .CLK(clk), .Q(ram[1102]) );
  DFFPOSX1 ram_reg_14__50_ ( .D(n5770), .CLK(clk), .Q(ram[1101]) );
  DFFPOSX1 ram_reg_14__51_ ( .D(n5769), .CLK(clk), .Q(ram[1100]) );
  DFFPOSX1 ram_reg_14__52_ ( .D(n5768), .CLK(clk), .Q(ram[1099]) );
  DFFPOSX1 ram_reg_14__53_ ( .D(n5767), .CLK(clk), .Q(ram[1098]) );
  DFFPOSX1 ram_reg_14__54_ ( .D(n5766), .CLK(clk), .Q(ram[1097]) );
  DFFPOSX1 ram_reg_14__55_ ( .D(n5765), .CLK(clk), .Q(ram[1096]) );
  DFFPOSX1 ram_reg_14__56_ ( .D(n5764), .CLK(clk), .Q(ram[1095]) );
  DFFPOSX1 ram_reg_14__57_ ( .D(n5763), .CLK(clk), .Q(ram[1094]) );
  DFFPOSX1 ram_reg_14__58_ ( .D(n5762), .CLK(clk), .Q(ram[1093]) );
  DFFPOSX1 ram_reg_14__59_ ( .D(n5761), .CLK(clk), .Q(ram[1092]) );
  DFFPOSX1 ram_reg_14__60_ ( .D(n5760), .CLK(clk), .Q(ram[1091]) );
  DFFPOSX1 ram_reg_14__61_ ( .D(n5759), .CLK(clk), .Q(ram[1090]) );
  DFFPOSX1 ram_reg_14__62_ ( .D(n5758), .CLK(clk), .Q(ram[1089]) );
  DFFPOSX1 ram_reg_14__63_ ( .D(n5757), .CLK(clk), .Q(ram[1088]) );
  DFFPOSX1 ram_reg_15__0_ ( .D(n5756), .CLK(clk), .Q(ram[1087]) );
  DFFPOSX1 ram_reg_15__1_ ( .D(n5755), .CLK(clk), .Q(ram[1086]) );
  DFFPOSX1 ram_reg_15__2_ ( .D(n5754), .CLK(clk), .Q(ram[1085]) );
  DFFPOSX1 ram_reg_15__3_ ( .D(n5753), .CLK(clk), .Q(ram[1084]) );
  DFFPOSX1 ram_reg_15__4_ ( .D(n5752), .CLK(clk), .Q(ram[1083]) );
  DFFPOSX1 ram_reg_15__5_ ( .D(n5751), .CLK(clk), .Q(ram[1082]) );
  DFFPOSX1 ram_reg_15__6_ ( .D(n5750), .CLK(clk), .Q(ram[1081]) );
  DFFPOSX1 ram_reg_15__7_ ( .D(n5749), .CLK(clk), .Q(ram[1080]) );
  DFFPOSX1 ram_reg_15__8_ ( .D(n5748), .CLK(clk), .Q(ram[1079]) );
  DFFPOSX1 ram_reg_15__9_ ( .D(n5747), .CLK(clk), .Q(ram[1078]) );
  DFFPOSX1 ram_reg_15__10_ ( .D(n5746), .CLK(clk), .Q(ram[1077]) );
  DFFPOSX1 ram_reg_15__11_ ( .D(n5745), .CLK(clk), .Q(ram[1076]) );
  DFFPOSX1 ram_reg_15__12_ ( .D(n5744), .CLK(clk), .Q(ram[1075]) );
  DFFPOSX1 ram_reg_15__13_ ( .D(n5743), .CLK(clk), .Q(ram[1074]) );
  DFFPOSX1 ram_reg_15__14_ ( .D(n5742), .CLK(clk), .Q(ram[1073]) );
  DFFPOSX1 ram_reg_15__15_ ( .D(n5741), .CLK(clk), .Q(ram[1072]) );
  DFFPOSX1 ram_reg_15__16_ ( .D(n5740), .CLK(clk), .Q(ram[1071]) );
  DFFPOSX1 ram_reg_15__17_ ( .D(n5739), .CLK(clk), .Q(ram[1070]) );
  DFFPOSX1 ram_reg_15__18_ ( .D(n5738), .CLK(clk), .Q(ram[1069]) );
  DFFPOSX1 ram_reg_15__19_ ( .D(n5737), .CLK(clk), .Q(ram[1068]) );
  DFFPOSX1 ram_reg_15__20_ ( .D(n5736), .CLK(clk), .Q(ram[1067]) );
  DFFPOSX1 ram_reg_15__21_ ( .D(n5735), .CLK(clk), .Q(ram[1066]) );
  DFFPOSX1 ram_reg_15__22_ ( .D(n5734), .CLK(clk), .Q(ram[1065]) );
  DFFPOSX1 ram_reg_15__23_ ( .D(n5733), .CLK(clk), .Q(ram[1064]) );
  DFFPOSX1 ram_reg_15__24_ ( .D(n5732), .CLK(clk), .Q(ram[1063]) );
  DFFPOSX1 ram_reg_15__25_ ( .D(n5731), .CLK(clk), .Q(ram[1062]) );
  DFFPOSX1 ram_reg_15__26_ ( .D(n5730), .CLK(clk), .Q(ram[1061]) );
  DFFPOSX1 ram_reg_15__27_ ( .D(n5729), .CLK(clk), .Q(ram[1060]) );
  DFFPOSX1 ram_reg_15__28_ ( .D(n5728), .CLK(clk), .Q(ram[1059]) );
  DFFPOSX1 ram_reg_15__29_ ( .D(n5727), .CLK(clk), .Q(ram[1058]) );
  DFFPOSX1 ram_reg_15__30_ ( .D(n5726), .CLK(clk), .Q(ram[1057]) );
  DFFPOSX1 ram_reg_15__31_ ( .D(n5725), .CLK(clk), .Q(ram[1056]) );
  DFFPOSX1 ram_reg_15__32_ ( .D(n5724), .CLK(clk), .Q(ram[1055]) );
  DFFPOSX1 ram_reg_15__33_ ( .D(n5723), .CLK(clk), .Q(ram[1054]) );
  DFFPOSX1 ram_reg_15__34_ ( .D(n5722), .CLK(clk), .Q(ram[1053]) );
  DFFPOSX1 ram_reg_15__35_ ( .D(n5721), .CLK(clk), .Q(ram[1052]) );
  DFFPOSX1 ram_reg_15__36_ ( .D(n5720), .CLK(clk), .Q(ram[1051]) );
  DFFPOSX1 ram_reg_15__37_ ( .D(n5719), .CLK(clk), .Q(ram[1050]) );
  DFFPOSX1 ram_reg_15__38_ ( .D(n5718), .CLK(clk), .Q(ram[1049]) );
  DFFPOSX1 ram_reg_15__39_ ( .D(n5717), .CLK(clk), .Q(ram[1048]) );
  DFFPOSX1 ram_reg_15__40_ ( .D(n5716), .CLK(clk), .Q(ram[1047]) );
  DFFPOSX1 ram_reg_15__41_ ( .D(n5715), .CLK(clk), .Q(ram[1046]) );
  DFFPOSX1 ram_reg_15__42_ ( .D(n5714), .CLK(clk), .Q(ram[1045]) );
  DFFPOSX1 ram_reg_15__43_ ( .D(n5713), .CLK(clk), .Q(ram[1044]) );
  DFFPOSX1 ram_reg_15__44_ ( .D(n5712), .CLK(clk), .Q(ram[1043]) );
  DFFPOSX1 ram_reg_15__45_ ( .D(n5711), .CLK(clk), .Q(ram[1042]) );
  DFFPOSX1 ram_reg_15__46_ ( .D(n5710), .CLK(clk), .Q(ram[1041]) );
  DFFPOSX1 ram_reg_15__47_ ( .D(n5709), .CLK(clk), .Q(ram[1040]) );
  DFFPOSX1 ram_reg_15__48_ ( .D(n5708), .CLK(clk), .Q(ram[1039]) );
  DFFPOSX1 ram_reg_15__49_ ( .D(n5707), .CLK(clk), .Q(ram[1038]) );
  DFFPOSX1 ram_reg_15__50_ ( .D(n5706), .CLK(clk), .Q(ram[1037]) );
  DFFPOSX1 ram_reg_15__51_ ( .D(n5705), .CLK(clk), .Q(ram[1036]) );
  DFFPOSX1 ram_reg_15__52_ ( .D(n5704), .CLK(clk), .Q(ram[1035]) );
  DFFPOSX1 ram_reg_15__53_ ( .D(n5703), .CLK(clk), .Q(ram[1034]) );
  DFFPOSX1 ram_reg_15__54_ ( .D(n5702), .CLK(clk), .Q(ram[1033]) );
  DFFPOSX1 ram_reg_15__55_ ( .D(n5701), .CLK(clk), .Q(ram[1032]) );
  DFFPOSX1 ram_reg_15__56_ ( .D(n5700), .CLK(clk), .Q(ram[1031]) );
  DFFPOSX1 ram_reg_15__57_ ( .D(n5699), .CLK(clk), .Q(ram[1030]) );
  DFFPOSX1 ram_reg_15__58_ ( .D(n5698), .CLK(clk), .Q(ram[1029]) );
  DFFPOSX1 ram_reg_15__59_ ( .D(n5697), .CLK(clk), .Q(ram[1028]) );
  DFFPOSX1 ram_reg_15__60_ ( .D(n5696), .CLK(clk), .Q(ram[1027]) );
  DFFPOSX1 ram_reg_15__61_ ( .D(n5695), .CLK(clk), .Q(ram[1026]) );
  DFFPOSX1 ram_reg_15__62_ ( .D(n5694), .CLK(clk), .Q(ram[1025]) );
  DFFPOSX1 ram_reg_15__63_ ( .D(n5693), .CLK(clk), .Q(ram[1024]) );
  DFFPOSX1 ram_reg_16__0_ ( .D(n5692), .CLK(clk), .Q(ram[1023]) );
  DFFPOSX1 ram_reg_16__1_ ( .D(n5691), .CLK(clk), .Q(ram[1022]) );
  DFFPOSX1 ram_reg_16__2_ ( .D(n5690), .CLK(clk), .Q(ram[1021]) );
  DFFPOSX1 ram_reg_16__3_ ( .D(n5689), .CLK(clk), .Q(ram[1020]) );
  DFFPOSX1 ram_reg_16__4_ ( .D(n5688), .CLK(clk), .Q(ram[1019]) );
  DFFPOSX1 ram_reg_16__5_ ( .D(n5687), .CLK(clk), .Q(ram[1018]) );
  DFFPOSX1 ram_reg_16__6_ ( .D(n5686), .CLK(clk), .Q(ram[1017]) );
  DFFPOSX1 ram_reg_16__7_ ( .D(n5685), .CLK(clk), .Q(ram[1016]) );
  DFFPOSX1 ram_reg_16__8_ ( .D(n5684), .CLK(clk), .Q(ram[1015]) );
  DFFPOSX1 ram_reg_16__9_ ( .D(n5683), .CLK(clk), .Q(ram[1014]) );
  DFFPOSX1 ram_reg_16__10_ ( .D(n5682), .CLK(clk), .Q(ram[1013]) );
  DFFPOSX1 ram_reg_16__11_ ( .D(n5681), .CLK(clk), .Q(ram[1012]) );
  DFFPOSX1 ram_reg_16__12_ ( .D(n5680), .CLK(clk), .Q(ram[1011]) );
  DFFPOSX1 ram_reg_16__13_ ( .D(n5679), .CLK(clk), .Q(ram[1010]) );
  DFFPOSX1 ram_reg_16__14_ ( .D(n5678), .CLK(clk), .Q(ram[1009]) );
  DFFPOSX1 ram_reg_16__15_ ( .D(n5677), .CLK(clk), .Q(ram[1008]) );
  DFFPOSX1 ram_reg_16__16_ ( .D(n5676), .CLK(clk), .Q(ram[1007]) );
  DFFPOSX1 ram_reg_16__17_ ( .D(n5675), .CLK(clk), .Q(ram[1006]) );
  DFFPOSX1 ram_reg_16__18_ ( .D(n5674), .CLK(clk), .Q(ram[1005]) );
  DFFPOSX1 ram_reg_16__19_ ( .D(n5673), .CLK(clk), .Q(ram[1004]) );
  DFFPOSX1 ram_reg_16__20_ ( .D(n5672), .CLK(clk), .Q(ram[1003]) );
  DFFPOSX1 ram_reg_16__21_ ( .D(n5671), .CLK(clk), .Q(ram[1002]) );
  DFFPOSX1 ram_reg_16__22_ ( .D(n5670), .CLK(clk), .Q(ram[1001]) );
  DFFPOSX1 ram_reg_16__23_ ( .D(n5669), .CLK(clk), .Q(ram[1000]) );
  DFFPOSX1 ram_reg_16__24_ ( .D(n5668), .CLK(clk), .Q(ram[999]) );
  DFFPOSX1 ram_reg_16__25_ ( .D(n5667), .CLK(clk), .Q(ram[998]) );
  DFFPOSX1 ram_reg_16__26_ ( .D(n5666), .CLK(clk), .Q(ram[997]) );
  DFFPOSX1 ram_reg_16__27_ ( .D(n5665), .CLK(clk), .Q(ram[996]) );
  DFFPOSX1 ram_reg_16__28_ ( .D(n5664), .CLK(clk), .Q(ram[995]) );
  DFFPOSX1 ram_reg_16__29_ ( .D(n5663), .CLK(clk), .Q(ram[994]) );
  DFFPOSX1 ram_reg_16__30_ ( .D(n5662), .CLK(clk), .Q(ram[993]) );
  DFFPOSX1 ram_reg_16__31_ ( .D(n5661), .CLK(clk), .Q(ram[992]) );
  DFFPOSX1 ram_reg_16__32_ ( .D(n5660), .CLK(clk), .Q(ram[991]) );
  DFFPOSX1 ram_reg_16__33_ ( .D(n5659), .CLK(clk), .Q(ram[990]) );
  DFFPOSX1 ram_reg_16__34_ ( .D(n5658), .CLK(clk), .Q(ram[989]) );
  DFFPOSX1 ram_reg_16__35_ ( .D(n5657), .CLK(clk), .Q(ram[988]) );
  DFFPOSX1 ram_reg_16__36_ ( .D(n5656), .CLK(clk), .Q(ram[987]) );
  DFFPOSX1 ram_reg_16__37_ ( .D(n5655), .CLK(clk), .Q(ram[986]) );
  DFFPOSX1 ram_reg_16__38_ ( .D(n5654), .CLK(clk), .Q(ram[985]) );
  DFFPOSX1 ram_reg_16__39_ ( .D(n5653), .CLK(clk), .Q(ram[984]) );
  DFFPOSX1 ram_reg_16__40_ ( .D(n5652), .CLK(clk), .Q(ram[983]) );
  DFFPOSX1 ram_reg_16__41_ ( .D(n5651), .CLK(clk), .Q(ram[982]) );
  DFFPOSX1 ram_reg_16__42_ ( .D(n5650), .CLK(clk), .Q(ram[981]) );
  DFFPOSX1 ram_reg_16__43_ ( .D(n5649), .CLK(clk), .Q(ram[980]) );
  DFFPOSX1 ram_reg_16__44_ ( .D(n5648), .CLK(clk), .Q(ram[979]) );
  DFFPOSX1 ram_reg_16__45_ ( .D(n5647), .CLK(clk), .Q(ram[978]) );
  DFFPOSX1 ram_reg_16__46_ ( .D(n5646), .CLK(clk), .Q(ram[977]) );
  DFFPOSX1 ram_reg_16__47_ ( .D(n5645), .CLK(clk), .Q(ram[976]) );
  DFFPOSX1 ram_reg_16__48_ ( .D(n5644), .CLK(clk), .Q(ram[975]) );
  DFFPOSX1 ram_reg_16__49_ ( .D(n5643), .CLK(clk), .Q(ram[974]) );
  DFFPOSX1 ram_reg_16__50_ ( .D(n5642), .CLK(clk), .Q(ram[973]) );
  DFFPOSX1 ram_reg_16__51_ ( .D(n5641), .CLK(clk), .Q(ram[972]) );
  DFFPOSX1 ram_reg_16__52_ ( .D(n5640), .CLK(clk), .Q(ram[971]) );
  DFFPOSX1 ram_reg_16__53_ ( .D(n5639), .CLK(clk), .Q(ram[970]) );
  DFFPOSX1 ram_reg_16__54_ ( .D(n5638), .CLK(clk), .Q(ram[969]) );
  DFFPOSX1 ram_reg_16__55_ ( .D(n5637), .CLK(clk), .Q(ram[968]) );
  DFFPOSX1 ram_reg_16__56_ ( .D(n5636), .CLK(clk), .Q(ram[967]) );
  DFFPOSX1 ram_reg_16__57_ ( .D(n5635), .CLK(clk), .Q(ram[966]) );
  DFFPOSX1 ram_reg_16__58_ ( .D(n5634), .CLK(clk), .Q(ram[965]) );
  DFFPOSX1 ram_reg_16__59_ ( .D(n5633), .CLK(clk), .Q(ram[964]) );
  DFFPOSX1 ram_reg_16__60_ ( .D(n5632), .CLK(clk), .Q(ram[963]) );
  DFFPOSX1 ram_reg_16__61_ ( .D(n5631), .CLK(clk), .Q(ram[962]) );
  DFFPOSX1 ram_reg_16__62_ ( .D(n5630), .CLK(clk), .Q(ram[961]) );
  DFFPOSX1 ram_reg_16__63_ ( .D(n5629), .CLK(clk), .Q(ram[960]) );
  DFFPOSX1 ram_reg_17__0_ ( .D(n5628), .CLK(clk), .Q(ram[959]) );
  DFFPOSX1 ram_reg_17__1_ ( .D(n5627), .CLK(clk), .Q(ram[958]) );
  DFFPOSX1 ram_reg_17__2_ ( .D(n5626), .CLK(clk), .Q(ram[957]) );
  DFFPOSX1 ram_reg_17__3_ ( .D(n5625), .CLK(clk), .Q(ram[956]) );
  DFFPOSX1 ram_reg_17__4_ ( .D(n5624), .CLK(clk), .Q(ram[955]) );
  DFFPOSX1 ram_reg_17__5_ ( .D(n5623), .CLK(clk), .Q(ram[954]) );
  DFFPOSX1 ram_reg_17__6_ ( .D(n5622), .CLK(clk), .Q(ram[953]) );
  DFFPOSX1 ram_reg_17__7_ ( .D(n5621), .CLK(clk), .Q(ram[952]) );
  DFFPOSX1 ram_reg_17__8_ ( .D(n5620), .CLK(clk), .Q(ram[951]) );
  DFFPOSX1 ram_reg_17__9_ ( .D(n5619), .CLK(clk), .Q(ram[950]) );
  DFFPOSX1 ram_reg_17__10_ ( .D(n5618), .CLK(clk), .Q(ram[949]) );
  DFFPOSX1 ram_reg_17__11_ ( .D(n5617), .CLK(clk), .Q(ram[948]) );
  DFFPOSX1 ram_reg_17__12_ ( .D(n5616), .CLK(clk), .Q(ram[947]) );
  DFFPOSX1 ram_reg_17__13_ ( .D(n5615), .CLK(clk), .Q(ram[946]) );
  DFFPOSX1 ram_reg_17__14_ ( .D(n5614), .CLK(clk), .Q(ram[945]) );
  DFFPOSX1 ram_reg_17__15_ ( .D(n5613), .CLK(clk), .Q(ram[944]) );
  DFFPOSX1 ram_reg_17__16_ ( .D(n5612), .CLK(clk), .Q(ram[943]) );
  DFFPOSX1 ram_reg_17__17_ ( .D(n5611), .CLK(clk), .Q(ram[942]) );
  DFFPOSX1 ram_reg_17__18_ ( .D(n5610), .CLK(clk), .Q(ram[941]) );
  DFFPOSX1 ram_reg_17__19_ ( .D(n5609), .CLK(clk), .Q(ram[940]) );
  DFFPOSX1 ram_reg_17__20_ ( .D(n5608), .CLK(clk), .Q(ram[939]) );
  DFFPOSX1 ram_reg_17__21_ ( .D(n5607), .CLK(clk), .Q(ram[938]) );
  DFFPOSX1 ram_reg_17__22_ ( .D(n5606), .CLK(clk), .Q(ram[937]) );
  DFFPOSX1 ram_reg_17__23_ ( .D(n5605), .CLK(clk), .Q(ram[936]) );
  DFFPOSX1 ram_reg_17__24_ ( .D(n5604), .CLK(clk), .Q(ram[935]) );
  DFFPOSX1 ram_reg_17__25_ ( .D(n5603), .CLK(clk), .Q(ram[934]) );
  DFFPOSX1 ram_reg_17__26_ ( .D(n5602), .CLK(clk), .Q(ram[933]) );
  DFFPOSX1 ram_reg_17__27_ ( .D(n5601), .CLK(clk), .Q(ram[932]) );
  DFFPOSX1 ram_reg_17__28_ ( .D(n5600), .CLK(clk), .Q(ram[931]) );
  DFFPOSX1 ram_reg_17__29_ ( .D(n5599), .CLK(clk), .Q(ram[930]) );
  DFFPOSX1 ram_reg_17__30_ ( .D(n5598), .CLK(clk), .Q(ram[929]) );
  DFFPOSX1 ram_reg_17__31_ ( .D(n5597), .CLK(clk), .Q(ram[928]) );
  DFFPOSX1 ram_reg_17__32_ ( .D(n5596), .CLK(clk), .Q(ram[927]) );
  DFFPOSX1 ram_reg_17__33_ ( .D(n5595), .CLK(clk), .Q(ram[926]) );
  DFFPOSX1 ram_reg_17__34_ ( .D(n5594), .CLK(clk), .Q(ram[925]) );
  DFFPOSX1 ram_reg_17__35_ ( .D(n5593), .CLK(clk), .Q(ram[924]) );
  DFFPOSX1 ram_reg_17__36_ ( .D(n5592), .CLK(clk), .Q(ram[923]) );
  DFFPOSX1 ram_reg_17__37_ ( .D(n5591), .CLK(clk), .Q(ram[922]) );
  DFFPOSX1 ram_reg_17__38_ ( .D(n5590), .CLK(clk), .Q(ram[921]) );
  DFFPOSX1 ram_reg_17__39_ ( .D(n5589), .CLK(clk), .Q(ram[920]) );
  DFFPOSX1 ram_reg_17__40_ ( .D(n5588), .CLK(clk), .Q(ram[919]) );
  DFFPOSX1 ram_reg_17__41_ ( .D(n5587), .CLK(clk), .Q(ram[918]) );
  DFFPOSX1 ram_reg_17__42_ ( .D(n5586), .CLK(clk), .Q(ram[917]) );
  DFFPOSX1 ram_reg_17__43_ ( .D(n5585), .CLK(clk), .Q(ram[916]) );
  DFFPOSX1 ram_reg_17__44_ ( .D(n5584), .CLK(clk), .Q(ram[915]) );
  DFFPOSX1 ram_reg_17__45_ ( .D(n5583), .CLK(clk), .Q(ram[914]) );
  DFFPOSX1 ram_reg_17__46_ ( .D(n5582), .CLK(clk), .Q(ram[913]) );
  DFFPOSX1 ram_reg_17__47_ ( .D(n5581), .CLK(clk), .Q(ram[912]) );
  DFFPOSX1 ram_reg_17__48_ ( .D(n5580), .CLK(clk), .Q(ram[911]) );
  DFFPOSX1 ram_reg_17__49_ ( .D(n5579), .CLK(clk), .Q(ram[910]) );
  DFFPOSX1 ram_reg_17__50_ ( .D(n5578), .CLK(clk), .Q(ram[909]) );
  DFFPOSX1 ram_reg_17__51_ ( .D(n5577), .CLK(clk), .Q(ram[908]) );
  DFFPOSX1 ram_reg_17__52_ ( .D(n5576), .CLK(clk), .Q(ram[907]) );
  DFFPOSX1 ram_reg_17__53_ ( .D(n5575), .CLK(clk), .Q(ram[906]) );
  DFFPOSX1 ram_reg_17__54_ ( .D(n5574), .CLK(clk), .Q(ram[905]) );
  DFFPOSX1 ram_reg_17__55_ ( .D(n5573), .CLK(clk), .Q(ram[904]) );
  DFFPOSX1 ram_reg_17__56_ ( .D(n5572), .CLK(clk), .Q(ram[903]) );
  DFFPOSX1 ram_reg_17__57_ ( .D(n5571), .CLK(clk), .Q(ram[902]) );
  DFFPOSX1 ram_reg_17__58_ ( .D(n5570), .CLK(clk), .Q(ram[901]) );
  DFFPOSX1 ram_reg_17__59_ ( .D(n5569), .CLK(clk), .Q(ram[900]) );
  DFFPOSX1 ram_reg_17__60_ ( .D(n5568), .CLK(clk), .Q(ram[899]) );
  DFFPOSX1 ram_reg_17__61_ ( .D(n5567), .CLK(clk), .Q(ram[898]) );
  DFFPOSX1 ram_reg_17__62_ ( .D(n5566), .CLK(clk), .Q(ram[897]) );
  DFFPOSX1 ram_reg_17__63_ ( .D(n5565), .CLK(clk), .Q(ram[896]) );
  DFFPOSX1 ram_reg_18__0_ ( .D(n5564), .CLK(clk), .Q(ram[895]) );
  DFFPOSX1 ram_reg_18__1_ ( .D(n5563), .CLK(clk), .Q(ram[894]) );
  DFFPOSX1 ram_reg_18__2_ ( .D(n5562), .CLK(clk), .Q(ram[893]) );
  DFFPOSX1 ram_reg_18__3_ ( .D(n5561), .CLK(clk), .Q(ram[892]) );
  DFFPOSX1 ram_reg_18__4_ ( .D(n5560), .CLK(clk), .Q(ram[891]) );
  DFFPOSX1 ram_reg_18__5_ ( .D(n5559), .CLK(clk), .Q(ram[890]) );
  DFFPOSX1 ram_reg_18__6_ ( .D(n5558), .CLK(clk), .Q(ram[889]) );
  DFFPOSX1 ram_reg_18__7_ ( .D(n5557), .CLK(clk), .Q(ram[888]) );
  DFFPOSX1 ram_reg_18__8_ ( .D(n5556), .CLK(clk), .Q(ram[887]) );
  DFFPOSX1 ram_reg_18__9_ ( .D(n5555), .CLK(clk), .Q(ram[886]) );
  DFFPOSX1 ram_reg_18__10_ ( .D(n5554), .CLK(clk), .Q(ram[885]) );
  DFFPOSX1 ram_reg_18__11_ ( .D(n5553), .CLK(clk), .Q(ram[884]) );
  DFFPOSX1 ram_reg_18__12_ ( .D(n5552), .CLK(clk), .Q(ram[883]) );
  DFFPOSX1 ram_reg_18__13_ ( .D(n5551), .CLK(clk), .Q(ram[882]) );
  DFFPOSX1 ram_reg_18__14_ ( .D(n5550), .CLK(clk), .Q(ram[881]) );
  DFFPOSX1 ram_reg_18__15_ ( .D(n5549), .CLK(clk), .Q(ram[880]) );
  DFFPOSX1 ram_reg_18__16_ ( .D(n5548), .CLK(clk), .Q(ram[879]) );
  DFFPOSX1 ram_reg_18__17_ ( .D(n5547), .CLK(clk), .Q(ram[878]) );
  DFFPOSX1 ram_reg_18__18_ ( .D(n5546), .CLK(clk), .Q(ram[877]) );
  DFFPOSX1 ram_reg_18__19_ ( .D(n5545), .CLK(clk), .Q(ram[876]) );
  DFFPOSX1 ram_reg_18__20_ ( .D(n5544), .CLK(clk), .Q(ram[875]) );
  DFFPOSX1 ram_reg_18__21_ ( .D(n5543), .CLK(clk), .Q(ram[874]) );
  DFFPOSX1 ram_reg_18__22_ ( .D(n5542), .CLK(clk), .Q(ram[873]) );
  DFFPOSX1 ram_reg_18__23_ ( .D(n5541), .CLK(clk), .Q(ram[872]) );
  DFFPOSX1 ram_reg_18__24_ ( .D(n5540), .CLK(clk), .Q(ram[871]) );
  DFFPOSX1 ram_reg_18__25_ ( .D(n5539), .CLK(clk), .Q(ram[870]) );
  DFFPOSX1 ram_reg_18__26_ ( .D(n5538), .CLK(clk), .Q(ram[869]) );
  DFFPOSX1 ram_reg_18__27_ ( .D(n5537), .CLK(clk), .Q(ram[868]) );
  DFFPOSX1 ram_reg_18__28_ ( .D(n5536), .CLK(clk), .Q(ram[867]) );
  DFFPOSX1 ram_reg_18__29_ ( .D(n5535), .CLK(clk), .Q(ram[866]) );
  DFFPOSX1 ram_reg_18__30_ ( .D(n5534), .CLK(clk), .Q(ram[865]) );
  DFFPOSX1 ram_reg_18__31_ ( .D(n5533), .CLK(clk), .Q(ram[864]) );
  DFFPOSX1 ram_reg_18__32_ ( .D(n5532), .CLK(clk), .Q(ram[863]) );
  DFFPOSX1 ram_reg_18__33_ ( .D(n5531), .CLK(clk), .Q(ram[862]) );
  DFFPOSX1 ram_reg_18__34_ ( .D(n5530), .CLK(clk), .Q(ram[861]) );
  DFFPOSX1 ram_reg_18__35_ ( .D(n5529), .CLK(clk), .Q(ram[860]) );
  DFFPOSX1 ram_reg_18__36_ ( .D(n5528), .CLK(clk), .Q(ram[859]) );
  DFFPOSX1 ram_reg_18__37_ ( .D(n5527), .CLK(clk), .Q(ram[858]) );
  DFFPOSX1 ram_reg_18__38_ ( .D(n5526), .CLK(clk), .Q(ram[857]) );
  DFFPOSX1 ram_reg_18__39_ ( .D(n5525), .CLK(clk), .Q(ram[856]) );
  DFFPOSX1 ram_reg_18__40_ ( .D(n5524), .CLK(clk), .Q(ram[855]) );
  DFFPOSX1 ram_reg_18__41_ ( .D(n5523), .CLK(clk), .Q(ram[854]) );
  DFFPOSX1 ram_reg_18__42_ ( .D(n5522), .CLK(clk), .Q(ram[853]) );
  DFFPOSX1 ram_reg_18__43_ ( .D(n5521), .CLK(clk), .Q(ram[852]) );
  DFFPOSX1 ram_reg_18__44_ ( .D(n5520), .CLK(clk), .Q(ram[851]) );
  DFFPOSX1 ram_reg_18__45_ ( .D(n5519), .CLK(clk), .Q(ram[850]) );
  DFFPOSX1 ram_reg_18__46_ ( .D(n5518), .CLK(clk), .Q(ram[849]) );
  DFFPOSX1 ram_reg_18__47_ ( .D(n5517), .CLK(clk), .Q(ram[848]) );
  DFFPOSX1 ram_reg_18__48_ ( .D(n5516), .CLK(clk), .Q(ram[847]) );
  DFFPOSX1 ram_reg_18__49_ ( .D(n5515), .CLK(clk), .Q(ram[846]) );
  DFFPOSX1 ram_reg_18__50_ ( .D(n5514), .CLK(clk), .Q(ram[845]) );
  DFFPOSX1 ram_reg_18__51_ ( .D(n5513), .CLK(clk), .Q(ram[844]) );
  DFFPOSX1 ram_reg_18__52_ ( .D(n5512), .CLK(clk), .Q(ram[843]) );
  DFFPOSX1 ram_reg_18__53_ ( .D(n5511), .CLK(clk), .Q(ram[842]) );
  DFFPOSX1 ram_reg_18__54_ ( .D(n5510), .CLK(clk), .Q(ram[841]) );
  DFFPOSX1 ram_reg_18__55_ ( .D(n5509), .CLK(clk), .Q(ram[840]) );
  DFFPOSX1 ram_reg_18__56_ ( .D(n5508), .CLK(clk), .Q(ram[839]) );
  DFFPOSX1 ram_reg_18__57_ ( .D(n5507), .CLK(clk), .Q(ram[838]) );
  DFFPOSX1 ram_reg_18__58_ ( .D(n5506), .CLK(clk), .Q(ram[837]) );
  DFFPOSX1 ram_reg_18__59_ ( .D(n5505), .CLK(clk), .Q(ram[836]) );
  DFFPOSX1 ram_reg_18__60_ ( .D(n5504), .CLK(clk), .Q(ram[835]) );
  DFFPOSX1 ram_reg_18__61_ ( .D(n5503), .CLK(clk), .Q(ram[834]) );
  DFFPOSX1 ram_reg_18__62_ ( .D(n5502), .CLK(clk), .Q(ram[833]) );
  DFFPOSX1 ram_reg_18__63_ ( .D(n5501), .CLK(clk), .Q(ram[832]) );
  DFFPOSX1 ram_reg_19__0_ ( .D(n5500), .CLK(clk), .Q(ram[831]) );
  DFFPOSX1 ram_reg_19__1_ ( .D(n5499), .CLK(clk), .Q(ram[830]) );
  DFFPOSX1 ram_reg_19__2_ ( .D(n5498), .CLK(clk), .Q(ram[829]) );
  DFFPOSX1 ram_reg_19__3_ ( .D(n5497), .CLK(clk), .Q(ram[828]) );
  DFFPOSX1 ram_reg_19__4_ ( .D(n5496), .CLK(clk), .Q(ram[827]) );
  DFFPOSX1 ram_reg_19__5_ ( .D(n5495), .CLK(clk), .Q(ram[826]) );
  DFFPOSX1 ram_reg_19__6_ ( .D(n5494), .CLK(clk), .Q(ram[825]) );
  DFFPOSX1 ram_reg_19__7_ ( .D(n5493), .CLK(clk), .Q(ram[824]) );
  DFFPOSX1 ram_reg_19__8_ ( .D(n5492), .CLK(clk), .Q(ram[823]) );
  DFFPOSX1 ram_reg_19__9_ ( .D(n5491), .CLK(clk), .Q(ram[822]) );
  DFFPOSX1 ram_reg_19__10_ ( .D(n5490), .CLK(clk), .Q(ram[821]) );
  DFFPOSX1 ram_reg_19__11_ ( .D(n5489), .CLK(clk), .Q(ram[820]) );
  DFFPOSX1 ram_reg_19__12_ ( .D(n5488), .CLK(clk), .Q(ram[819]) );
  DFFPOSX1 ram_reg_19__13_ ( .D(n5487), .CLK(clk), .Q(ram[818]) );
  DFFPOSX1 ram_reg_19__14_ ( .D(n5486), .CLK(clk), .Q(ram[817]) );
  DFFPOSX1 ram_reg_19__15_ ( .D(n5485), .CLK(clk), .Q(ram[816]) );
  DFFPOSX1 ram_reg_19__16_ ( .D(n5484), .CLK(clk), .Q(ram[815]) );
  DFFPOSX1 ram_reg_19__17_ ( .D(n5483), .CLK(clk), .Q(ram[814]) );
  DFFPOSX1 ram_reg_19__18_ ( .D(n5482), .CLK(clk), .Q(ram[813]) );
  DFFPOSX1 ram_reg_19__19_ ( .D(n5481), .CLK(clk), .Q(ram[812]) );
  DFFPOSX1 ram_reg_19__20_ ( .D(n5480), .CLK(clk), .Q(ram[811]) );
  DFFPOSX1 ram_reg_19__21_ ( .D(n5479), .CLK(clk), .Q(ram[810]) );
  DFFPOSX1 ram_reg_19__22_ ( .D(n5478), .CLK(clk), .Q(ram[809]) );
  DFFPOSX1 ram_reg_19__23_ ( .D(n5477), .CLK(clk), .Q(ram[808]) );
  DFFPOSX1 ram_reg_19__24_ ( .D(n5476), .CLK(clk), .Q(ram[807]) );
  DFFPOSX1 ram_reg_19__25_ ( .D(n5475), .CLK(clk), .Q(ram[806]) );
  DFFPOSX1 ram_reg_19__26_ ( .D(n5474), .CLK(clk), .Q(ram[805]) );
  DFFPOSX1 ram_reg_19__27_ ( .D(n5473), .CLK(clk), .Q(ram[804]) );
  DFFPOSX1 ram_reg_19__28_ ( .D(n5472), .CLK(clk), .Q(ram[803]) );
  DFFPOSX1 ram_reg_19__29_ ( .D(n5471), .CLK(clk), .Q(ram[802]) );
  DFFPOSX1 ram_reg_19__30_ ( .D(n5470), .CLK(clk), .Q(ram[801]) );
  DFFPOSX1 ram_reg_19__31_ ( .D(n5469), .CLK(clk), .Q(ram[800]) );
  DFFPOSX1 ram_reg_19__32_ ( .D(n5468), .CLK(clk), .Q(ram[799]) );
  DFFPOSX1 ram_reg_19__33_ ( .D(n5467), .CLK(clk), .Q(ram[798]) );
  DFFPOSX1 ram_reg_19__34_ ( .D(n5466), .CLK(clk), .Q(ram[797]) );
  DFFPOSX1 ram_reg_19__35_ ( .D(n5465), .CLK(clk), .Q(ram[796]) );
  DFFPOSX1 ram_reg_19__36_ ( .D(n5464), .CLK(clk), .Q(ram[795]) );
  DFFPOSX1 ram_reg_19__37_ ( .D(n5463), .CLK(clk), .Q(ram[794]) );
  DFFPOSX1 ram_reg_19__38_ ( .D(n5462), .CLK(clk), .Q(ram[793]) );
  DFFPOSX1 ram_reg_19__39_ ( .D(n5461), .CLK(clk), .Q(ram[792]) );
  DFFPOSX1 ram_reg_19__40_ ( .D(n5460), .CLK(clk), .Q(ram[791]) );
  DFFPOSX1 ram_reg_19__41_ ( .D(n5459), .CLK(clk), .Q(ram[790]) );
  DFFPOSX1 ram_reg_19__42_ ( .D(n5458), .CLK(clk), .Q(ram[789]) );
  DFFPOSX1 ram_reg_19__43_ ( .D(n5457), .CLK(clk), .Q(ram[788]) );
  DFFPOSX1 ram_reg_19__44_ ( .D(n5456), .CLK(clk), .Q(ram[787]) );
  DFFPOSX1 ram_reg_19__45_ ( .D(n5455), .CLK(clk), .Q(ram[786]) );
  DFFPOSX1 ram_reg_19__46_ ( .D(n5454), .CLK(clk), .Q(ram[785]) );
  DFFPOSX1 ram_reg_19__47_ ( .D(n5453), .CLK(clk), .Q(ram[784]) );
  DFFPOSX1 ram_reg_19__48_ ( .D(n5452), .CLK(clk), .Q(ram[783]) );
  DFFPOSX1 ram_reg_19__49_ ( .D(n5451), .CLK(clk), .Q(ram[782]) );
  DFFPOSX1 ram_reg_19__50_ ( .D(n5450), .CLK(clk), .Q(ram[781]) );
  DFFPOSX1 ram_reg_19__51_ ( .D(n5449), .CLK(clk), .Q(ram[780]) );
  DFFPOSX1 ram_reg_19__52_ ( .D(n5448), .CLK(clk), .Q(ram[779]) );
  DFFPOSX1 ram_reg_19__53_ ( .D(n5447), .CLK(clk), .Q(ram[778]) );
  DFFPOSX1 ram_reg_19__54_ ( .D(n5446), .CLK(clk), .Q(ram[777]) );
  DFFPOSX1 ram_reg_19__55_ ( .D(n5445), .CLK(clk), .Q(ram[776]) );
  DFFPOSX1 ram_reg_19__56_ ( .D(n5444), .CLK(clk), .Q(ram[775]) );
  DFFPOSX1 ram_reg_19__57_ ( .D(n5443), .CLK(clk), .Q(ram[774]) );
  DFFPOSX1 ram_reg_19__58_ ( .D(n5442), .CLK(clk), .Q(ram[773]) );
  DFFPOSX1 ram_reg_19__59_ ( .D(n5441), .CLK(clk), .Q(ram[772]) );
  DFFPOSX1 ram_reg_19__60_ ( .D(n5440), .CLK(clk), .Q(ram[771]) );
  DFFPOSX1 ram_reg_19__61_ ( .D(n5439), .CLK(clk), .Q(ram[770]) );
  DFFPOSX1 ram_reg_19__62_ ( .D(n5438), .CLK(clk), .Q(ram[769]) );
  DFFPOSX1 ram_reg_19__63_ ( .D(n5437), .CLK(clk), .Q(ram[768]) );
  DFFPOSX1 ram_reg_20__0_ ( .D(n5436), .CLK(clk), .Q(ram[767]) );
  DFFPOSX1 ram_reg_20__1_ ( .D(n5435), .CLK(clk), .Q(ram[766]) );
  DFFPOSX1 ram_reg_20__2_ ( .D(n5434), .CLK(clk), .Q(ram[765]) );
  DFFPOSX1 ram_reg_20__3_ ( .D(n5433), .CLK(clk), .Q(ram[764]) );
  DFFPOSX1 ram_reg_20__4_ ( .D(n5432), .CLK(clk), .Q(ram[763]) );
  DFFPOSX1 ram_reg_20__5_ ( .D(n5431), .CLK(clk), .Q(ram[762]) );
  DFFPOSX1 ram_reg_20__6_ ( .D(n5430), .CLK(clk), .Q(ram[761]) );
  DFFPOSX1 ram_reg_20__7_ ( .D(n5429), .CLK(clk), .Q(ram[760]) );
  DFFPOSX1 ram_reg_20__8_ ( .D(n5428), .CLK(clk), .Q(ram[759]) );
  DFFPOSX1 ram_reg_20__9_ ( .D(n5427), .CLK(clk), .Q(ram[758]) );
  DFFPOSX1 ram_reg_20__10_ ( .D(n5426), .CLK(clk), .Q(ram[757]) );
  DFFPOSX1 ram_reg_20__11_ ( .D(n5425), .CLK(clk), .Q(ram[756]) );
  DFFPOSX1 ram_reg_20__12_ ( .D(n5424), .CLK(clk), .Q(ram[755]) );
  DFFPOSX1 ram_reg_20__13_ ( .D(n5423), .CLK(clk), .Q(ram[754]) );
  DFFPOSX1 ram_reg_20__14_ ( .D(n5422), .CLK(clk), .Q(ram[753]) );
  DFFPOSX1 ram_reg_20__15_ ( .D(n5421), .CLK(clk), .Q(ram[752]) );
  DFFPOSX1 ram_reg_20__16_ ( .D(n5420), .CLK(clk), .Q(ram[751]) );
  DFFPOSX1 ram_reg_20__17_ ( .D(n5419), .CLK(clk), .Q(ram[750]) );
  DFFPOSX1 ram_reg_20__18_ ( .D(n5418), .CLK(clk), .Q(ram[749]) );
  DFFPOSX1 ram_reg_20__19_ ( .D(n5417), .CLK(clk), .Q(ram[748]) );
  DFFPOSX1 ram_reg_20__20_ ( .D(n5416), .CLK(clk), .Q(ram[747]) );
  DFFPOSX1 ram_reg_20__21_ ( .D(n5415), .CLK(clk), .Q(ram[746]) );
  DFFPOSX1 ram_reg_20__22_ ( .D(n5414), .CLK(clk), .Q(ram[745]) );
  DFFPOSX1 ram_reg_20__23_ ( .D(n5413), .CLK(clk), .Q(ram[744]) );
  DFFPOSX1 ram_reg_20__24_ ( .D(n5412), .CLK(clk), .Q(ram[743]) );
  DFFPOSX1 ram_reg_20__25_ ( .D(n5411), .CLK(clk), .Q(ram[742]) );
  DFFPOSX1 ram_reg_20__26_ ( .D(n5410), .CLK(clk), .Q(ram[741]) );
  DFFPOSX1 ram_reg_20__27_ ( .D(n5409), .CLK(clk), .Q(ram[740]) );
  DFFPOSX1 ram_reg_20__28_ ( .D(n5408), .CLK(clk), .Q(ram[739]) );
  DFFPOSX1 ram_reg_20__29_ ( .D(n5407), .CLK(clk), .Q(ram[738]) );
  DFFPOSX1 ram_reg_20__30_ ( .D(n5406), .CLK(clk), .Q(ram[737]) );
  DFFPOSX1 ram_reg_20__31_ ( .D(n5405), .CLK(clk), .Q(ram[736]) );
  DFFPOSX1 ram_reg_20__32_ ( .D(n5404), .CLK(clk), .Q(ram[735]) );
  DFFPOSX1 ram_reg_20__33_ ( .D(n5403), .CLK(clk), .Q(ram[734]) );
  DFFPOSX1 ram_reg_20__34_ ( .D(n5402), .CLK(clk), .Q(ram[733]) );
  DFFPOSX1 ram_reg_20__35_ ( .D(n5401), .CLK(clk), .Q(ram[732]) );
  DFFPOSX1 ram_reg_20__36_ ( .D(n5400), .CLK(clk), .Q(ram[731]) );
  DFFPOSX1 ram_reg_20__37_ ( .D(n5399), .CLK(clk), .Q(ram[730]) );
  DFFPOSX1 ram_reg_20__38_ ( .D(n5398), .CLK(clk), .Q(ram[729]) );
  DFFPOSX1 ram_reg_20__39_ ( .D(n5397), .CLK(clk), .Q(ram[728]) );
  DFFPOSX1 ram_reg_20__40_ ( .D(n5396), .CLK(clk), .Q(ram[727]) );
  DFFPOSX1 ram_reg_20__41_ ( .D(n5395), .CLK(clk), .Q(ram[726]) );
  DFFPOSX1 ram_reg_20__42_ ( .D(n5394), .CLK(clk), .Q(ram[725]) );
  DFFPOSX1 ram_reg_20__43_ ( .D(n5393), .CLK(clk), .Q(ram[724]) );
  DFFPOSX1 ram_reg_20__44_ ( .D(n5392), .CLK(clk), .Q(ram[723]) );
  DFFPOSX1 ram_reg_20__45_ ( .D(n5391), .CLK(clk), .Q(ram[722]) );
  DFFPOSX1 ram_reg_20__46_ ( .D(n5390), .CLK(clk), .Q(ram[721]) );
  DFFPOSX1 ram_reg_20__47_ ( .D(n5389), .CLK(clk), .Q(ram[720]) );
  DFFPOSX1 ram_reg_20__48_ ( .D(n5388), .CLK(clk), .Q(ram[719]) );
  DFFPOSX1 ram_reg_20__49_ ( .D(n5387), .CLK(clk), .Q(ram[718]) );
  DFFPOSX1 ram_reg_20__50_ ( .D(n5386), .CLK(clk), .Q(ram[717]) );
  DFFPOSX1 ram_reg_20__51_ ( .D(n5385), .CLK(clk), .Q(ram[716]) );
  DFFPOSX1 ram_reg_20__52_ ( .D(n5384), .CLK(clk), .Q(ram[715]) );
  DFFPOSX1 ram_reg_20__53_ ( .D(n5383), .CLK(clk), .Q(ram[714]) );
  DFFPOSX1 ram_reg_20__54_ ( .D(n5382), .CLK(clk), .Q(ram[713]) );
  DFFPOSX1 ram_reg_20__55_ ( .D(n5381), .CLK(clk), .Q(ram[712]) );
  DFFPOSX1 ram_reg_20__56_ ( .D(n5380), .CLK(clk), .Q(ram[711]) );
  DFFPOSX1 ram_reg_20__57_ ( .D(n5379), .CLK(clk), .Q(ram[710]) );
  DFFPOSX1 ram_reg_20__58_ ( .D(n5378), .CLK(clk), .Q(ram[709]) );
  DFFPOSX1 ram_reg_20__59_ ( .D(n5377), .CLK(clk), .Q(ram[708]) );
  DFFPOSX1 ram_reg_20__60_ ( .D(n5376), .CLK(clk), .Q(ram[707]) );
  DFFPOSX1 ram_reg_20__61_ ( .D(n5375), .CLK(clk), .Q(ram[706]) );
  DFFPOSX1 ram_reg_20__62_ ( .D(n5374), .CLK(clk), .Q(ram[705]) );
  DFFPOSX1 ram_reg_20__63_ ( .D(n5373), .CLK(clk), .Q(ram[704]) );
  DFFPOSX1 ram_reg_21__0_ ( .D(n5372), .CLK(clk), .Q(ram[703]) );
  DFFPOSX1 ram_reg_21__1_ ( .D(n5371), .CLK(clk), .Q(ram[702]) );
  DFFPOSX1 ram_reg_21__2_ ( .D(n5370), .CLK(clk), .Q(ram[701]) );
  DFFPOSX1 ram_reg_21__3_ ( .D(n5369), .CLK(clk), .Q(ram[700]) );
  DFFPOSX1 ram_reg_21__4_ ( .D(n5368), .CLK(clk), .Q(ram[699]) );
  DFFPOSX1 ram_reg_21__5_ ( .D(n5367), .CLK(clk), .Q(ram[698]) );
  DFFPOSX1 ram_reg_21__6_ ( .D(n5366), .CLK(clk), .Q(ram[697]) );
  DFFPOSX1 ram_reg_21__7_ ( .D(n5365), .CLK(clk), .Q(ram[696]) );
  DFFPOSX1 ram_reg_21__8_ ( .D(n5364), .CLK(clk), .Q(ram[695]) );
  DFFPOSX1 ram_reg_21__9_ ( .D(n5363), .CLK(clk), .Q(ram[694]) );
  DFFPOSX1 ram_reg_21__10_ ( .D(n5362), .CLK(clk), .Q(ram[693]) );
  DFFPOSX1 ram_reg_21__11_ ( .D(n5361), .CLK(clk), .Q(ram[692]) );
  DFFPOSX1 ram_reg_21__12_ ( .D(n5360), .CLK(clk), .Q(ram[691]) );
  DFFPOSX1 ram_reg_21__13_ ( .D(n5359), .CLK(clk), .Q(ram[690]) );
  DFFPOSX1 ram_reg_21__14_ ( .D(n5358), .CLK(clk), .Q(ram[689]) );
  DFFPOSX1 ram_reg_21__15_ ( .D(n5357), .CLK(clk), .Q(ram[688]) );
  DFFPOSX1 ram_reg_21__16_ ( .D(n5356), .CLK(clk), .Q(ram[687]) );
  DFFPOSX1 ram_reg_21__17_ ( .D(n5355), .CLK(clk), .Q(ram[686]) );
  DFFPOSX1 ram_reg_21__18_ ( .D(n5354), .CLK(clk), .Q(ram[685]) );
  DFFPOSX1 ram_reg_21__19_ ( .D(n5353), .CLK(clk), .Q(ram[684]) );
  DFFPOSX1 ram_reg_21__20_ ( .D(n5352), .CLK(clk), .Q(ram[683]) );
  DFFPOSX1 ram_reg_21__21_ ( .D(n5351), .CLK(clk), .Q(ram[682]) );
  DFFPOSX1 ram_reg_21__22_ ( .D(n5350), .CLK(clk), .Q(ram[681]) );
  DFFPOSX1 ram_reg_21__23_ ( .D(n5349), .CLK(clk), .Q(ram[680]) );
  DFFPOSX1 ram_reg_21__24_ ( .D(n5348), .CLK(clk), .Q(ram[679]) );
  DFFPOSX1 ram_reg_21__25_ ( .D(n5347), .CLK(clk), .Q(ram[678]) );
  DFFPOSX1 ram_reg_21__26_ ( .D(n5346), .CLK(clk), .Q(ram[677]) );
  DFFPOSX1 ram_reg_21__27_ ( .D(n5345), .CLK(clk), .Q(ram[676]) );
  DFFPOSX1 ram_reg_21__28_ ( .D(n5344), .CLK(clk), .Q(ram[675]) );
  DFFPOSX1 ram_reg_21__29_ ( .D(n5343), .CLK(clk), .Q(ram[674]) );
  DFFPOSX1 ram_reg_21__30_ ( .D(n5342), .CLK(clk), .Q(ram[673]) );
  DFFPOSX1 ram_reg_21__31_ ( .D(n5341), .CLK(clk), .Q(ram[672]) );
  DFFPOSX1 ram_reg_21__32_ ( .D(n5340), .CLK(clk), .Q(ram[671]) );
  DFFPOSX1 ram_reg_21__33_ ( .D(n5339), .CLK(clk), .Q(ram[670]) );
  DFFPOSX1 ram_reg_21__34_ ( .D(n5338), .CLK(clk), .Q(ram[669]) );
  DFFPOSX1 ram_reg_21__35_ ( .D(n5337), .CLK(clk), .Q(ram[668]) );
  DFFPOSX1 ram_reg_21__36_ ( .D(n5336), .CLK(clk), .Q(ram[667]) );
  DFFPOSX1 ram_reg_21__37_ ( .D(n5335), .CLK(clk), .Q(ram[666]) );
  DFFPOSX1 ram_reg_21__38_ ( .D(n5334), .CLK(clk), .Q(ram[665]) );
  DFFPOSX1 ram_reg_21__39_ ( .D(n5333), .CLK(clk), .Q(ram[664]) );
  DFFPOSX1 ram_reg_21__40_ ( .D(n5332), .CLK(clk), .Q(ram[663]) );
  DFFPOSX1 ram_reg_21__41_ ( .D(n5331), .CLK(clk), .Q(ram[662]) );
  DFFPOSX1 ram_reg_21__42_ ( .D(n5330), .CLK(clk), .Q(ram[661]) );
  DFFPOSX1 ram_reg_21__43_ ( .D(n5329), .CLK(clk), .Q(ram[660]) );
  DFFPOSX1 ram_reg_21__44_ ( .D(n5328), .CLK(clk), .Q(ram[659]) );
  DFFPOSX1 ram_reg_21__45_ ( .D(n5327), .CLK(clk), .Q(ram[658]) );
  DFFPOSX1 ram_reg_21__46_ ( .D(n5326), .CLK(clk), .Q(ram[657]) );
  DFFPOSX1 ram_reg_21__47_ ( .D(n5325), .CLK(clk), .Q(ram[656]) );
  DFFPOSX1 ram_reg_21__48_ ( .D(n5324), .CLK(clk), .Q(ram[655]) );
  DFFPOSX1 ram_reg_21__49_ ( .D(n5323), .CLK(clk), .Q(ram[654]) );
  DFFPOSX1 ram_reg_21__50_ ( .D(n5322), .CLK(clk), .Q(ram[653]) );
  DFFPOSX1 ram_reg_21__51_ ( .D(n5321), .CLK(clk), .Q(ram[652]) );
  DFFPOSX1 ram_reg_21__52_ ( .D(n5320), .CLK(clk), .Q(ram[651]) );
  DFFPOSX1 ram_reg_21__53_ ( .D(n5319), .CLK(clk), .Q(ram[650]) );
  DFFPOSX1 ram_reg_21__54_ ( .D(n5318), .CLK(clk), .Q(ram[649]) );
  DFFPOSX1 ram_reg_21__55_ ( .D(n5317), .CLK(clk), .Q(ram[648]) );
  DFFPOSX1 ram_reg_21__56_ ( .D(n5316), .CLK(clk), .Q(ram[647]) );
  DFFPOSX1 ram_reg_21__57_ ( .D(n5315), .CLK(clk), .Q(ram[646]) );
  DFFPOSX1 ram_reg_21__58_ ( .D(n5314), .CLK(clk), .Q(ram[645]) );
  DFFPOSX1 ram_reg_21__59_ ( .D(n5313), .CLK(clk), .Q(ram[644]) );
  DFFPOSX1 ram_reg_21__60_ ( .D(n5312), .CLK(clk), .Q(ram[643]) );
  DFFPOSX1 ram_reg_21__61_ ( .D(n5311), .CLK(clk), .Q(ram[642]) );
  DFFPOSX1 ram_reg_21__62_ ( .D(n5310), .CLK(clk), .Q(ram[641]) );
  DFFPOSX1 ram_reg_21__63_ ( .D(n5309), .CLK(clk), .Q(ram[640]) );
  DFFPOSX1 ram_reg_22__0_ ( .D(n5308), .CLK(clk), .Q(ram[639]) );
  DFFPOSX1 ram_reg_22__1_ ( .D(n5307), .CLK(clk), .Q(ram[638]) );
  DFFPOSX1 ram_reg_22__2_ ( .D(n5306), .CLK(clk), .Q(ram[637]) );
  DFFPOSX1 ram_reg_22__3_ ( .D(n5305), .CLK(clk), .Q(ram[636]) );
  DFFPOSX1 ram_reg_22__4_ ( .D(n5304), .CLK(clk), .Q(ram[635]) );
  DFFPOSX1 ram_reg_22__5_ ( .D(n5303), .CLK(clk), .Q(ram[634]) );
  DFFPOSX1 ram_reg_22__6_ ( .D(n5302), .CLK(clk), .Q(ram[633]) );
  DFFPOSX1 ram_reg_22__7_ ( .D(n5301), .CLK(clk), .Q(ram[632]) );
  DFFPOSX1 ram_reg_22__8_ ( .D(n5300), .CLK(clk), .Q(ram[631]) );
  DFFPOSX1 ram_reg_22__9_ ( .D(n5299), .CLK(clk), .Q(ram[630]) );
  DFFPOSX1 ram_reg_22__10_ ( .D(n5298), .CLK(clk), .Q(ram[629]) );
  DFFPOSX1 ram_reg_22__11_ ( .D(n5297), .CLK(clk), .Q(ram[628]) );
  DFFPOSX1 ram_reg_22__12_ ( .D(n5296), .CLK(clk), .Q(ram[627]) );
  DFFPOSX1 ram_reg_22__13_ ( .D(n5295), .CLK(clk), .Q(ram[626]) );
  DFFPOSX1 ram_reg_22__14_ ( .D(n5294), .CLK(clk), .Q(ram[625]) );
  DFFPOSX1 ram_reg_22__15_ ( .D(n5293), .CLK(clk), .Q(ram[624]) );
  DFFPOSX1 ram_reg_22__16_ ( .D(n5292), .CLK(clk), .Q(ram[623]) );
  DFFPOSX1 ram_reg_22__17_ ( .D(n5291), .CLK(clk), .Q(ram[622]) );
  DFFPOSX1 ram_reg_22__18_ ( .D(n5290), .CLK(clk), .Q(ram[621]) );
  DFFPOSX1 ram_reg_22__19_ ( .D(n5289), .CLK(clk), .Q(ram[620]) );
  DFFPOSX1 ram_reg_22__20_ ( .D(n5288), .CLK(clk), .Q(ram[619]) );
  DFFPOSX1 ram_reg_22__21_ ( .D(n5287), .CLK(clk), .Q(ram[618]) );
  DFFPOSX1 ram_reg_22__22_ ( .D(n5286), .CLK(clk), .Q(ram[617]) );
  DFFPOSX1 ram_reg_22__23_ ( .D(n5285), .CLK(clk), .Q(ram[616]) );
  DFFPOSX1 ram_reg_22__24_ ( .D(n5284), .CLK(clk), .Q(ram[615]) );
  DFFPOSX1 ram_reg_22__25_ ( .D(n5283), .CLK(clk), .Q(ram[614]) );
  DFFPOSX1 ram_reg_22__26_ ( .D(n5282), .CLK(clk), .Q(ram[613]) );
  DFFPOSX1 ram_reg_22__27_ ( .D(n5281), .CLK(clk), .Q(ram[612]) );
  DFFPOSX1 ram_reg_22__28_ ( .D(n5280), .CLK(clk), .Q(ram[611]) );
  DFFPOSX1 ram_reg_22__29_ ( .D(n5279), .CLK(clk), .Q(ram[610]) );
  DFFPOSX1 ram_reg_22__30_ ( .D(n5278), .CLK(clk), .Q(ram[609]) );
  DFFPOSX1 ram_reg_22__31_ ( .D(n5277), .CLK(clk), .Q(ram[608]) );
  DFFPOSX1 ram_reg_22__32_ ( .D(n5276), .CLK(clk), .Q(ram[607]) );
  DFFPOSX1 ram_reg_22__33_ ( .D(n5275), .CLK(clk), .Q(ram[606]) );
  DFFPOSX1 ram_reg_22__34_ ( .D(n5274), .CLK(clk), .Q(ram[605]) );
  DFFPOSX1 ram_reg_22__35_ ( .D(n5273), .CLK(clk), .Q(ram[604]) );
  DFFPOSX1 ram_reg_22__36_ ( .D(n5272), .CLK(clk), .Q(ram[603]) );
  DFFPOSX1 ram_reg_22__37_ ( .D(n5271), .CLK(clk), .Q(ram[602]) );
  DFFPOSX1 ram_reg_22__38_ ( .D(n5270), .CLK(clk), .Q(ram[601]) );
  DFFPOSX1 ram_reg_22__39_ ( .D(n5269), .CLK(clk), .Q(ram[600]) );
  DFFPOSX1 ram_reg_22__40_ ( .D(n5268), .CLK(clk), .Q(ram[599]) );
  DFFPOSX1 ram_reg_22__41_ ( .D(n5267), .CLK(clk), .Q(ram[598]) );
  DFFPOSX1 ram_reg_22__42_ ( .D(n5266), .CLK(clk), .Q(ram[597]) );
  DFFPOSX1 ram_reg_22__43_ ( .D(n5265), .CLK(clk), .Q(ram[596]) );
  DFFPOSX1 ram_reg_22__44_ ( .D(n5264), .CLK(clk), .Q(ram[595]) );
  DFFPOSX1 ram_reg_22__45_ ( .D(n5263), .CLK(clk), .Q(ram[594]) );
  DFFPOSX1 ram_reg_22__46_ ( .D(n5262), .CLK(clk), .Q(ram[593]) );
  DFFPOSX1 ram_reg_22__47_ ( .D(n5261), .CLK(clk), .Q(ram[592]) );
  DFFPOSX1 ram_reg_22__48_ ( .D(n5260), .CLK(clk), .Q(ram[591]) );
  DFFPOSX1 ram_reg_22__49_ ( .D(n5259), .CLK(clk), .Q(ram[590]) );
  DFFPOSX1 ram_reg_22__50_ ( .D(n5258), .CLK(clk), .Q(ram[589]) );
  DFFPOSX1 ram_reg_22__51_ ( .D(n5257), .CLK(clk), .Q(ram[588]) );
  DFFPOSX1 ram_reg_22__52_ ( .D(n5256), .CLK(clk), .Q(ram[587]) );
  DFFPOSX1 ram_reg_22__53_ ( .D(n5255), .CLK(clk), .Q(ram[586]) );
  DFFPOSX1 ram_reg_22__54_ ( .D(n5254), .CLK(clk), .Q(ram[585]) );
  DFFPOSX1 ram_reg_22__55_ ( .D(n5253), .CLK(clk), .Q(ram[584]) );
  DFFPOSX1 ram_reg_22__56_ ( .D(n5252), .CLK(clk), .Q(ram[583]) );
  DFFPOSX1 ram_reg_22__57_ ( .D(n5251), .CLK(clk), .Q(ram[582]) );
  DFFPOSX1 ram_reg_22__58_ ( .D(n5250), .CLK(clk), .Q(ram[581]) );
  DFFPOSX1 ram_reg_22__59_ ( .D(n5249), .CLK(clk), .Q(ram[580]) );
  DFFPOSX1 ram_reg_22__60_ ( .D(n5248), .CLK(clk), .Q(ram[579]) );
  DFFPOSX1 ram_reg_22__61_ ( .D(n5247), .CLK(clk), .Q(ram[578]) );
  DFFPOSX1 ram_reg_22__62_ ( .D(n5246), .CLK(clk), .Q(ram[577]) );
  DFFPOSX1 ram_reg_22__63_ ( .D(n5245), .CLK(clk), .Q(ram[576]) );
  DFFPOSX1 ram_reg_23__0_ ( .D(n5244), .CLK(clk), .Q(ram[575]) );
  DFFPOSX1 ram_reg_23__1_ ( .D(n5243), .CLK(clk), .Q(ram[574]) );
  DFFPOSX1 ram_reg_23__2_ ( .D(n5242), .CLK(clk), .Q(ram[573]) );
  DFFPOSX1 ram_reg_23__3_ ( .D(n5241), .CLK(clk), .Q(ram[572]) );
  DFFPOSX1 ram_reg_23__4_ ( .D(n5240), .CLK(clk), .Q(ram[571]) );
  DFFPOSX1 ram_reg_23__5_ ( .D(n5239), .CLK(clk), .Q(ram[570]) );
  DFFPOSX1 ram_reg_23__6_ ( .D(n5238), .CLK(clk), .Q(ram[569]) );
  DFFPOSX1 ram_reg_23__7_ ( .D(n5237), .CLK(clk), .Q(ram[568]) );
  DFFPOSX1 ram_reg_23__8_ ( .D(n5236), .CLK(clk), .Q(ram[567]) );
  DFFPOSX1 ram_reg_23__9_ ( .D(n5235), .CLK(clk), .Q(ram[566]) );
  DFFPOSX1 ram_reg_23__10_ ( .D(n5234), .CLK(clk), .Q(ram[565]) );
  DFFPOSX1 ram_reg_23__11_ ( .D(n5233), .CLK(clk), .Q(ram[564]) );
  DFFPOSX1 ram_reg_23__12_ ( .D(n5232), .CLK(clk), .Q(ram[563]) );
  DFFPOSX1 ram_reg_23__13_ ( .D(n5231), .CLK(clk), .Q(ram[562]) );
  DFFPOSX1 ram_reg_23__14_ ( .D(n5230), .CLK(clk), .Q(ram[561]) );
  DFFPOSX1 ram_reg_23__15_ ( .D(n5229), .CLK(clk), .Q(ram[560]) );
  DFFPOSX1 ram_reg_23__16_ ( .D(n5228), .CLK(clk), .Q(ram[559]) );
  DFFPOSX1 ram_reg_23__17_ ( .D(n5227), .CLK(clk), .Q(ram[558]) );
  DFFPOSX1 ram_reg_23__18_ ( .D(n5226), .CLK(clk), .Q(ram[557]) );
  DFFPOSX1 ram_reg_23__19_ ( .D(n5225), .CLK(clk), .Q(ram[556]) );
  DFFPOSX1 ram_reg_23__20_ ( .D(n5224), .CLK(clk), .Q(ram[555]) );
  DFFPOSX1 ram_reg_23__21_ ( .D(n5223), .CLK(clk), .Q(ram[554]) );
  DFFPOSX1 ram_reg_23__22_ ( .D(n5222), .CLK(clk), .Q(ram[553]) );
  DFFPOSX1 ram_reg_23__23_ ( .D(n5221), .CLK(clk), .Q(ram[552]) );
  DFFPOSX1 ram_reg_23__24_ ( .D(n5220), .CLK(clk), .Q(ram[551]) );
  DFFPOSX1 ram_reg_23__25_ ( .D(n5219), .CLK(clk), .Q(ram[550]) );
  DFFPOSX1 ram_reg_23__26_ ( .D(n5218), .CLK(clk), .Q(ram[549]) );
  DFFPOSX1 ram_reg_23__27_ ( .D(n5217), .CLK(clk), .Q(ram[548]) );
  DFFPOSX1 ram_reg_23__28_ ( .D(n5216), .CLK(clk), .Q(ram[547]) );
  DFFPOSX1 ram_reg_23__29_ ( .D(n5215), .CLK(clk), .Q(ram[546]) );
  DFFPOSX1 ram_reg_23__30_ ( .D(n5214), .CLK(clk), .Q(ram[545]) );
  DFFPOSX1 ram_reg_23__31_ ( .D(n5213), .CLK(clk), .Q(ram[544]) );
  DFFPOSX1 ram_reg_23__32_ ( .D(n5212), .CLK(clk), .Q(ram[543]) );
  DFFPOSX1 ram_reg_23__33_ ( .D(n5211), .CLK(clk), .Q(ram[542]) );
  DFFPOSX1 ram_reg_23__34_ ( .D(n5210), .CLK(clk), .Q(ram[541]) );
  DFFPOSX1 ram_reg_23__35_ ( .D(n5209), .CLK(clk), .Q(ram[540]) );
  DFFPOSX1 ram_reg_23__36_ ( .D(n5208), .CLK(clk), .Q(ram[539]) );
  DFFPOSX1 ram_reg_23__37_ ( .D(n5207), .CLK(clk), .Q(ram[538]) );
  DFFPOSX1 ram_reg_23__38_ ( .D(n5206), .CLK(clk), .Q(ram[537]) );
  DFFPOSX1 ram_reg_23__39_ ( .D(n5205), .CLK(clk), .Q(ram[536]) );
  DFFPOSX1 ram_reg_23__40_ ( .D(n5204), .CLK(clk), .Q(ram[535]) );
  DFFPOSX1 ram_reg_23__41_ ( .D(n5203), .CLK(clk), .Q(ram[534]) );
  DFFPOSX1 ram_reg_23__42_ ( .D(n5202), .CLK(clk), .Q(ram[533]) );
  DFFPOSX1 ram_reg_23__43_ ( .D(n5201), .CLK(clk), .Q(ram[532]) );
  DFFPOSX1 ram_reg_23__44_ ( .D(n5200), .CLK(clk), .Q(ram[531]) );
  DFFPOSX1 ram_reg_23__45_ ( .D(n5199), .CLK(clk), .Q(ram[530]) );
  DFFPOSX1 ram_reg_23__46_ ( .D(n5198), .CLK(clk), .Q(ram[529]) );
  DFFPOSX1 ram_reg_23__47_ ( .D(n5197), .CLK(clk), .Q(ram[528]) );
  DFFPOSX1 ram_reg_23__48_ ( .D(n5196), .CLK(clk), .Q(ram[527]) );
  DFFPOSX1 ram_reg_23__49_ ( .D(n5195), .CLK(clk), .Q(ram[526]) );
  DFFPOSX1 ram_reg_23__50_ ( .D(n5194), .CLK(clk), .Q(ram[525]) );
  DFFPOSX1 ram_reg_23__51_ ( .D(n5193), .CLK(clk), .Q(ram[524]) );
  DFFPOSX1 ram_reg_23__52_ ( .D(n5192), .CLK(clk), .Q(ram[523]) );
  DFFPOSX1 ram_reg_23__53_ ( .D(n5191), .CLK(clk), .Q(ram[522]) );
  DFFPOSX1 ram_reg_23__54_ ( .D(n5190), .CLK(clk), .Q(ram[521]) );
  DFFPOSX1 ram_reg_23__55_ ( .D(n5189), .CLK(clk), .Q(ram[520]) );
  DFFPOSX1 ram_reg_23__56_ ( .D(n5188), .CLK(clk), .Q(ram[519]) );
  DFFPOSX1 ram_reg_23__57_ ( .D(n5187), .CLK(clk), .Q(ram[518]) );
  DFFPOSX1 ram_reg_23__58_ ( .D(n5186), .CLK(clk), .Q(ram[517]) );
  DFFPOSX1 ram_reg_23__59_ ( .D(n5185), .CLK(clk), .Q(ram[516]) );
  DFFPOSX1 ram_reg_23__60_ ( .D(n5184), .CLK(clk), .Q(ram[515]) );
  DFFPOSX1 ram_reg_23__61_ ( .D(n5183), .CLK(clk), .Q(ram[514]) );
  DFFPOSX1 ram_reg_23__62_ ( .D(n5182), .CLK(clk), .Q(ram[513]) );
  DFFPOSX1 ram_reg_23__63_ ( .D(n5181), .CLK(clk), .Q(ram[512]) );
  DFFPOSX1 ram_reg_24__0_ ( .D(n5180), .CLK(clk), .Q(ram[511]) );
  DFFPOSX1 ram_reg_24__1_ ( .D(n5179), .CLK(clk), .Q(ram[510]) );
  DFFPOSX1 ram_reg_24__2_ ( .D(n5178), .CLK(clk), .Q(ram[509]) );
  DFFPOSX1 ram_reg_24__3_ ( .D(n5177), .CLK(clk), .Q(ram[508]) );
  DFFPOSX1 ram_reg_24__4_ ( .D(n5176), .CLK(clk), .Q(ram[507]) );
  DFFPOSX1 ram_reg_24__5_ ( .D(n5175), .CLK(clk), .Q(ram[506]) );
  DFFPOSX1 ram_reg_24__6_ ( .D(n5174), .CLK(clk), .Q(ram[505]) );
  DFFPOSX1 ram_reg_24__7_ ( .D(n5173), .CLK(clk), .Q(ram[504]) );
  DFFPOSX1 ram_reg_24__8_ ( .D(n5172), .CLK(clk), .Q(ram[503]) );
  DFFPOSX1 ram_reg_24__9_ ( .D(n5171), .CLK(clk), .Q(ram[502]) );
  DFFPOSX1 ram_reg_24__10_ ( .D(n5170), .CLK(clk), .Q(ram[501]) );
  DFFPOSX1 ram_reg_24__11_ ( .D(n5169), .CLK(clk), .Q(ram[500]) );
  DFFPOSX1 ram_reg_24__12_ ( .D(n5168), .CLK(clk), .Q(ram[499]) );
  DFFPOSX1 ram_reg_24__13_ ( .D(n5167), .CLK(clk), .Q(ram[498]) );
  DFFPOSX1 ram_reg_24__14_ ( .D(n5166), .CLK(clk), .Q(ram[497]) );
  DFFPOSX1 ram_reg_24__15_ ( .D(n5165), .CLK(clk), .Q(ram[496]) );
  DFFPOSX1 ram_reg_24__16_ ( .D(n5164), .CLK(clk), .Q(ram[495]) );
  DFFPOSX1 ram_reg_24__17_ ( .D(n5163), .CLK(clk), .Q(ram[494]) );
  DFFPOSX1 ram_reg_24__18_ ( .D(n5162), .CLK(clk), .Q(ram[493]) );
  DFFPOSX1 ram_reg_24__19_ ( .D(n5161), .CLK(clk), .Q(ram[492]) );
  DFFPOSX1 ram_reg_24__20_ ( .D(n5160), .CLK(clk), .Q(ram[491]) );
  DFFPOSX1 ram_reg_24__21_ ( .D(n5159), .CLK(clk), .Q(ram[490]) );
  DFFPOSX1 ram_reg_24__22_ ( .D(n5158), .CLK(clk), .Q(ram[489]) );
  DFFPOSX1 ram_reg_24__23_ ( .D(n5157), .CLK(clk), .Q(ram[488]) );
  DFFPOSX1 ram_reg_24__24_ ( .D(n5156), .CLK(clk), .Q(ram[487]) );
  DFFPOSX1 ram_reg_24__25_ ( .D(n5155), .CLK(clk), .Q(ram[486]) );
  DFFPOSX1 ram_reg_24__26_ ( .D(n5154), .CLK(clk), .Q(ram[485]) );
  DFFPOSX1 ram_reg_24__27_ ( .D(n5153), .CLK(clk), .Q(ram[484]) );
  DFFPOSX1 ram_reg_24__28_ ( .D(n5152), .CLK(clk), .Q(ram[483]) );
  DFFPOSX1 ram_reg_24__29_ ( .D(n5151), .CLK(clk), .Q(ram[482]) );
  DFFPOSX1 ram_reg_24__30_ ( .D(n5150), .CLK(clk), .Q(ram[481]) );
  DFFPOSX1 ram_reg_24__31_ ( .D(n5149), .CLK(clk), .Q(ram[480]) );
  DFFPOSX1 ram_reg_24__32_ ( .D(n5148), .CLK(clk), .Q(ram[479]) );
  DFFPOSX1 ram_reg_24__33_ ( .D(n5147), .CLK(clk), .Q(ram[478]) );
  DFFPOSX1 ram_reg_24__34_ ( .D(n5146), .CLK(clk), .Q(ram[477]) );
  DFFPOSX1 ram_reg_24__35_ ( .D(n5145), .CLK(clk), .Q(ram[476]) );
  DFFPOSX1 ram_reg_24__36_ ( .D(n5144), .CLK(clk), .Q(ram[475]) );
  DFFPOSX1 ram_reg_24__37_ ( .D(n5143), .CLK(clk), .Q(ram[474]) );
  DFFPOSX1 ram_reg_24__38_ ( .D(n5142), .CLK(clk), .Q(ram[473]) );
  DFFPOSX1 ram_reg_24__39_ ( .D(n5141), .CLK(clk), .Q(ram[472]) );
  DFFPOSX1 ram_reg_24__40_ ( .D(n5140), .CLK(clk), .Q(ram[471]) );
  DFFPOSX1 ram_reg_24__41_ ( .D(n5139), .CLK(clk), .Q(ram[470]) );
  DFFPOSX1 ram_reg_24__42_ ( .D(n5138), .CLK(clk), .Q(ram[469]) );
  DFFPOSX1 ram_reg_24__43_ ( .D(n5137), .CLK(clk), .Q(ram[468]) );
  DFFPOSX1 ram_reg_24__44_ ( .D(n5136), .CLK(clk), .Q(ram[467]) );
  DFFPOSX1 ram_reg_24__45_ ( .D(n5135), .CLK(clk), .Q(ram[466]) );
  DFFPOSX1 ram_reg_24__46_ ( .D(n5134), .CLK(clk), .Q(ram[465]) );
  DFFPOSX1 ram_reg_24__47_ ( .D(n5133), .CLK(clk), .Q(ram[464]) );
  DFFPOSX1 ram_reg_24__48_ ( .D(n5132), .CLK(clk), .Q(ram[463]) );
  DFFPOSX1 ram_reg_24__49_ ( .D(n5131), .CLK(clk), .Q(ram[462]) );
  DFFPOSX1 ram_reg_24__50_ ( .D(n5130), .CLK(clk), .Q(ram[461]) );
  DFFPOSX1 ram_reg_24__51_ ( .D(n5129), .CLK(clk), .Q(ram[460]) );
  DFFPOSX1 ram_reg_24__52_ ( .D(n5128), .CLK(clk), .Q(ram[459]) );
  DFFPOSX1 ram_reg_24__53_ ( .D(n5127), .CLK(clk), .Q(ram[458]) );
  DFFPOSX1 ram_reg_24__54_ ( .D(n5126), .CLK(clk), .Q(ram[457]) );
  DFFPOSX1 ram_reg_24__55_ ( .D(n5125), .CLK(clk), .Q(ram[456]) );
  DFFPOSX1 ram_reg_24__56_ ( .D(n5124), .CLK(clk), .Q(ram[455]) );
  DFFPOSX1 ram_reg_24__57_ ( .D(n5123), .CLK(clk), .Q(ram[454]) );
  DFFPOSX1 ram_reg_24__58_ ( .D(n5122), .CLK(clk), .Q(ram[453]) );
  DFFPOSX1 ram_reg_24__59_ ( .D(n5121), .CLK(clk), .Q(ram[452]) );
  DFFPOSX1 ram_reg_24__60_ ( .D(n5120), .CLK(clk), .Q(ram[451]) );
  DFFPOSX1 ram_reg_24__61_ ( .D(n5119), .CLK(clk), .Q(ram[450]) );
  DFFPOSX1 ram_reg_24__62_ ( .D(n5118), .CLK(clk), .Q(ram[449]) );
  DFFPOSX1 ram_reg_24__63_ ( .D(n5117), .CLK(clk), .Q(ram[448]) );
  DFFPOSX1 ram_reg_25__0_ ( .D(n5116), .CLK(clk), .Q(ram[447]) );
  DFFPOSX1 ram_reg_25__1_ ( .D(n5115), .CLK(clk), .Q(ram[446]) );
  DFFPOSX1 ram_reg_25__2_ ( .D(n5114), .CLK(clk), .Q(ram[445]) );
  DFFPOSX1 ram_reg_25__3_ ( .D(n5113), .CLK(clk), .Q(ram[444]) );
  DFFPOSX1 ram_reg_25__4_ ( .D(n5112), .CLK(clk), .Q(ram[443]) );
  DFFPOSX1 ram_reg_25__5_ ( .D(n5111), .CLK(clk), .Q(ram[442]) );
  DFFPOSX1 ram_reg_25__6_ ( .D(n5110), .CLK(clk), .Q(ram[441]) );
  DFFPOSX1 ram_reg_25__7_ ( .D(n5109), .CLK(clk), .Q(ram[440]) );
  DFFPOSX1 ram_reg_25__8_ ( .D(n5108), .CLK(clk), .Q(ram[439]) );
  DFFPOSX1 ram_reg_25__9_ ( .D(n5107), .CLK(clk), .Q(ram[438]) );
  DFFPOSX1 ram_reg_25__10_ ( .D(n5106), .CLK(clk), .Q(ram[437]) );
  DFFPOSX1 ram_reg_25__11_ ( .D(n5105), .CLK(clk), .Q(ram[436]) );
  DFFPOSX1 ram_reg_25__12_ ( .D(n5104), .CLK(clk), .Q(ram[435]) );
  DFFPOSX1 ram_reg_25__13_ ( .D(n5103), .CLK(clk), .Q(ram[434]) );
  DFFPOSX1 ram_reg_25__14_ ( .D(n5102), .CLK(clk), .Q(ram[433]) );
  DFFPOSX1 ram_reg_25__15_ ( .D(n5101), .CLK(clk), .Q(ram[432]) );
  DFFPOSX1 ram_reg_25__16_ ( .D(n5100), .CLK(clk), .Q(ram[431]) );
  DFFPOSX1 ram_reg_25__17_ ( .D(n5099), .CLK(clk), .Q(ram[430]) );
  DFFPOSX1 ram_reg_25__18_ ( .D(n5098), .CLK(clk), .Q(ram[429]) );
  DFFPOSX1 ram_reg_25__19_ ( .D(n5097), .CLK(clk), .Q(ram[428]) );
  DFFPOSX1 ram_reg_25__20_ ( .D(n5096), .CLK(clk), .Q(ram[427]) );
  DFFPOSX1 ram_reg_25__21_ ( .D(n5095), .CLK(clk), .Q(ram[426]) );
  DFFPOSX1 ram_reg_25__22_ ( .D(n5094), .CLK(clk), .Q(ram[425]) );
  DFFPOSX1 ram_reg_25__23_ ( .D(n5093), .CLK(clk), .Q(ram[424]) );
  DFFPOSX1 ram_reg_25__24_ ( .D(n5092), .CLK(clk), .Q(ram[423]) );
  DFFPOSX1 ram_reg_25__25_ ( .D(n5091), .CLK(clk), .Q(ram[422]) );
  DFFPOSX1 ram_reg_25__26_ ( .D(n5090), .CLK(clk), .Q(ram[421]) );
  DFFPOSX1 ram_reg_25__27_ ( .D(n5089), .CLK(clk), .Q(ram[420]) );
  DFFPOSX1 ram_reg_25__28_ ( .D(n5088), .CLK(clk), .Q(ram[419]) );
  DFFPOSX1 ram_reg_25__29_ ( .D(n5087), .CLK(clk), .Q(ram[418]) );
  DFFPOSX1 ram_reg_25__30_ ( .D(n5086), .CLK(clk), .Q(ram[417]) );
  DFFPOSX1 ram_reg_25__31_ ( .D(n5085), .CLK(clk), .Q(ram[416]) );
  DFFPOSX1 ram_reg_25__32_ ( .D(n5084), .CLK(clk), .Q(ram[415]) );
  DFFPOSX1 ram_reg_25__33_ ( .D(n5083), .CLK(clk), .Q(ram[414]) );
  DFFPOSX1 ram_reg_25__34_ ( .D(n5082), .CLK(clk), .Q(ram[413]) );
  DFFPOSX1 ram_reg_25__35_ ( .D(n5081), .CLK(clk), .Q(ram[412]) );
  DFFPOSX1 ram_reg_25__36_ ( .D(n5080), .CLK(clk), .Q(ram[411]) );
  DFFPOSX1 ram_reg_25__37_ ( .D(n5079), .CLK(clk), .Q(ram[410]) );
  DFFPOSX1 ram_reg_25__38_ ( .D(n5078), .CLK(clk), .Q(ram[409]) );
  DFFPOSX1 ram_reg_25__39_ ( .D(n5077), .CLK(clk), .Q(ram[408]) );
  DFFPOSX1 ram_reg_25__40_ ( .D(n5076), .CLK(clk), .Q(ram[407]) );
  DFFPOSX1 ram_reg_25__41_ ( .D(n5075), .CLK(clk), .Q(ram[406]) );
  DFFPOSX1 ram_reg_25__42_ ( .D(n5074), .CLK(clk), .Q(ram[405]) );
  DFFPOSX1 ram_reg_25__43_ ( .D(n5073), .CLK(clk), .Q(ram[404]) );
  DFFPOSX1 ram_reg_25__44_ ( .D(n5072), .CLK(clk), .Q(ram[403]) );
  DFFPOSX1 ram_reg_25__45_ ( .D(n5071), .CLK(clk), .Q(ram[402]) );
  DFFPOSX1 ram_reg_25__46_ ( .D(n5070), .CLK(clk), .Q(ram[401]) );
  DFFPOSX1 ram_reg_25__47_ ( .D(n5069), .CLK(clk), .Q(ram[400]) );
  DFFPOSX1 ram_reg_25__48_ ( .D(n5068), .CLK(clk), .Q(ram[399]) );
  DFFPOSX1 ram_reg_25__49_ ( .D(n5067), .CLK(clk), .Q(ram[398]) );
  DFFPOSX1 ram_reg_25__50_ ( .D(n5066), .CLK(clk), .Q(ram[397]) );
  DFFPOSX1 ram_reg_25__51_ ( .D(n5065), .CLK(clk), .Q(ram[396]) );
  DFFPOSX1 ram_reg_25__52_ ( .D(n5064), .CLK(clk), .Q(ram[395]) );
  DFFPOSX1 ram_reg_25__53_ ( .D(n5063), .CLK(clk), .Q(ram[394]) );
  DFFPOSX1 ram_reg_25__54_ ( .D(n5062), .CLK(clk), .Q(ram[393]) );
  DFFPOSX1 ram_reg_25__55_ ( .D(n5061), .CLK(clk), .Q(ram[392]) );
  DFFPOSX1 ram_reg_25__56_ ( .D(n5060), .CLK(clk), .Q(ram[391]) );
  DFFPOSX1 ram_reg_25__57_ ( .D(n5059), .CLK(clk), .Q(ram[390]) );
  DFFPOSX1 ram_reg_25__58_ ( .D(n5058), .CLK(clk), .Q(ram[389]) );
  DFFPOSX1 ram_reg_25__59_ ( .D(n5057), .CLK(clk), .Q(ram[388]) );
  DFFPOSX1 ram_reg_25__60_ ( .D(n5056), .CLK(clk), .Q(ram[387]) );
  DFFPOSX1 ram_reg_25__61_ ( .D(n5055), .CLK(clk), .Q(ram[386]) );
  DFFPOSX1 ram_reg_25__62_ ( .D(n5054), .CLK(clk), .Q(ram[385]) );
  DFFPOSX1 ram_reg_25__63_ ( .D(n5053), .CLK(clk), .Q(ram[384]) );
  DFFPOSX1 ram_reg_26__0_ ( .D(n5052), .CLK(clk), .Q(ram[383]) );
  DFFPOSX1 ram_reg_26__1_ ( .D(n5051), .CLK(clk), .Q(ram[382]) );
  DFFPOSX1 ram_reg_26__2_ ( .D(n5050), .CLK(clk), .Q(ram[381]) );
  DFFPOSX1 ram_reg_26__3_ ( .D(n5049), .CLK(clk), .Q(ram[380]) );
  DFFPOSX1 ram_reg_26__4_ ( .D(n5048), .CLK(clk), .Q(ram[379]) );
  DFFPOSX1 ram_reg_26__5_ ( .D(n5047), .CLK(clk), .Q(ram[378]) );
  DFFPOSX1 ram_reg_26__6_ ( .D(n5046), .CLK(clk), .Q(ram[377]) );
  DFFPOSX1 ram_reg_26__7_ ( .D(n5045), .CLK(clk), .Q(ram[376]) );
  DFFPOSX1 ram_reg_26__8_ ( .D(n5044), .CLK(clk), .Q(ram[375]) );
  DFFPOSX1 ram_reg_26__9_ ( .D(n5043), .CLK(clk), .Q(ram[374]) );
  DFFPOSX1 ram_reg_26__10_ ( .D(n5042), .CLK(clk), .Q(ram[373]) );
  DFFPOSX1 ram_reg_26__11_ ( .D(n5041), .CLK(clk), .Q(ram[372]) );
  DFFPOSX1 ram_reg_26__12_ ( .D(n5040), .CLK(clk), .Q(ram[371]) );
  DFFPOSX1 ram_reg_26__13_ ( .D(n5039), .CLK(clk), .Q(ram[370]) );
  DFFPOSX1 ram_reg_26__14_ ( .D(n5038), .CLK(clk), .Q(ram[369]) );
  DFFPOSX1 ram_reg_26__15_ ( .D(n5037), .CLK(clk), .Q(ram[368]) );
  DFFPOSX1 ram_reg_26__16_ ( .D(n5036), .CLK(clk), .Q(ram[367]) );
  DFFPOSX1 ram_reg_26__17_ ( .D(n5035), .CLK(clk), .Q(ram[366]) );
  DFFPOSX1 ram_reg_26__18_ ( .D(n5034), .CLK(clk), .Q(ram[365]) );
  DFFPOSX1 ram_reg_26__19_ ( .D(n5033), .CLK(clk), .Q(ram[364]) );
  DFFPOSX1 ram_reg_26__20_ ( .D(n5032), .CLK(clk), .Q(ram[363]) );
  DFFPOSX1 ram_reg_26__21_ ( .D(n5031), .CLK(clk), .Q(ram[362]) );
  DFFPOSX1 ram_reg_26__22_ ( .D(n5030), .CLK(clk), .Q(ram[361]) );
  DFFPOSX1 ram_reg_26__23_ ( .D(n5029), .CLK(clk), .Q(ram[360]) );
  DFFPOSX1 ram_reg_26__24_ ( .D(n5028), .CLK(clk), .Q(ram[359]) );
  DFFPOSX1 ram_reg_26__25_ ( .D(n5027), .CLK(clk), .Q(ram[358]) );
  DFFPOSX1 ram_reg_26__26_ ( .D(n5026), .CLK(clk), .Q(ram[357]) );
  DFFPOSX1 ram_reg_26__27_ ( .D(n5025), .CLK(clk), .Q(ram[356]) );
  DFFPOSX1 ram_reg_26__28_ ( .D(n5024), .CLK(clk), .Q(ram[355]) );
  DFFPOSX1 ram_reg_26__29_ ( .D(n5023), .CLK(clk), .Q(ram[354]) );
  DFFPOSX1 ram_reg_26__30_ ( .D(n5022), .CLK(clk), .Q(ram[353]) );
  DFFPOSX1 ram_reg_26__31_ ( .D(n5021), .CLK(clk), .Q(ram[352]) );
  DFFPOSX1 ram_reg_26__32_ ( .D(n5020), .CLK(clk), .Q(ram[351]) );
  DFFPOSX1 ram_reg_26__33_ ( .D(n5019), .CLK(clk), .Q(ram[350]) );
  DFFPOSX1 ram_reg_26__34_ ( .D(n5018), .CLK(clk), .Q(ram[349]) );
  DFFPOSX1 ram_reg_26__35_ ( .D(n5017), .CLK(clk), .Q(ram[348]) );
  DFFPOSX1 ram_reg_26__36_ ( .D(n5016), .CLK(clk), .Q(ram[347]) );
  DFFPOSX1 ram_reg_26__37_ ( .D(n5015), .CLK(clk), .Q(ram[346]) );
  DFFPOSX1 ram_reg_26__38_ ( .D(n5014), .CLK(clk), .Q(ram[345]) );
  DFFPOSX1 ram_reg_26__39_ ( .D(n5013), .CLK(clk), .Q(ram[344]) );
  DFFPOSX1 ram_reg_26__40_ ( .D(n5012), .CLK(clk), .Q(ram[343]) );
  DFFPOSX1 ram_reg_26__41_ ( .D(n5011), .CLK(clk), .Q(ram[342]) );
  DFFPOSX1 ram_reg_26__42_ ( .D(n5010), .CLK(clk), .Q(ram[341]) );
  DFFPOSX1 ram_reg_26__43_ ( .D(n5009), .CLK(clk), .Q(ram[340]) );
  DFFPOSX1 ram_reg_26__44_ ( .D(n5008), .CLK(clk), .Q(ram[339]) );
  DFFPOSX1 ram_reg_26__45_ ( .D(n5007), .CLK(clk), .Q(ram[338]) );
  DFFPOSX1 ram_reg_26__46_ ( .D(n5006), .CLK(clk), .Q(ram[337]) );
  DFFPOSX1 ram_reg_26__47_ ( .D(n5005), .CLK(clk), .Q(ram[336]) );
  DFFPOSX1 ram_reg_26__48_ ( .D(n5004), .CLK(clk), .Q(ram[335]) );
  DFFPOSX1 ram_reg_26__49_ ( .D(n5003), .CLK(clk), .Q(ram[334]) );
  DFFPOSX1 ram_reg_26__50_ ( .D(n5002), .CLK(clk), .Q(ram[333]) );
  DFFPOSX1 ram_reg_26__51_ ( .D(n5001), .CLK(clk), .Q(ram[332]) );
  DFFPOSX1 ram_reg_26__52_ ( .D(n5000), .CLK(clk), .Q(ram[331]) );
  DFFPOSX1 ram_reg_26__53_ ( .D(n4999), .CLK(clk), .Q(ram[330]) );
  DFFPOSX1 ram_reg_26__54_ ( .D(n4998), .CLK(clk), .Q(ram[329]) );
  DFFPOSX1 ram_reg_26__55_ ( .D(n4997), .CLK(clk), .Q(ram[328]) );
  DFFPOSX1 ram_reg_26__56_ ( .D(n4996), .CLK(clk), .Q(ram[327]) );
  DFFPOSX1 ram_reg_26__57_ ( .D(n4995), .CLK(clk), .Q(ram[326]) );
  DFFPOSX1 ram_reg_26__58_ ( .D(n4994), .CLK(clk), .Q(ram[325]) );
  DFFPOSX1 ram_reg_26__59_ ( .D(n4993), .CLK(clk), .Q(ram[324]) );
  DFFPOSX1 ram_reg_26__60_ ( .D(n4992), .CLK(clk), .Q(ram[323]) );
  DFFPOSX1 ram_reg_26__61_ ( .D(n4991), .CLK(clk), .Q(ram[322]) );
  DFFPOSX1 ram_reg_26__62_ ( .D(n4990), .CLK(clk), .Q(ram[321]) );
  DFFPOSX1 ram_reg_26__63_ ( .D(n4989), .CLK(clk), .Q(ram[320]) );
  DFFPOSX1 ram_reg_27__0_ ( .D(n4988), .CLK(clk), .Q(ram[319]) );
  DFFPOSX1 ram_reg_27__1_ ( .D(n4987), .CLK(clk), .Q(ram[318]) );
  DFFPOSX1 ram_reg_27__2_ ( .D(n4986), .CLK(clk), .Q(ram[317]) );
  DFFPOSX1 ram_reg_27__3_ ( .D(n4985), .CLK(clk), .Q(ram[316]) );
  DFFPOSX1 ram_reg_27__4_ ( .D(n4984), .CLK(clk), .Q(ram[315]) );
  DFFPOSX1 ram_reg_27__5_ ( .D(n4983), .CLK(clk), .Q(ram[314]) );
  DFFPOSX1 ram_reg_27__6_ ( .D(n4982), .CLK(clk), .Q(ram[313]) );
  DFFPOSX1 ram_reg_27__7_ ( .D(n4981), .CLK(clk), .Q(ram[312]) );
  DFFPOSX1 ram_reg_27__8_ ( .D(n4980), .CLK(clk), .Q(ram[311]) );
  DFFPOSX1 ram_reg_27__9_ ( .D(n4979), .CLK(clk), .Q(ram[310]) );
  DFFPOSX1 ram_reg_27__10_ ( .D(n4978), .CLK(clk), .Q(ram[309]) );
  DFFPOSX1 ram_reg_27__11_ ( .D(n4977), .CLK(clk), .Q(ram[308]) );
  DFFPOSX1 ram_reg_27__12_ ( .D(n4976), .CLK(clk), .Q(ram[307]) );
  DFFPOSX1 ram_reg_27__13_ ( .D(n4975), .CLK(clk), .Q(ram[306]) );
  DFFPOSX1 ram_reg_27__14_ ( .D(n4974), .CLK(clk), .Q(ram[305]) );
  DFFPOSX1 ram_reg_27__15_ ( .D(n4973), .CLK(clk), .Q(ram[304]) );
  DFFPOSX1 ram_reg_27__16_ ( .D(n4972), .CLK(clk), .Q(ram[303]) );
  DFFPOSX1 ram_reg_27__17_ ( .D(n4971), .CLK(clk), .Q(ram[302]) );
  DFFPOSX1 ram_reg_27__18_ ( .D(n4970), .CLK(clk), .Q(ram[301]) );
  DFFPOSX1 ram_reg_27__19_ ( .D(n4969), .CLK(clk), .Q(ram[300]) );
  DFFPOSX1 ram_reg_27__20_ ( .D(n4968), .CLK(clk), .Q(ram[299]) );
  DFFPOSX1 ram_reg_27__21_ ( .D(n4967), .CLK(clk), .Q(ram[298]) );
  DFFPOSX1 ram_reg_27__22_ ( .D(n4966), .CLK(clk), .Q(ram[297]) );
  DFFPOSX1 ram_reg_27__23_ ( .D(n4965), .CLK(clk), .Q(ram[296]) );
  DFFPOSX1 ram_reg_27__24_ ( .D(n4964), .CLK(clk), .Q(ram[295]) );
  DFFPOSX1 ram_reg_27__25_ ( .D(n4963), .CLK(clk), .Q(ram[294]) );
  DFFPOSX1 ram_reg_27__26_ ( .D(n4962), .CLK(clk), .Q(ram[293]) );
  DFFPOSX1 ram_reg_27__27_ ( .D(n4961), .CLK(clk), .Q(ram[292]) );
  DFFPOSX1 ram_reg_27__28_ ( .D(n4960), .CLK(clk), .Q(ram[291]) );
  DFFPOSX1 ram_reg_27__29_ ( .D(n4959), .CLK(clk), .Q(ram[290]) );
  DFFPOSX1 ram_reg_27__30_ ( .D(n4958), .CLK(clk), .Q(ram[289]) );
  DFFPOSX1 ram_reg_27__31_ ( .D(n4957), .CLK(clk), .Q(ram[288]) );
  DFFPOSX1 ram_reg_27__32_ ( .D(n4956), .CLK(clk), .Q(ram[287]) );
  DFFPOSX1 ram_reg_27__33_ ( .D(n4955), .CLK(clk), .Q(ram[286]) );
  DFFPOSX1 ram_reg_27__34_ ( .D(n4954), .CLK(clk), .Q(ram[285]) );
  DFFPOSX1 ram_reg_27__35_ ( .D(n4953), .CLK(clk), .Q(ram[284]) );
  DFFPOSX1 ram_reg_27__36_ ( .D(n4952), .CLK(clk), .Q(ram[283]) );
  DFFPOSX1 ram_reg_27__37_ ( .D(n4951), .CLK(clk), .Q(ram[282]) );
  DFFPOSX1 ram_reg_27__38_ ( .D(n4950), .CLK(clk), .Q(ram[281]) );
  DFFPOSX1 ram_reg_27__39_ ( .D(n4949), .CLK(clk), .Q(ram[280]) );
  DFFPOSX1 ram_reg_27__40_ ( .D(n4948), .CLK(clk), .Q(ram[279]) );
  DFFPOSX1 ram_reg_27__41_ ( .D(n4947), .CLK(clk), .Q(ram[278]) );
  DFFPOSX1 ram_reg_27__42_ ( .D(n4946), .CLK(clk), .Q(ram[277]) );
  DFFPOSX1 ram_reg_27__43_ ( .D(n4945), .CLK(clk), .Q(ram[276]) );
  DFFPOSX1 ram_reg_27__44_ ( .D(n4944), .CLK(clk), .Q(ram[275]) );
  DFFPOSX1 ram_reg_27__45_ ( .D(n4943), .CLK(clk), .Q(ram[274]) );
  DFFPOSX1 ram_reg_27__46_ ( .D(n4942), .CLK(clk), .Q(ram[273]) );
  DFFPOSX1 ram_reg_27__47_ ( .D(n4941), .CLK(clk), .Q(ram[272]) );
  DFFPOSX1 ram_reg_27__48_ ( .D(n4940), .CLK(clk), .Q(ram[271]) );
  DFFPOSX1 ram_reg_27__49_ ( .D(n4939), .CLK(clk), .Q(ram[270]) );
  DFFPOSX1 ram_reg_27__50_ ( .D(n4938), .CLK(clk), .Q(ram[269]) );
  DFFPOSX1 ram_reg_27__51_ ( .D(n4937), .CLK(clk), .Q(ram[268]) );
  DFFPOSX1 ram_reg_27__52_ ( .D(n4936), .CLK(clk), .Q(ram[267]) );
  DFFPOSX1 ram_reg_27__53_ ( .D(n4935), .CLK(clk), .Q(ram[266]) );
  DFFPOSX1 ram_reg_27__54_ ( .D(n4934), .CLK(clk), .Q(ram[265]) );
  DFFPOSX1 ram_reg_27__55_ ( .D(n4933), .CLK(clk), .Q(ram[264]) );
  DFFPOSX1 ram_reg_27__56_ ( .D(n4932), .CLK(clk), .Q(ram[263]) );
  DFFPOSX1 ram_reg_27__57_ ( .D(n4931), .CLK(clk), .Q(ram[262]) );
  DFFPOSX1 ram_reg_27__58_ ( .D(n4930), .CLK(clk), .Q(ram[261]) );
  DFFPOSX1 ram_reg_27__59_ ( .D(n4929), .CLK(clk), .Q(ram[260]) );
  DFFPOSX1 ram_reg_27__60_ ( .D(n4928), .CLK(clk), .Q(ram[259]) );
  DFFPOSX1 ram_reg_27__61_ ( .D(n4927), .CLK(clk), .Q(ram[258]) );
  DFFPOSX1 ram_reg_27__62_ ( .D(n4926), .CLK(clk), .Q(ram[257]) );
  DFFPOSX1 ram_reg_27__63_ ( .D(n4925), .CLK(clk), .Q(ram[256]) );
  DFFPOSX1 ram_reg_28__0_ ( .D(n4924), .CLK(clk), .Q(ram[255]) );
  DFFPOSX1 ram_reg_28__1_ ( .D(n4923), .CLK(clk), .Q(ram[254]) );
  DFFPOSX1 ram_reg_28__2_ ( .D(n4922), .CLK(clk), .Q(ram[253]) );
  DFFPOSX1 ram_reg_28__3_ ( .D(n4921), .CLK(clk), .Q(ram[252]) );
  DFFPOSX1 ram_reg_28__4_ ( .D(n4920), .CLK(clk), .Q(ram[251]) );
  DFFPOSX1 ram_reg_28__5_ ( .D(n4919), .CLK(clk), .Q(ram[250]) );
  DFFPOSX1 ram_reg_28__6_ ( .D(n4918), .CLK(clk), .Q(ram[249]) );
  DFFPOSX1 ram_reg_28__7_ ( .D(n4917), .CLK(clk), .Q(ram[248]) );
  DFFPOSX1 ram_reg_28__8_ ( .D(n4916), .CLK(clk), .Q(ram[247]) );
  DFFPOSX1 ram_reg_28__9_ ( .D(n4915), .CLK(clk), .Q(ram[246]) );
  DFFPOSX1 ram_reg_28__10_ ( .D(n4914), .CLK(clk), .Q(ram[245]) );
  DFFPOSX1 ram_reg_28__11_ ( .D(n4913), .CLK(clk), .Q(ram[244]) );
  DFFPOSX1 ram_reg_28__12_ ( .D(n4912), .CLK(clk), .Q(ram[243]) );
  DFFPOSX1 ram_reg_28__13_ ( .D(n4911), .CLK(clk), .Q(ram[242]) );
  DFFPOSX1 ram_reg_28__14_ ( .D(n4910), .CLK(clk), .Q(ram[241]) );
  DFFPOSX1 ram_reg_28__15_ ( .D(n4909), .CLK(clk), .Q(ram[240]) );
  DFFPOSX1 ram_reg_28__16_ ( .D(n4908), .CLK(clk), .Q(ram[239]) );
  DFFPOSX1 ram_reg_28__17_ ( .D(n4907), .CLK(clk), .Q(ram[238]) );
  DFFPOSX1 ram_reg_28__18_ ( .D(n4906), .CLK(clk), .Q(ram[237]) );
  DFFPOSX1 ram_reg_28__19_ ( .D(n4905), .CLK(clk), .Q(ram[236]) );
  DFFPOSX1 ram_reg_28__20_ ( .D(n4904), .CLK(clk), .Q(ram[235]) );
  DFFPOSX1 ram_reg_28__21_ ( .D(n4903), .CLK(clk), .Q(ram[234]) );
  DFFPOSX1 ram_reg_28__22_ ( .D(n4902), .CLK(clk), .Q(ram[233]) );
  DFFPOSX1 ram_reg_28__23_ ( .D(n4901), .CLK(clk), .Q(ram[232]) );
  DFFPOSX1 ram_reg_28__24_ ( .D(n4900), .CLK(clk), .Q(ram[231]) );
  DFFPOSX1 ram_reg_28__25_ ( .D(n4899), .CLK(clk), .Q(ram[230]) );
  DFFPOSX1 ram_reg_28__26_ ( .D(n4898), .CLK(clk), .Q(ram[229]) );
  DFFPOSX1 ram_reg_28__27_ ( .D(n4897), .CLK(clk), .Q(ram[228]) );
  DFFPOSX1 ram_reg_28__28_ ( .D(n4896), .CLK(clk), .Q(ram[227]) );
  DFFPOSX1 ram_reg_28__29_ ( .D(n4895), .CLK(clk), .Q(ram[226]) );
  DFFPOSX1 ram_reg_28__30_ ( .D(n4894), .CLK(clk), .Q(ram[225]) );
  DFFPOSX1 ram_reg_28__31_ ( .D(n4893), .CLK(clk), .Q(ram[224]) );
  DFFPOSX1 ram_reg_28__32_ ( .D(n4892), .CLK(clk), .Q(ram[223]) );
  DFFPOSX1 ram_reg_28__33_ ( .D(n4891), .CLK(clk), .Q(ram[222]) );
  DFFPOSX1 ram_reg_28__34_ ( .D(n4890), .CLK(clk), .Q(ram[221]) );
  DFFPOSX1 ram_reg_28__35_ ( .D(n4889), .CLK(clk), .Q(ram[220]) );
  DFFPOSX1 ram_reg_28__36_ ( .D(n4888), .CLK(clk), .Q(ram[219]) );
  DFFPOSX1 ram_reg_28__37_ ( .D(n4887), .CLK(clk), .Q(ram[218]) );
  DFFPOSX1 ram_reg_28__38_ ( .D(n4886), .CLK(clk), .Q(ram[217]) );
  DFFPOSX1 ram_reg_28__39_ ( .D(n4885), .CLK(clk), .Q(ram[216]) );
  DFFPOSX1 ram_reg_28__40_ ( .D(n4884), .CLK(clk), .Q(ram[215]) );
  DFFPOSX1 ram_reg_28__41_ ( .D(n4883), .CLK(clk), .Q(ram[214]) );
  DFFPOSX1 ram_reg_28__42_ ( .D(n4882), .CLK(clk), .Q(ram[213]) );
  DFFPOSX1 ram_reg_28__43_ ( .D(n4881), .CLK(clk), .Q(ram[212]) );
  DFFPOSX1 ram_reg_28__44_ ( .D(n4880), .CLK(clk), .Q(ram[211]) );
  DFFPOSX1 ram_reg_28__45_ ( .D(n4879), .CLK(clk), .Q(ram[210]) );
  DFFPOSX1 ram_reg_28__46_ ( .D(n4878), .CLK(clk), .Q(ram[209]) );
  DFFPOSX1 ram_reg_28__47_ ( .D(n4877), .CLK(clk), .Q(ram[208]) );
  DFFPOSX1 ram_reg_28__48_ ( .D(n4876), .CLK(clk), .Q(ram[207]) );
  DFFPOSX1 ram_reg_28__49_ ( .D(n4875), .CLK(clk), .Q(ram[206]) );
  DFFPOSX1 ram_reg_28__50_ ( .D(n4874), .CLK(clk), .Q(ram[205]) );
  DFFPOSX1 ram_reg_28__51_ ( .D(n4873), .CLK(clk), .Q(ram[204]) );
  DFFPOSX1 ram_reg_28__52_ ( .D(n4872), .CLK(clk), .Q(ram[203]) );
  DFFPOSX1 ram_reg_28__53_ ( .D(n4871), .CLK(clk), .Q(ram[202]) );
  DFFPOSX1 ram_reg_28__54_ ( .D(n4870), .CLK(clk), .Q(ram[201]) );
  DFFPOSX1 ram_reg_28__55_ ( .D(n4869), .CLK(clk), .Q(ram[200]) );
  DFFPOSX1 ram_reg_28__56_ ( .D(n4868), .CLK(clk), .Q(ram[199]) );
  DFFPOSX1 ram_reg_28__57_ ( .D(n4867), .CLK(clk), .Q(ram[198]) );
  DFFPOSX1 ram_reg_28__58_ ( .D(n4866), .CLK(clk), .Q(ram[197]) );
  DFFPOSX1 ram_reg_28__59_ ( .D(n4865), .CLK(clk), .Q(ram[196]) );
  DFFPOSX1 ram_reg_28__60_ ( .D(n4864), .CLK(clk), .Q(ram[195]) );
  DFFPOSX1 ram_reg_28__61_ ( .D(n4863), .CLK(clk), .Q(ram[194]) );
  DFFPOSX1 ram_reg_28__62_ ( .D(n4862), .CLK(clk), .Q(ram[193]) );
  DFFPOSX1 ram_reg_28__63_ ( .D(n4861), .CLK(clk), .Q(ram[192]) );
  DFFPOSX1 ram_reg_29__0_ ( .D(n4860), .CLK(clk), .Q(ram[191]) );
  DFFPOSX1 ram_reg_29__1_ ( .D(n4859), .CLK(clk), .Q(ram[190]) );
  DFFPOSX1 ram_reg_29__2_ ( .D(n4858), .CLK(clk), .Q(ram[189]) );
  DFFPOSX1 ram_reg_29__3_ ( .D(n4857), .CLK(clk), .Q(ram[188]) );
  DFFPOSX1 ram_reg_29__4_ ( .D(n4856), .CLK(clk), .Q(ram[187]) );
  DFFPOSX1 ram_reg_29__5_ ( .D(n4855), .CLK(clk), .Q(ram[186]) );
  DFFPOSX1 ram_reg_29__6_ ( .D(n4854), .CLK(clk), .Q(ram[185]) );
  DFFPOSX1 ram_reg_29__7_ ( .D(n4853), .CLK(clk), .Q(ram[184]) );
  DFFPOSX1 ram_reg_29__8_ ( .D(n4852), .CLK(clk), .Q(ram[183]) );
  DFFPOSX1 ram_reg_29__9_ ( .D(n4851), .CLK(clk), .Q(ram[182]) );
  DFFPOSX1 ram_reg_29__10_ ( .D(n4850), .CLK(clk), .Q(ram[181]) );
  DFFPOSX1 ram_reg_29__11_ ( .D(n4849), .CLK(clk), .Q(ram[180]) );
  DFFPOSX1 ram_reg_29__12_ ( .D(n4848), .CLK(clk), .Q(ram[179]) );
  DFFPOSX1 ram_reg_29__13_ ( .D(n4847), .CLK(clk), .Q(ram[178]) );
  DFFPOSX1 ram_reg_29__14_ ( .D(n4846), .CLK(clk), .Q(ram[177]) );
  DFFPOSX1 ram_reg_29__15_ ( .D(n4845), .CLK(clk), .Q(ram[176]) );
  DFFPOSX1 ram_reg_29__16_ ( .D(n4844), .CLK(clk), .Q(ram[175]) );
  DFFPOSX1 ram_reg_29__17_ ( .D(n4843), .CLK(clk), .Q(ram[174]) );
  DFFPOSX1 ram_reg_29__18_ ( .D(n4842), .CLK(clk), .Q(ram[173]) );
  DFFPOSX1 ram_reg_29__19_ ( .D(n4841), .CLK(clk), .Q(ram[172]) );
  DFFPOSX1 ram_reg_29__20_ ( .D(n4840), .CLK(clk), .Q(ram[171]) );
  DFFPOSX1 ram_reg_29__21_ ( .D(n4839), .CLK(clk), .Q(ram[170]) );
  DFFPOSX1 ram_reg_29__22_ ( .D(n4838), .CLK(clk), .Q(ram[169]) );
  DFFPOSX1 ram_reg_29__23_ ( .D(n4837), .CLK(clk), .Q(ram[168]) );
  DFFPOSX1 ram_reg_29__24_ ( .D(n4836), .CLK(clk), .Q(ram[167]) );
  DFFPOSX1 ram_reg_29__25_ ( .D(n4835), .CLK(clk), .Q(ram[166]) );
  DFFPOSX1 ram_reg_29__26_ ( .D(n4834), .CLK(clk), .Q(ram[165]) );
  DFFPOSX1 ram_reg_29__27_ ( .D(n4833), .CLK(clk), .Q(ram[164]) );
  DFFPOSX1 ram_reg_29__28_ ( .D(n4832), .CLK(clk), .Q(ram[163]) );
  DFFPOSX1 ram_reg_29__29_ ( .D(n4831), .CLK(clk), .Q(ram[162]) );
  DFFPOSX1 ram_reg_29__30_ ( .D(n4830), .CLK(clk), .Q(ram[161]) );
  DFFPOSX1 ram_reg_29__31_ ( .D(n4829), .CLK(clk), .Q(ram[160]) );
  DFFPOSX1 ram_reg_29__32_ ( .D(n4828), .CLK(clk), .Q(ram[159]) );
  DFFPOSX1 ram_reg_29__33_ ( .D(n4827), .CLK(clk), .Q(ram[158]) );
  DFFPOSX1 ram_reg_29__34_ ( .D(n4826), .CLK(clk), .Q(ram[157]) );
  DFFPOSX1 ram_reg_29__35_ ( .D(n4825), .CLK(clk), .Q(ram[156]) );
  DFFPOSX1 ram_reg_29__36_ ( .D(n4824), .CLK(clk), .Q(ram[155]) );
  DFFPOSX1 ram_reg_29__37_ ( .D(n4823), .CLK(clk), .Q(ram[154]) );
  DFFPOSX1 ram_reg_29__38_ ( .D(n4822), .CLK(clk), .Q(ram[153]) );
  DFFPOSX1 ram_reg_29__39_ ( .D(n4821), .CLK(clk), .Q(ram[152]) );
  DFFPOSX1 ram_reg_29__40_ ( .D(n4820), .CLK(clk), .Q(ram[151]) );
  DFFPOSX1 ram_reg_29__41_ ( .D(n4819), .CLK(clk), .Q(ram[150]) );
  DFFPOSX1 ram_reg_29__42_ ( .D(n4818), .CLK(clk), .Q(ram[149]) );
  DFFPOSX1 ram_reg_29__43_ ( .D(n4817), .CLK(clk), .Q(ram[148]) );
  DFFPOSX1 ram_reg_29__44_ ( .D(n4816), .CLK(clk), .Q(ram[147]) );
  DFFPOSX1 ram_reg_29__45_ ( .D(n4815), .CLK(clk), .Q(ram[146]) );
  DFFPOSX1 ram_reg_29__46_ ( .D(n4814), .CLK(clk), .Q(ram[145]) );
  DFFPOSX1 ram_reg_29__47_ ( .D(n4813), .CLK(clk), .Q(ram[144]) );
  DFFPOSX1 ram_reg_29__48_ ( .D(n4812), .CLK(clk), .Q(ram[143]) );
  DFFPOSX1 ram_reg_29__49_ ( .D(n4811), .CLK(clk), .Q(ram[142]) );
  DFFPOSX1 ram_reg_29__50_ ( .D(n4810), .CLK(clk), .Q(ram[141]) );
  DFFPOSX1 ram_reg_29__51_ ( .D(n4809), .CLK(clk), .Q(ram[140]) );
  DFFPOSX1 ram_reg_29__52_ ( .D(n4808), .CLK(clk), .Q(ram[139]) );
  DFFPOSX1 ram_reg_29__53_ ( .D(n4807), .CLK(clk), .Q(ram[138]) );
  DFFPOSX1 ram_reg_29__54_ ( .D(n4806), .CLK(clk), .Q(ram[137]) );
  DFFPOSX1 ram_reg_29__55_ ( .D(n4805), .CLK(clk), .Q(ram[136]) );
  DFFPOSX1 ram_reg_29__56_ ( .D(n4804), .CLK(clk), .Q(ram[135]) );
  DFFPOSX1 ram_reg_29__57_ ( .D(n4803), .CLK(clk), .Q(ram[134]) );
  DFFPOSX1 ram_reg_29__58_ ( .D(n4802), .CLK(clk), .Q(ram[133]) );
  DFFPOSX1 ram_reg_29__59_ ( .D(n4801), .CLK(clk), .Q(ram[132]) );
  DFFPOSX1 ram_reg_29__60_ ( .D(n4800), .CLK(clk), .Q(ram[131]) );
  DFFPOSX1 ram_reg_29__61_ ( .D(n4799), .CLK(clk), .Q(ram[130]) );
  DFFPOSX1 ram_reg_29__62_ ( .D(n4798), .CLK(clk), .Q(ram[129]) );
  DFFPOSX1 ram_reg_29__63_ ( .D(n4797), .CLK(clk), .Q(ram[128]) );
  DFFPOSX1 ram_reg_30__0_ ( .D(n4796), .CLK(clk), .Q(ram[127]) );
  DFFPOSX1 ram_reg_30__1_ ( .D(n4795), .CLK(clk), .Q(ram[126]) );
  DFFPOSX1 ram_reg_30__2_ ( .D(n4794), .CLK(clk), .Q(ram[125]) );
  DFFPOSX1 ram_reg_30__3_ ( .D(n4793), .CLK(clk), .Q(ram[124]) );
  DFFPOSX1 ram_reg_30__4_ ( .D(n4792), .CLK(clk), .Q(ram[123]) );
  DFFPOSX1 ram_reg_30__5_ ( .D(n4791), .CLK(clk), .Q(ram[122]) );
  DFFPOSX1 ram_reg_30__6_ ( .D(n4790), .CLK(clk), .Q(ram[121]) );
  DFFPOSX1 ram_reg_30__7_ ( .D(n4789), .CLK(clk), .Q(ram[120]) );
  DFFPOSX1 ram_reg_30__8_ ( .D(n4788), .CLK(clk), .Q(ram[119]) );
  DFFPOSX1 ram_reg_30__9_ ( .D(n4787), .CLK(clk), .Q(ram[118]) );
  DFFPOSX1 ram_reg_30__10_ ( .D(n4786), .CLK(clk), .Q(ram[117]) );
  DFFPOSX1 ram_reg_30__11_ ( .D(n4785), .CLK(clk), .Q(ram[116]) );
  DFFPOSX1 ram_reg_30__12_ ( .D(n4784), .CLK(clk), .Q(ram[115]) );
  DFFPOSX1 ram_reg_30__13_ ( .D(n4783), .CLK(clk), .Q(ram[114]) );
  DFFPOSX1 ram_reg_30__14_ ( .D(n4782), .CLK(clk), .Q(ram[113]) );
  DFFPOSX1 ram_reg_30__15_ ( .D(n4781), .CLK(clk), .Q(ram[112]) );
  DFFPOSX1 ram_reg_30__16_ ( .D(n4780), .CLK(clk), .Q(ram[111]) );
  DFFPOSX1 ram_reg_30__17_ ( .D(n4779), .CLK(clk), .Q(ram[110]) );
  DFFPOSX1 ram_reg_30__18_ ( .D(n4778), .CLK(clk), .Q(ram[109]) );
  DFFPOSX1 ram_reg_30__19_ ( .D(n4777), .CLK(clk), .Q(ram[108]) );
  DFFPOSX1 ram_reg_30__20_ ( .D(n4776), .CLK(clk), .Q(ram[107]) );
  DFFPOSX1 ram_reg_30__21_ ( .D(n4775), .CLK(clk), .Q(ram[106]) );
  DFFPOSX1 ram_reg_30__22_ ( .D(n4774), .CLK(clk), .Q(ram[105]) );
  DFFPOSX1 ram_reg_30__23_ ( .D(n4773), .CLK(clk), .Q(ram[104]) );
  DFFPOSX1 ram_reg_30__24_ ( .D(n4772), .CLK(clk), .Q(ram[103]) );
  DFFPOSX1 ram_reg_30__25_ ( .D(n4771), .CLK(clk), .Q(ram[102]) );
  DFFPOSX1 ram_reg_30__26_ ( .D(n4770), .CLK(clk), .Q(ram[101]) );
  DFFPOSX1 ram_reg_30__27_ ( .D(n4769), .CLK(clk), .Q(ram[100]) );
  DFFPOSX1 ram_reg_30__28_ ( .D(n4768), .CLK(clk), .Q(ram[99]) );
  DFFPOSX1 ram_reg_30__29_ ( .D(n4767), .CLK(clk), .Q(ram[98]) );
  DFFPOSX1 ram_reg_30__30_ ( .D(n4766), .CLK(clk), .Q(ram[97]) );
  DFFPOSX1 ram_reg_30__31_ ( .D(n4765), .CLK(clk), .Q(ram[96]) );
  DFFPOSX1 ram_reg_30__32_ ( .D(n4764), .CLK(clk), .Q(ram[95]) );
  DFFPOSX1 ram_reg_30__33_ ( .D(n4763), .CLK(clk), .Q(ram[94]) );
  DFFPOSX1 ram_reg_30__34_ ( .D(n4762), .CLK(clk), .Q(ram[93]) );
  DFFPOSX1 ram_reg_30__35_ ( .D(n4761), .CLK(clk), .Q(ram[92]) );
  DFFPOSX1 ram_reg_30__36_ ( .D(n4760), .CLK(clk), .Q(ram[91]) );
  DFFPOSX1 ram_reg_30__37_ ( .D(n4759), .CLK(clk), .Q(ram[90]) );
  DFFPOSX1 ram_reg_30__38_ ( .D(n4758), .CLK(clk), .Q(ram[89]) );
  DFFPOSX1 ram_reg_30__39_ ( .D(n4757), .CLK(clk), .Q(ram[88]) );
  DFFPOSX1 ram_reg_30__40_ ( .D(n4756), .CLK(clk), .Q(ram[87]) );
  DFFPOSX1 ram_reg_30__41_ ( .D(n4755), .CLK(clk), .Q(ram[86]) );
  DFFPOSX1 ram_reg_30__42_ ( .D(n4754), .CLK(clk), .Q(ram[85]) );
  DFFPOSX1 ram_reg_30__43_ ( .D(n4753), .CLK(clk), .Q(ram[84]) );
  DFFPOSX1 ram_reg_30__44_ ( .D(n4752), .CLK(clk), .Q(ram[83]) );
  DFFPOSX1 ram_reg_30__45_ ( .D(n4751), .CLK(clk), .Q(ram[82]) );
  DFFPOSX1 ram_reg_30__46_ ( .D(n4750), .CLK(clk), .Q(ram[81]) );
  DFFPOSX1 ram_reg_30__47_ ( .D(n4749), .CLK(clk), .Q(ram[80]) );
  DFFPOSX1 ram_reg_30__48_ ( .D(n4748), .CLK(clk), .Q(ram[79]) );
  DFFPOSX1 ram_reg_30__49_ ( .D(n4747), .CLK(clk), .Q(ram[78]) );
  DFFPOSX1 ram_reg_30__50_ ( .D(n4746), .CLK(clk), .Q(ram[77]) );
  DFFPOSX1 ram_reg_30__51_ ( .D(n4745), .CLK(clk), .Q(ram[76]) );
  DFFPOSX1 ram_reg_30__52_ ( .D(n4744), .CLK(clk), .Q(ram[75]) );
  DFFPOSX1 ram_reg_30__53_ ( .D(n4743), .CLK(clk), .Q(ram[74]) );
  DFFPOSX1 ram_reg_30__54_ ( .D(n4742), .CLK(clk), .Q(ram[73]) );
  DFFPOSX1 ram_reg_30__55_ ( .D(n4741), .CLK(clk), .Q(ram[72]) );
  DFFPOSX1 ram_reg_30__56_ ( .D(n4740), .CLK(clk), .Q(ram[71]) );
  DFFPOSX1 ram_reg_30__57_ ( .D(n4739), .CLK(clk), .Q(ram[70]) );
  DFFPOSX1 ram_reg_30__58_ ( .D(n4738), .CLK(clk), .Q(ram[69]) );
  DFFPOSX1 ram_reg_30__59_ ( .D(n4737), .CLK(clk), .Q(ram[68]) );
  DFFPOSX1 ram_reg_30__60_ ( .D(n4736), .CLK(clk), .Q(ram[67]) );
  DFFPOSX1 ram_reg_30__61_ ( .D(n4735), .CLK(clk), .Q(ram[66]) );
  DFFPOSX1 ram_reg_30__62_ ( .D(n4734), .CLK(clk), .Q(ram[65]) );
  DFFPOSX1 ram_reg_30__63_ ( .D(n4733), .CLK(clk), .Q(ram[64]) );
  DFFPOSX1 ram_reg_31__0_ ( .D(n4732), .CLK(clk), .Q(ram[63]) );
  DFFPOSX1 ram_reg_31__1_ ( .D(n4731), .CLK(clk), .Q(ram[62]) );
  DFFPOSX1 ram_reg_31__2_ ( .D(n4730), .CLK(clk), .Q(ram[61]) );
  DFFPOSX1 ram_reg_31__3_ ( .D(n4729), .CLK(clk), .Q(ram[60]) );
  DFFPOSX1 ram_reg_31__4_ ( .D(n4728), .CLK(clk), .Q(ram[59]) );
  DFFPOSX1 ram_reg_31__5_ ( .D(n4727), .CLK(clk), .Q(ram[58]) );
  DFFPOSX1 ram_reg_31__6_ ( .D(n4726), .CLK(clk), .Q(ram[57]) );
  DFFPOSX1 ram_reg_31__7_ ( .D(n4725), .CLK(clk), .Q(ram[56]) );
  DFFPOSX1 ram_reg_31__8_ ( .D(n4724), .CLK(clk), .Q(ram[55]) );
  DFFPOSX1 ram_reg_31__9_ ( .D(n4723), .CLK(clk), .Q(ram[54]) );
  DFFPOSX1 ram_reg_31__10_ ( .D(n4722), .CLK(clk), .Q(ram[53]) );
  DFFPOSX1 ram_reg_31__11_ ( .D(n4721), .CLK(clk), .Q(ram[52]) );
  DFFPOSX1 ram_reg_31__12_ ( .D(n4720), .CLK(clk), .Q(ram[51]) );
  DFFPOSX1 ram_reg_31__13_ ( .D(n4719), .CLK(clk), .Q(ram[50]) );
  DFFPOSX1 ram_reg_31__14_ ( .D(n4718), .CLK(clk), .Q(ram[49]) );
  DFFPOSX1 ram_reg_31__15_ ( .D(n4717), .CLK(clk), .Q(ram[48]) );
  DFFPOSX1 ram_reg_31__16_ ( .D(n4716), .CLK(clk), .Q(ram[47]) );
  DFFPOSX1 ram_reg_31__17_ ( .D(n4715), .CLK(clk), .Q(ram[46]) );
  DFFPOSX1 ram_reg_31__18_ ( .D(n4714), .CLK(clk), .Q(ram[45]) );
  DFFPOSX1 ram_reg_31__19_ ( .D(n4713), .CLK(clk), .Q(ram[44]) );
  DFFPOSX1 ram_reg_31__20_ ( .D(n4712), .CLK(clk), .Q(ram[43]) );
  DFFPOSX1 ram_reg_31__21_ ( .D(n4711), .CLK(clk), .Q(ram[42]) );
  DFFPOSX1 ram_reg_31__22_ ( .D(n4710), .CLK(clk), .Q(ram[41]) );
  DFFPOSX1 ram_reg_31__23_ ( .D(n4709), .CLK(clk), .Q(ram[40]) );
  DFFPOSX1 ram_reg_31__24_ ( .D(n4708), .CLK(clk), .Q(ram[39]) );
  DFFPOSX1 ram_reg_31__25_ ( .D(n4707), .CLK(clk), .Q(ram[38]) );
  DFFPOSX1 ram_reg_31__26_ ( .D(n4706), .CLK(clk), .Q(ram[37]) );
  DFFPOSX1 ram_reg_31__27_ ( .D(n4705), .CLK(clk), .Q(ram[36]) );
  DFFPOSX1 ram_reg_31__28_ ( .D(n4704), .CLK(clk), .Q(ram[35]) );
  DFFPOSX1 ram_reg_31__29_ ( .D(n4703), .CLK(clk), .Q(ram[34]) );
  DFFPOSX1 ram_reg_31__30_ ( .D(n4702), .CLK(clk), .Q(ram[33]) );
  DFFPOSX1 ram_reg_31__31_ ( .D(n4701), .CLK(clk), .Q(ram[32]) );
  DFFPOSX1 ram_reg_31__32_ ( .D(n4700), .CLK(clk), .Q(ram[31]) );
  DFFPOSX1 ram_reg_31__33_ ( .D(n4699), .CLK(clk), .Q(ram[30]) );
  DFFPOSX1 ram_reg_31__34_ ( .D(n4698), .CLK(clk), .Q(ram[29]) );
  DFFPOSX1 ram_reg_31__35_ ( .D(n4697), .CLK(clk), .Q(ram[28]) );
  DFFPOSX1 ram_reg_31__36_ ( .D(n4696), .CLK(clk), .Q(ram[27]) );
  DFFPOSX1 ram_reg_31__37_ ( .D(n4695), .CLK(clk), .Q(ram[26]) );
  DFFPOSX1 ram_reg_31__38_ ( .D(n4694), .CLK(clk), .Q(ram[25]) );
  DFFPOSX1 ram_reg_31__39_ ( .D(n4693), .CLK(clk), .Q(ram[24]) );
  DFFPOSX1 ram_reg_31__40_ ( .D(n4692), .CLK(clk), .Q(ram[23]) );
  DFFPOSX1 ram_reg_31__41_ ( .D(n4691), .CLK(clk), .Q(ram[22]) );
  DFFPOSX1 ram_reg_31__42_ ( .D(n4690), .CLK(clk), .Q(ram[21]) );
  DFFPOSX1 ram_reg_31__43_ ( .D(n4689), .CLK(clk), .Q(ram[20]) );
  DFFPOSX1 ram_reg_31__44_ ( .D(n4688), .CLK(clk), .Q(ram[19]) );
  DFFPOSX1 ram_reg_31__45_ ( .D(n4687), .CLK(clk), .Q(ram[18]) );
  DFFPOSX1 ram_reg_31__46_ ( .D(n4686), .CLK(clk), .Q(ram[17]) );
  DFFPOSX1 ram_reg_31__47_ ( .D(n4685), .CLK(clk), .Q(ram[16]) );
  DFFPOSX1 ram_reg_31__48_ ( .D(n4684), .CLK(clk), .Q(ram[15]) );
  DFFPOSX1 ram_reg_31__49_ ( .D(n4683), .CLK(clk), .Q(ram[14]) );
  DFFPOSX1 ram_reg_31__50_ ( .D(n4682), .CLK(clk), .Q(ram[13]) );
  DFFPOSX1 ram_reg_31__51_ ( .D(n4681), .CLK(clk), .Q(ram[12]) );
  DFFPOSX1 ram_reg_31__52_ ( .D(n4680), .CLK(clk), .Q(ram[11]) );
  DFFPOSX1 ram_reg_31__53_ ( .D(n4679), .CLK(clk), .Q(ram[10]) );
  DFFPOSX1 ram_reg_31__54_ ( .D(n4678), .CLK(clk), .Q(ram[9]) );
  DFFPOSX1 ram_reg_31__55_ ( .D(n4677), .CLK(clk), .Q(ram[8]) );
  DFFPOSX1 ram_reg_31__56_ ( .D(n4676), .CLK(clk), .Q(ram[7]) );
  DFFPOSX1 ram_reg_31__57_ ( .D(n4675), .CLK(clk), .Q(ram[6]) );
  DFFPOSX1 ram_reg_31__58_ ( .D(n4674), .CLK(clk), .Q(ram[5]) );
  DFFPOSX1 ram_reg_31__59_ ( .D(n4673), .CLK(clk), .Q(ram[4]) );
  DFFPOSX1 ram_reg_31__60_ ( .D(n4672), .CLK(clk), .Q(ram[3]) );
  DFFPOSX1 ram_reg_31__61_ ( .D(n4671), .CLK(clk), .Q(ram[2]) );
  DFFPOSX1 ram_reg_31__62_ ( .D(n4670), .CLK(clk), .Q(ram[1]) );
  DFFPOSX1 ram_reg_31__63_ ( .D(n4669), .CLK(clk), .Q(ram[0]) );
  NAND3X1 U3366 ( .A(n10959), .B(n10961), .C(n10957), .Y(n2517) );
  NAND3X1 U3497 ( .A(n10961), .B(n10958), .C(n10959), .Y(n2584) );
  NAND3X1 U3628 ( .A(n10961), .B(n10960), .C(n10957), .Y(n2651) );
  NAND3X1 U3759 ( .A(n10960), .B(n10958), .C(n10961), .Y(n2718) );
  NAND3X1 U3890 ( .A(n10959), .B(n10962), .C(n10957), .Y(n2785) );
  NAND3X1 U4021 ( .A(n10962), .B(n10958), .C(n10959), .Y(n2852) );
  NAND3X1 U4153 ( .A(n10962), .B(n10960), .C(n10957), .Y(n2919) );
  XNOR2X1 U4283 ( .A(read2_addr[3]), .B(n10959), .Y(n4578) );
  XNOR2X1 U4284 ( .A(read2_addr[0]), .B(n4150), .Y(n4577) );
  XNOR2X1 U4285 ( .A(read2_addr[1]), .B(n10963), .Y(n4576) );
  XNOR2X1 U4287 ( .A(read2_addr[2]), .B(n10961), .Y(n4580) );
  XNOR2X1 U4288 ( .A(read2_addr[4]), .B(n10957), .Y(n4579) );
  XNOR2X1 U4487 ( .A(read1_addr[3]), .B(n10959), .Y(n4664) );
  XNOR2X1 U4488 ( .A(read1_addr[0]), .B(n4150), .Y(n4663) );
  XNOR2X1 U4489 ( .A(read1_addr[1]), .B(n10963), .Y(n4662) );
  XNOR2X1 U4491 ( .A(read1_addr[2]), .B(n10961), .Y(n4666) );
  NAND3X1 U4492 ( .A(n10965), .B(n10964), .C(n13229), .Y(n4667) );
  NAND3X1 U4493 ( .A(n10960), .B(n10958), .C(n10962), .Y(n2986) );
  XNOR2X1 U4494 ( .A(read1_addr[4]), .B(n10957), .Y(n4665) );
  INVX2 U3 ( .A(n11110), .Y(n10763) );
  INVX2 U4 ( .A(n11110), .Y(n10764) );
  OR2X2 U5 ( .A(n4), .B(n2150), .Y(n11110) );
  AND2X1 U6 ( .A(write_en), .B(n2), .Y(n4508) );
  AND2X1 U7 ( .A(n1836), .B(n11016), .Y(n2155) );
  AND2X1 U8 ( .A(n2152), .B(n11016), .Y(n2156) );
  AND2X1 U9 ( .A(n11005), .B(n1836), .Y(n2154) );
  AND2X1 U10 ( .A(n11005), .B(n2152), .Y(n2157) );
  OR2X1 U11 ( .A(n3), .B(n2151), .Y(n11043) );
  BUFX2 U12 ( .A(Din[23]), .Y(n1) );
  AND2X1 U13 ( .A(n11112), .B(n11840), .Y(n11905) );
  AND2X1 U14 ( .A(n11112), .B(n12369), .Y(n12434) );
  AND2X1 U15 ( .A(n11112), .B(n12435), .Y(n12500) );
  AND2X1 U16 ( .A(n11112), .B(n12567), .Y(n12632) );
  AND2X1 U17 ( .A(n11112), .B(n12700), .Y(n12765) );
  AND2X1 U18 ( .A(n11112), .B(n12766), .Y(n12831) );
  AND2X1 U19 ( .A(n11112), .B(n12832), .Y(n12897) );
  AND2X1 U20 ( .A(n11112), .B(n12898), .Y(n12963) );
  AND2X1 U21 ( .A(n11112), .B(n13097), .Y(n13225) );
  BUFX2 U22 ( .A(n4667), .Y(n2) );
  BUFX2 U23 ( .A(n10968), .Y(n3) );
  BUFX2 U24 ( .A(n11046), .Y(n4) );
  AND2X1 U25 ( .A(n11112), .B(n12038), .Y(n12103) );
  AND2X1 U26 ( .A(n11112), .B(n11245), .Y(n11310) );
  AND2X1 U27 ( .A(ram[1980]), .B(n10952), .Y(n13218) );
  INVX1 U28 ( .A(n13218), .Y(n5) );
  AND2X1 U29 ( .A(ram[1967]), .B(n10952), .Y(n13192) );
  INVX1 U30 ( .A(n13192), .Y(n6) );
  AND2X1 U31 ( .A(ram[1954]), .B(n10952), .Y(n13166) );
  INVX1 U32 ( .A(n13166), .Y(n7) );
  AND2X1 U33 ( .A(ram[1941]), .B(n10952), .Y(n13140) );
  INVX1 U34 ( .A(n13140), .Y(n8) );
  AND2X1 U35 ( .A(ram[1929]), .B(n10952), .Y(n13116) );
  INVX1 U36 ( .A(n13116), .Y(n9) );
  AND2X1 U37 ( .A(ram[1917]), .B(n10824), .Y(n13092) );
  INVX1 U38 ( .A(n13092), .Y(n10) );
  AND2X1 U39 ( .A(ram[1904]), .B(n10824), .Y(n13079) );
  INVX1 U40 ( .A(n13079), .Y(n11) );
  AND2X1 U41 ( .A(ram[1891]), .B(n10824), .Y(n13066) );
  INVX1 U42 ( .A(n13066), .Y(n12) );
  AND2X1 U43 ( .A(ram[1878]), .B(n10824), .Y(n13053) );
  INVX1 U44 ( .A(n13053), .Y(n13) );
  AND2X1 U45 ( .A(ram[1866]), .B(n10824), .Y(n13041) );
  INVX1 U46 ( .A(n13041), .Y(n14) );
  AND2X1 U47 ( .A(ram[1854]), .B(n10822), .Y(n13027) );
  INVX1 U48 ( .A(n13027), .Y(n15) );
  AND2X1 U49 ( .A(ram[1841]), .B(n10822), .Y(n13014) );
  INVX1 U50 ( .A(n13014), .Y(n16) );
  AND2X1 U51 ( .A(ram[1828]), .B(n10822), .Y(n13001) );
  INVX1 U52 ( .A(n13001), .Y(n17) );
  AND2X1 U53 ( .A(ram[1815]), .B(n10822), .Y(n12988) );
  INVX1 U54 ( .A(n12988), .Y(n18) );
  AND2X1 U55 ( .A(ram[1803]), .B(n10822), .Y(n12976) );
  INVX1 U56 ( .A(n12976), .Y(n34) );
  AND2X1 U57 ( .A(ram[1791]), .B(n10820), .Y(n12962) );
  INVX1 U58 ( .A(n12962), .Y(n35) );
  AND2X1 U59 ( .A(ram[1778]), .B(n10820), .Y(n12949) );
  INVX1 U60 ( .A(n12949), .Y(n36) );
  AND2X1 U61 ( .A(ram[1765]), .B(n10820), .Y(n12936) );
  INVX1 U62 ( .A(n12936), .Y(n37) );
  AND2X1 U63 ( .A(ram[1752]), .B(n10820), .Y(n12923) );
  INVX1 U64 ( .A(n12923), .Y(n38) );
  AND2X1 U65 ( .A(ram[1527]), .B(n10812), .Y(n12690) );
  INVX1 U66 ( .A(n12690), .Y(n39) );
  AND2X1 U67 ( .A(ram[1514]), .B(n10812), .Y(n12677) );
  INVX1 U68 ( .A(n12677), .Y(n40) );
  AND2X1 U69 ( .A(ram[1501]), .B(n10812), .Y(n12664) );
  INVX1 U70 ( .A(n12664), .Y(n41) );
  AND2X1 U71 ( .A(ram[1488]), .B(n10812), .Y(n12651) );
  INVX1 U72 ( .A(n12651), .Y(n42) );
  AND2X1 U73 ( .A(ram[1476]), .B(n10812), .Y(n12639) );
  INVX1 U74 ( .A(n12639), .Y(n43) );
  AND2X1 U75 ( .A(ram[1464]), .B(n10810), .Y(n12624) );
  INVX1 U76 ( .A(n12624), .Y(n44) );
  AND2X1 U77 ( .A(ram[1451]), .B(n10810), .Y(n12611) );
  INVX1 U78 ( .A(n12611), .Y(n45) );
  AND2X1 U79 ( .A(ram[1438]), .B(n10810), .Y(n12598) );
  INVX1 U80 ( .A(n12598), .Y(n46) );
  AND2X1 U81 ( .A(ram[1425]), .B(n10810), .Y(n12585) );
  INVX1 U82 ( .A(n12585), .Y(n47) );
  AND2X1 U83 ( .A(ram[1413]), .B(n10810), .Y(n12573) );
  INVX1 U84 ( .A(n12573), .Y(n48) );
  AND2X1 U85 ( .A(ram[1401]), .B(n10808), .Y(n12559) );
  INVX1 U86 ( .A(n12559), .Y(n49) );
  AND2X1 U87 ( .A(ram[1388]), .B(n10808), .Y(n12546) );
  INVX1 U88 ( .A(n12546), .Y(n50) );
  AND2X1 U89 ( .A(ram[1375]), .B(n10808), .Y(n12533) );
  INVX1 U90 ( .A(n12533), .Y(n51) );
  AND2X1 U91 ( .A(ram[1362]), .B(n10808), .Y(n12520) );
  INVX1 U92 ( .A(n12520), .Y(n52) );
  AND2X1 U93 ( .A(ram[1350]), .B(n10808), .Y(n12508) );
  INVX1 U94 ( .A(n12508), .Y(n53) );
  AND2X1 U95 ( .A(ram[1338]), .B(n10806), .Y(n12494) );
  INVX1 U96 ( .A(n12494), .Y(n54) );
  AND2X1 U97 ( .A(ram[1325]), .B(n10806), .Y(n12481) );
  INVX1 U98 ( .A(n12481), .Y(n55) );
  AND2X1 U99 ( .A(ram[1312]), .B(n10806), .Y(n12468) );
  INVX1 U100 ( .A(n12468), .Y(n120) );
  AND2X1 U101 ( .A(ram[1299]), .B(n10806), .Y(n12455) );
  INVX1 U102 ( .A(n12455), .Y(n121) );
  AND2X1 U103 ( .A(ram[1287]), .B(n10806), .Y(n12443) );
  INVX1 U104 ( .A(n12443), .Y(n122) );
  AND2X1 U105 ( .A(ram[1275]), .B(n10804), .Y(n12429) );
  INVX1 U106 ( .A(n12429), .Y(n187) );
  AND2X1 U107 ( .A(ram[1262]), .B(n10804), .Y(n12416) );
  INVX1 U108 ( .A(n12416), .Y(n188) );
  AND2X1 U109 ( .A(ram[1249]), .B(n10804), .Y(n12403) );
  INVX1 U110 ( .A(n12403), .Y(n189) );
  AND2X1 U111 ( .A(ram[1236]), .B(n10804), .Y(n12390) );
  INVX1 U112 ( .A(n12390), .Y(n190) );
  AND2X1 U113 ( .A(ram[1224]), .B(n10804), .Y(n12378) );
  INVX1 U114 ( .A(n12378), .Y(n191) );
  AND2X1 U115 ( .A(ram[1212]), .B(n10802), .Y(n12364) );
  INVX1 U116 ( .A(n12364), .Y(n192) );
  AND2X1 U117 ( .A(ram[1199]), .B(n10802), .Y(n12351) );
  INVX1 U118 ( .A(n12351), .Y(n193) );
  AND2X1 U119 ( .A(ram[1186]), .B(n10802), .Y(n12338) );
  INVX1 U120 ( .A(n12338), .Y(n194) );
  AND2X1 U121 ( .A(ram[1173]), .B(n10802), .Y(n12325) );
  INVX1 U122 ( .A(n12325), .Y(n195) );
  AND2X1 U123 ( .A(ram[1161]), .B(n10802), .Y(n12313) );
  INVX1 U124 ( .A(n12313), .Y(n196) );
  AND2X1 U125 ( .A(ram[1149]), .B(n10800), .Y(n12299) );
  INVX1 U126 ( .A(n12299), .Y(n197) );
  AND2X1 U127 ( .A(ram[1136]), .B(n10800), .Y(n12286) );
  INVX1 U128 ( .A(n12286), .Y(n198) );
  AND2X1 U129 ( .A(ram[1123]), .B(n10800), .Y(n12273) );
  INVX1 U130 ( .A(n12273), .Y(n199) );
  AND2X1 U131 ( .A(ram[1110]), .B(n10800), .Y(n12260) );
  INVX1 U132 ( .A(n12260), .Y(n200) );
  AND2X1 U133 ( .A(ram[1098]), .B(n10800), .Y(n12248) );
  INVX1 U134 ( .A(n12248), .Y(n201) );
  AND2X1 U135 ( .A(ram[1086]), .B(n10798), .Y(n12234) );
  INVX1 U136 ( .A(n12234), .Y(n202) );
  AND2X1 U137 ( .A(ram[1073]), .B(n10798), .Y(n12221) );
  INVX1 U138 ( .A(n12221), .Y(n203) );
  AND2X1 U139 ( .A(ram[1060]), .B(n10798), .Y(n12208) );
  INVX1 U140 ( .A(n12208), .Y(n204) );
  AND2X1 U141 ( .A(ram[1047]), .B(n10798), .Y(n12195) );
  INVX1 U142 ( .A(n12195), .Y(n205) );
  AND2X1 U143 ( .A(ram[1035]), .B(n10798), .Y(n12183) );
  INVX1 U144 ( .A(n12183), .Y(n206) );
  AND2X1 U145 ( .A(ram[1023]), .B(n10796), .Y(n12169) );
  INVX1 U146 ( .A(n12169), .Y(n207) );
  AND2X1 U147 ( .A(ram[1010]), .B(n10796), .Y(n12156) );
  INVX1 U148 ( .A(n12156), .Y(n208) );
  AND2X1 U149 ( .A(ram[997]), .B(n10796), .Y(n12143) );
  INVX1 U150 ( .A(n12143), .Y(n209) );
  AND2X1 U151 ( .A(ram[984]), .B(n10796), .Y(n12130) );
  INVX1 U152 ( .A(n12130), .Y(n210) );
  AND2X1 U153 ( .A(ram[759]), .B(n10788), .Y(n11896) );
  INVX1 U154 ( .A(n11896), .Y(n211) );
  AND2X1 U155 ( .A(ram[746]), .B(n10788), .Y(n11883) );
  INVX1 U156 ( .A(n11883), .Y(n212) );
  AND2X1 U157 ( .A(ram[733]), .B(n10788), .Y(n11870) );
  INVX1 U158 ( .A(n11870), .Y(n213) );
  AND2X1 U159 ( .A(ram[720]), .B(n10788), .Y(n11857) );
  INVX1 U160 ( .A(n11857), .Y(n214) );
  AND2X1 U161 ( .A(ram[708]), .B(n10788), .Y(n11845) );
  INVX1 U162 ( .A(n11845), .Y(n215) );
  AND2X1 U163 ( .A(ram[696]), .B(n10786), .Y(n11831) );
  INVX1 U164 ( .A(n11831), .Y(n216) );
  AND2X1 U165 ( .A(ram[683]), .B(n10786), .Y(n11818) );
  INVX1 U166 ( .A(n11818), .Y(n217) );
  AND2X1 U167 ( .A(ram[670]), .B(n10786), .Y(n11805) );
  INVX1 U168 ( .A(n11805), .Y(n218) );
  AND2X1 U169 ( .A(ram[657]), .B(n10786), .Y(n11792) );
  INVX1 U170 ( .A(n11792), .Y(n219) );
  AND2X1 U171 ( .A(ram[645]), .B(n10786), .Y(n11780) );
  INVX1 U172 ( .A(n11780), .Y(n220) );
  AND2X1 U173 ( .A(ram[633]), .B(n10784), .Y(n11766) );
  INVX1 U174 ( .A(n11766), .Y(n221) );
  AND2X1 U175 ( .A(ram[620]), .B(n10784), .Y(n11753) );
  INVX1 U176 ( .A(n11753), .Y(n222) );
  AND2X1 U177 ( .A(ram[607]), .B(n10784), .Y(n11740) );
  INVX1 U178 ( .A(n11740), .Y(n223) );
  AND2X1 U179 ( .A(ram[594]), .B(n10784), .Y(n11727) );
  INVX1 U180 ( .A(n11727), .Y(n224) );
  AND2X1 U181 ( .A(ram[582]), .B(n10784), .Y(n11715) );
  INVX1 U182 ( .A(n11715), .Y(n225) );
  AND2X1 U183 ( .A(ram[570]), .B(n10782), .Y(n11701) );
  INVX1 U184 ( .A(n11701), .Y(n226) );
  AND2X1 U185 ( .A(ram[557]), .B(n10782), .Y(n11688) );
  INVX1 U186 ( .A(n11688), .Y(n227) );
  AND2X1 U187 ( .A(ram[544]), .B(n10782), .Y(n11675) );
  INVX1 U188 ( .A(n11675), .Y(n228) );
  AND2X1 U189 ( .A(ram[531]), .B(n10782), .Y(n11662) );
  INVX1 U190 ( .A(n11662), .Y(n229) );
  AND2X1 U191 ( .A(ram[519]), .B(n10782), .Y(n11650) );
  INVX1 U192 ( .A(n11650), .Y(n230) );
  AND2X1 U193 ( .A(ram[507]), .B(n10780), .Y(n11636) );
  INVX1 U194 ( .A(n11636), .Y(n231) );
  AND2X1 U195 ( .A(ram[494]), .B(n10780), .Y(n11623) );
  INVX1 U196 ( .A(n11623), .Y(n232) );
  AND2X1 U197 ( .A(ram[481]), .B(n10780), .Y(n11610) );
  INVX1 U198 ( .A(n11610), .Y(n233) );
  AND2X1 U199 ( .A(ram[468]), .B(n10780), .Y(n11597) );
  INVX1 U200 ( .A(n11597), .Y(n234) );
  AND2X1 U201 ( .A(ram[456]), .B(n10780), .Y(n11585) );
  INVX1 U202 ( .A(n11585), .Y(n235) );
  AND2X1 U203 ( .A(ram[444]), .B(n10778), .Y(n11570) );
  INVX1 U204 ( .A(n11570), .Y(n236) );
  AND2X1 U205 ( .A(ram[431]), .B(n10778), .Y(n11557) );
  INVX1 U206 ( .A(n11557), .Y(n237) );
  AND2X1 U207 ( .A(ram[418]), .B(n10778), .Y(n11544) );
  INVX1 U208 ( .A(n11544), .Y(n238) );
  AND2X1 U209 ( .A(ram[405]), .B(n10778), .Y(n11531) );
  INVX1 U210 ( .A(n11531), .Y(n239) );
  AND2X1 U211 ( .A(ram[393]), .B(n10778), .Y(n11519) );
  INVX1 U212 ( .A(n11519), .Y(n240) );
  AND2X1 U213 ( .A(ram[381]), .B(n10776), .Y(n11505) );
  INVX1 U214 ( .A(n11505), .Y(n241) );
  AND2X1 U215 ( .A(ram[368]), .B(n10776), .Y(n11492) );
  INVX1 U216 ( .A(n11492), .Y(n242) );
  AND2X1 U217 ( .A(ram[355]), .B(n10776), .Y(n11479) );
  INVX1 U218 ( .A(n11479), .Y(n243) );
  AND2X1 U219 ( .A(ram[342]), .B(n10776), .Y(n11466) );
  INVX1 U220 ( .A(n11466), .Y(n244) );
  AND2X1 U221 ( .A(ram[330]), .B(n10776), .Y(n11454) );
  INVX1 U222 ( .A(n11454), .Y(n245) );
  AND2X1 U223 ( .A(ram[318]), .B(n10774), .Y(n11440) );
  INVX1 U224 ( .A(n11440), .Y(n246) );
  AND2X1 U225 ( .A(ram[305]), .B(n10774), .Y(n11427) );
  INVX1 U226 ( .A(n11427), .Y(n247) );
  AND2X1 U227 ( .A(ram[292]), .B(n10774), .Y(n11414) );
  INVX1 U228 ( .A(n11414), .Y(n248) );
  AND2X1 U229 ( .A(ram[279]), .B(n10774), .Y(n11401) );
  INVX1 U230 ( .A(n11401), .Y(n249) );
  AND2X1 U231 ( .A(ram[267]), .B(n10774), .Y(n11389) );
  INVX1 U232 ( .A(n11389), .Y(n250) );
  AND2X1 U233 ( .A(ram[255]), .B(n10772), .Y(n11375) );
  INVX1 U234 ( .A(n11375), .Y(n251) );
  AND2X1 U235 ( .A(ram[242]), .B(n10772), .Y(n11362) );
  INVX1 U236 ( .A(n11362), .Y(n252) );
  AND2X1 U237 ( .A(ram[229]), .B(n10772), .Y(n11349) );
  INVX1 U238 ( .A(n11349), .Y(n253) );
  AND2X1 U239 ( .A(ram[216]), .B(n10772), .Y(n11336) );
  INVX1 U240 ( .A(n11336), .Y(n254) );
  AND2X1 U241 ( .A(n11112), .B(n12105), .Y(n12170) );
  AND2X1 U242 ( .A(n11112), .B(n11311), .Y(n11376) );
  AND2X1 U243 ( .A(ram[1979]), .B(n10952), .Y(n13216) );
  INVX1 U244 ( .A(n13216), .Y(n255) );
  AND2X1 U245 ( .A(ram[1966]), .B(n10952), .Y(n13190) );
  INVX1 U246 ( .A(n13190), .Y(n256) );
  AND2X1 U247 ( .A(ram[1953]), .B(n10952), .Y(n13164) );
  INVX1 U248 ( .A(n13164), .Y(n257) );
  AND2X1 U249 ( .A(ram[1940]), .B(n10952), .Y(n13138) );
  INVX1 U250 ( .A(n13138), .Y(n258) );
  AND2X1 U251 ( .A(ram[1928]), .B(n10952), .Y(n13114) );
  INVX1 U252 ( .A(n13114), .Y(n259) );
  AND2X1 U253 ( .A(ram[1918]), .B(n10824), .Y(n13093) );
  INVX1 U254 ( .A(n13093), .Y(n260) );
  AND2X1 U255 ( .A(ram[1905]), .B(n10824), .Y(n13080) );
  INVX1 U256 ( .A(n13080), .Y(n261) );
  AND2X1 U257 ( .A(ram[1892]), .B(n10824), .Y(n13067) );
  INVX1 U258 ( .A(n13067), .Y(n262) );
  AND2X1 U259 ( .A(ram[1879]), .B(n10824), .Y(n13054) );
  INVX1 U260 ( .A(n13054), .Y(n263) );
  AND2X1 U261 ( .A(ram[1867]), .B(n10824), .Y(n13042) );
  INVX1 U262 ( .A(n13042), .Y(n264) );
  AND2X1 U263 ( .A(ram[1853]), .B(n10822), .Y(n13026) );
  INVX1 U264 ( .A(n13026), .Y(n265) );
  AND2X1 U265 ( .A(ram[1840]), .B(n10822), .Y(n13013) );
  INVX1 U266 ( .A(n13013), .Y(n266) );
  AND2X1 U267 ( .A(ram[1827]), .B(n10822), .Y(n13000) );
  INVX1 U268 ( .A(n13000), .Y(n267) );
  AND2X1 U269 ( .A(ram[1814]), .B(n10822), .Y(n12987) );
  INVX1 U270 ( .A(n12987), .Y(n268) );
  AND2X1 U271 ( .A(ram[1802]), .B(n10822), .Y(n12975) );
  INVX1 U272 ( .A(n12975), .Y(n269) );
  AND2X1 U273 ( .A(ram[1727]), .B(n10818), .Y(n12896) );
  INVX1 U274 ( .A(n12896), .Y(n270) );
  AND2X1 U275 ( .A(ram[1714]), .B(n10818), .Y(n12883) );
  INVX1 U276 ( .A(n12883), .Y(n271) );
  AND2X1 U277 ( .A(ram[1701]), .B(n10818), .Y(n12870) );
  INVX1 U278 ( .A(n12870), .Y(n272) );
  AND2X1 U279 ( .A(ram[1688]), .B(n10818), .Y(n12857) );
  INVX1 U280 ( .A(n12857), .Y(n273) );
  AND2X1 U281 ( .A(ram[1528]), .B(n10812), .Y(n12691) );
  INVX1 U282 ( .A(n12691), .Y(n274) );
  AND2X1 U283 ( .A(ram[1515]), .B(n10812), .Y(n12678) );
  INVX1 U284 ( .A(n12678), .Y(n275) );
  AND2X1 U285 ( .A(ram[1502]), .B(n10812), .Y(n12665) );
  INVX1 U286 ( .A(n12665), .Y(n276) );
  AND2X1 U287 ( .A(ram[1489]), .B(n10812), .Y(n12652) );
  INVX1 U288 ( .A(n12652), .Y(n277) );
  AND2X1 U289 ( .A(ram[1477]), .B(n10812), .Y(n12640) );
  INVX1 U290 ( .A(n12640), .Y(n278) );
  AND2X1 U291 ( .A(ram[1463]), .B(n10810), .Y(n12623) );
  INVX1 U292 ( .A(n12623), .Y(n279) );
  AND2X1 U293 ( .A(ram[1450]), .B(n10810), .Y(n12610) );
  INVX1 U294 ( .A(n12610), .Y(n280) );
  AND2X1 U295 ( .A(ram[1437]), .B(n10810), .Y(n12597) );
  INVX1 U296 ( .A(n12597), .Y(n281) );
  AND2X1 U297 ( .A(ram[1424]), .B(n10810), .Y(n12584) );
  INVX1 U298 ( .A(n12584), .Y(n282) );
  AND2X1 U299 ( .A(ram[1412]), .B(n10810), .Y(n12572) );
  INVX1 U300 ( .A(n12572), .Y(n283) );
  AND2X1 U301 ( .A(ram[1402]), .B(n10808), .Y(n12560) );
  INVX1 U302 ( .A(n12560), .Y(n284) );
  AND2X1 U303 ( .A(ram[1389]), .B(n10808), .Y(n12547) );
  INVX1 U304 ( .A(n12547), .Y(n285) );
  AND2X1 U305 ( .A(ram[1376]), .B(n10808), .Y(n12534) );
  INVX1 U306 ( .A(n12534), .Y(n286) );
  AND2X1 U307 ( .A(ram[1363]), .B(n10808), .Y(n12521) );
  INVX1 U308 ( .A(n12521), .Y(n287) );
  AND2X1 U309 ( .A(ram[1351]), .B(n10808), .Y(n12509) );
  INVX1 U310 ( .A(n12509), .Y(n288) );
  AND2X1 U311 ( .A(ram[1337]), .B(n10806), .Y(n12493) );
  INVX1 U312 ( .A(n12493), .Y(n289) );
  AND2X1 U313 ( .A(ram[1324]), .B(n10806), .Y(n12480) );
  INVX1 U314 ( .A(n12480), .Y(n290) );
  AND2X1 U315 ( .A(ram[1311]), .B(n10806), .Y(n12467) );
  INVX1 U316 ( .A(n12467), .Y(n291) );
  AND2X1 U317 ( .A(ram[1298]), .B(n10806), .Y(n12454) );
  INVX1 U318 ( .A(n12454), .Y(n292) );
  AND2X1 U319 ( .A(ram[1286]), .B(n10806), .Y(n12442) );
  INVX1 U320 ( .A(n12442), .Y(n293) );
  AND2X1 U321 ( .A(ram[1276]), .B(n10804), .Y(n12430) );
  INVX1 U322 ( .A(n12430), .Y(n294) );
  AND2X1 U323 ( .A(ram[1263]), .B(n10804), .Y(n12417) );
  INVX1 U324 ( .A(n12417), .Y(n295) );
  AND2X1 U325 ( .A(ram[1250]), .B(n10804), .Y(n12404) );
  INVX1 U326 ( .A(n12404), .Y(n296) );
  AND2X1 U327 ( .A(ram[1237]), .B(n10804), .Y(n12391) );
  INVX1 U328 ( .A(n12391), .Y(n297) );
  AND2X1 U329 ( .A(ram[1225]), .B(n10804), .Y(n12379) );
  INVX1 U330 ( .A(n12379), .Y(n298) );
  AND2X1 U331 ( .A(ram[1211]), .B(n10802), .Y(n12363) );
  INVX1 U332 ( .A(n12363), .Y(n299) );
  AND2X1 U333 ( .A(ram[1198]), .B(n10802), .Y(n12350) );
  INVX1 U334 ( .A(n12350), .Y(n300) );
  AND2X1 U335 ( .A(ram[1185]), .B(n10802), .Y(n12337) );
  INVX1 U336 ( .A(n12337), .Y(n301) );
  AND2X1 U337 ( .A(ram[1172]), .B(n10802), .Y(n12324) );
  INVX1 U338 ( .A(n12324), .Y(n302) );
  AND2X1 U339 ( .A(ram[1160]), .B(n10802), .Y(n12312) );
  INVX1 U340 ( .A(n12312), .Y(n303) );
  AND2X1 U341 ( .A(ram[1150]), .B(n10800), .Y(n12300) );
  INVX1 U342 ( .A(n12300), .Y(n304) );
  AND2X1 U343 ( .A(ram[1137]), .B(n10800), .Y(n12287) );
  INVX1 U344 ( .A(n12287), .Y(n305) );
  AND2X1 U345 ( .A(ram[1124]), .B(n10800), .Y(n12274) );
  INVX1 U346 ( .A(n12274), .Y(n306) );
  AND2X1 U347 ( .A(ram[1111]), .B(n10800), .Y(n12261) );
  INVX1 U348 ( .A(n12261), .Y(n307) );
  AND2X1 U349 ( .A(ram[1099]), .B(n10800), .Y(n12249) );
  INVX1 U350 ( .A(n12249), .Y(n308) );
  AND2X1 U351 ( .A(ram[1085]), .B(n10798), .Y(n12233) );
  INVX1 U352 ( .A(n12233), .Y(n309) );
  AND2X1 U353 ( .A(ram[1072]), .B(n10798), .Y(n12220) );
  INVX1 U354 ( .A(n12220), .Y(n310) );
  AND2X1 U355 ( .A(ram[1059]), .B(n10798), .Y(n12207) );
  INVX1 U356 ( .A(n12207), .Y(n311) );
  AND2X1 U357 ( .A(ram[1046]), .B(n10798), .Y(n12194) );
  INVX1 U358 ( .A(n12194), .Y(n312) );
  AND2X1 U359 ( .A(ram[1034]), .B(n10798), .Y(n12182) );
  INVX1 U360 ( .A(n12182), .Y(n313) );
  AND2X1 U361 ( .A(ram[959]), .B(n10794), .Y(n12102) );
  INVX1 U362 ( .A(n12102), .Y(n314) );
  AND2X1 U363 ( .A(ram[946]), .B(n10794), .Y(n12089) );
  INVX1 U364 ( .A(n12089), .Y(n315) );
  AND2X1 U365 ( .A(ram[933]), .B(n10794), .Y(n12076) );
  INVX1 U366 ( .A(n12076), .Y(n316) );
  AND2X1 U367 ( .A(ram[920]), .B(n10794), .Y(n12063) );
  INVX1 U368 ( .A(n12063), .Y(n317) );
  AND2X1 U369 ( .A(ram[760]), .B(n10788), .Y(n11897) );
  INVX1 U370 ( .A(n11897), .Y(n318) );
  AND2X1 U371 ( .A(ram[747]), .B(n10788), .Y(n11884) );
  INVX1 U372 ( .A(n11884), .Y(n319) );
  AND2X1 U373 ( .A(ram[734]), .B(n10788), .Y(n11871) );
  INVX1 U374 ( .A(n11871), .Y(n320) );
  AND2X1 U375 ( .A(ram[721]), .B(n10788), .Y(n11858) );
  INVX1 U376 ( .A(n11858), .Y(n321) );
  AND2X1 U377 ( .A(ram[709]), .B(n10788), .Y(n11846) );
  INVX1 U378 ( .A(n11846), .Y(n322) );
  AND2X1 U379 ( .A(ram[695]), .B(n10786), .Y(n11830) );
  INVX1 U380 ( .A(n11830), .Y(n323) );
  AND2X1 U381 ( .A(ram[682]), .B(n10786), .Y(n11817) );
  INVX1 U382 ( .A(n11817), .Y(n324) );
  AND2X1 U383 ( .A(ram[669]), .B(n10786), .Y(n11804) );
  INVX1 U384 ( .A(n11804), .Y(n325) );
  AND2X1 U385 ( .A(ram[656]), .B(n10786), .Y(n11791) );
  INVX1 U386 ( .A(n11791), .Y(n326) );
  AND2X1 U387 ( .A(ram[644]), .B(n10786), .Y(n11779) );
  INVX1 U388 ( .A(n11779), .Y(n327) );
  AND2X1 U389 ( .A(ram[634]), .B(n10784), .Y(n11767) );
  INVX1 U390 ( .A(n11767), .Y(n328) );
  AND2X1 U391 ( .A(ram[621]), .B(n10784), .Y(n11754) );
  INVX1 U392 ( .A(n11754), .Y(n329) );
  AND2X1 U393 ( .A(ram[608]), .B(n10784), .Y(n11741) );
  INVX1 U394 ( .A(n11741), .Y(n330) );
  AND2X1 U395 ( .A(ram[595]), .B(n10784), .Y(n11728) );
  INVX1 U396 ( .A(n11728), .Y(n331) );
  AND2X1 U397 ( .A(ram[583]), .B(n10784), .Y(n11716) );
  INVX1 U398 ( .A(n11716), .Y(n332) );
  AND2X1 U399 ( .A(ram[569]), .B(n10782), .Y(n11700) );
  INVX1 U400 ( .A(n11700), .Y(n333) );
  AND2X1 U401 ( .A(ram[556]), .B(n10782), .Y(n11687) );
  INVX1 U402 ( .A(n11687), .Y(n334) );
  AND2X1 U403 ( .A(ram[543]), .B(n10782), .Y(n11674) );
  INVX1 U404 ( .A(n11674), .Y(n335) );
  AND2X1 U405 ( .A(ram[530]), .B(n10782), .Y(n11661) );
  INVX1 U406 ( .A(n11661), .Y(n336) );
  AND2X1 U407 ( .A(ram[518]), .B(n10782), .Y(n11649) );
  INVX1 U408 ( .A(n11649), .Y(n337) );
  AND2X1 U409 ( .A(ram[508]), .B(n10780), .Y(n11637) );
  INVX1 U410 ( .A(n11637), .Y(n338) );
  AND2X1 U411 ( .A(ram[495]), .B(n10780), .Y(n11624) );
  INVX1 U412 ( .A(n11624), .Y(n339) );
  AND2X1 U413 ( .A(ram[482]), .B(n10780), .Y(n11611) );
  INVX1 U414 ( .A(n11611), .Y(n340) );
  AND2X1 U415 ( .A(ram[469]), .B(n10780), .Y(n11598) );
  INVX1 U416 ( .A(n11598), .Y(n341) );
  AND2X1 U417 ( .A(ram[457]), .B(n10780), .Y(n11586) );
  INVX1 U418 ( .A(n11586), .Y(n342) );
  AND2X1 U419 ( .A(ram[443]), .B(n10778), .Y(n11569) );
  INVX1 U420 ( .A(n11569), .Y(n343) );
  AND2X1 U421 ( .A(ram[430]), .B(n10778), .Y(n11556) );
  INVX1 U422 ( .A(n11556), .Y(n344) );
  AND2X1 U423 ( .A(ram[417]), .B(n10778), .Y(n11543) );
  INVX1 U424 ( .A(n11543), .Y(n345) );
  AND2X1 U425 ( .A(ram[404]), .B(n10778), .Y(n11530) );
  INVX1 U426 ( .A(n11530), .Y(n346) );
  AND2X1 U427 ( .A(ram[392]), .B(n10778), .Y(n11518) );
  INVX1 U428 ( .A(n11518), .Y(n347) );
  AND2X1 U429 ( .A(ram[382]), .B(n10776), .Y(n11506) );
  INVX1 U430 ( .A(n11506), .Y(n348) );
  AND2X1 U431 ( .A(ram[369]), .B(n10776), .Y(n11493) );
  INVX1 U432 ( .A(n11493), .Y(n349) );
  AND2X1 U433 ( .A(ram[356]), .B(n10776), .Y(n11480) );
  INVX1 U434 ( .A(n11480), .Y(n350) );
  AND2X1 U435 ( .A(ram[343]), .B(n10776), .Y(n11467) );
  INVX1 U436 ( .A(n11467), .Y(n351) );
  AND2X1 U437 ( .A(ram[331]), .B(n10776), .Y(n11455) );
  INVX1 U438 ( .A(n11455), .Y(n352) );
  AND2X1 U439 ( .A(ram[317]), .B(n10774), .Y(n11439) );
  INVX1 U440 ( .A(n11439), .Y(n353) );
  AND2X1 U441 ( .A(ram[304]), .B(n10774), .Y(n11426) );
  INVX1 U442 ( .A(n11426), .Y(n354) );
  AND2X1 U443 ( .A(ram[291]), .B(n10774), .Y(n11413) );
  INVX1 U444 ( .A(n11413), .Y(n355) );
  AND2X1 U445 ( .A(ram[278]), .B(n10774), .Y(n11400) );
  INVX1 U446 ( .A(n11400), .Y(n356) );
  AND2X1 U447 ( .A(ram[266]), .B(n10774), .Y(n11388) );
  INVX1 U448 ( .A(n11388), .Y(n357) );
  AND2X1 U449 ( .A(ram[191]), .B(n10770), .Y(n11309) );
  INVX1 U450 ( .A(n11309), .Y(n358) );
  AND2X1 U451 ( .A(ram[178]), .B(n10770), .Y(n11296) );
  INVX1 U452 ( .A(n11296), .Y(n359) );
  AND2X1 U453 ( .A(ram[165]), .B(n10770), .Y(n11283) );
  INVX1 U454 ( .A(n11283), .Y(n360) );
  AND2X1 U455 ( .A(ram[152]), .B(n10770), .Y(n11270) );
  INVX1 U456 ( .A(n11270), .Y(n361) );
  AND2X1 U457 ( .A(n11112), .B(n11906), .Y(n11971) );
  AND2X1 U458 ( .A(n11112), .B(n11113), .Y(n11178) );
  AND2X1 U459 ( .A(ram[1982]), .B(n10952), .Y(n13222) );
  INVX1 U460 ( .A(n13222), .Y(n362) );
  AND2X1 U461 ( .A(ram[1969]), .B(n10952), .Y(n13196) );
  INVX1 U462 ( .A(n13196), .Y(n363) );
  AND2X1 U463 ( .A(ram[1956]), .B(n10952), .Y(n13170) );
  INVX1 U464 ( .A(n13170), .Y(n364) );
  AND2X1 U465 ( .A(ram[1943]), .B(n10952), .Y(n13144) );
  INVX1 U466 ( .A(n13144), .Y(n365) );
  AND2X1 U467 ( .A(ram[1931]), .B(n10952), .Y(n13120) );
  INVX1 U468 ( .A(n13120), .Y(n366) );
  AND2X1 U469 ( .A(ram[1915]), .B(n10824), .Y(n13090) );
  INVX1 U470 ( .A(n13090), .Y(n367) );
  AND2X1 U471 ( .A(ram[1902]), .B(n10824), .Y(n13077) );
  INVX1 U472 ( .A(n13077), .Y(n368) );
  AND2X1 U473 ( .A(ram[1889]), .B(n10824), .Y(n13064) );
  INVX1 U474 ( .A(n13064), .Y(n369) );
  AND2X1 U475 ( .A(ram[1876]), .B(n10824), .Y(n13051) );
  INVX1 U476 ( .A(n13051), .Y(n370) );
  AND2X1 U477 ( .A(ram[1864]), .B(n10824), .Y(n13039) );
  INVX1 U478 ( .A(n13039), .Y(n371) );
  AND2X1 U479 ( .A(ram[1852]), .B(n10822), .Y(n13025) );
  INVX1 U480 ( .A(n13025), .Y(n372) );
  AND2X1 U481 ( .A(ram[1839]), .B(n10822), .Y(n13012) );
  INVX1 U482 ( .A(n13012), .Y(n373) );
  AND2X1 U483 ( .A(ram[1826]), .B(n10822), .Y(n12999) );
  INVX1 U484 ( .A(n12999), .Y(n374) );
  AND2X1 U485 ( .A(ram[1813]), .B(n10822), .Y(n12986) );
  INVX1 U486 ( .A(n12986), .Y(n375) );
  AND2X1 U487 ( .A(ram[1801]), .B(n10822), .Y(n12974) );
  INVX1 U488 ( .A(n12974), .Y(n376) );
  AND2X1 U489 ( .A(ram[1663]), .B(n10816), .Y(n12830) );
  INVX1 U490 ( .A(n12830), .Y(n377) );
  AND2X1 U491 ( .A(ram[1650]), .B(n10816), .Y(n12817) );
  INVX1 U492 ( .A(n12817), .Y(n378) );
  AND2X1 U493 ( .A(ram[1637]), .B(n10816), .Y(n12804) );
  INVX1 U494 ( .A(n12804), .Y(n379) );
  AND2X1 U495 ( .A(ram[1624]), .B(n10816), .Y(n12791) );
  INVX1 U496 ( .A(n12791), .Y(n380) );
  AND2X1 U497 ( .A(ram[1529]), .B(n10812), .Y(n12692) );
  INVX1 U498 ( .A(n12692), .Y(n381) );
  AND2X1 U499 ( .A(ram[1516]), .B(n10812), .Y(n12679) );
  INVX1 U500 ( .A(n12679), .Y(n382) );
  AND2X1 U501 ( .A(ram[1503]), .B(n10812), .Y(n12666) );
  INVX1 U502 ( .A(n12666), .Y(n383) );
  AND2X1 U503 ( .A(ram[1490]), .B(n10812), .Y(n12653) );
  INVX1 U504 ( .A(n12653), .Y(n384) );
  AND2X1 U505 ( .A(ram[1478]), .B(n10812), .Y(n12641) );
  INVX1 U506 ( .A(n12641), .Y(n385) );
  AND2X1 U507 ( .A(ram[1466]), .B(n10810), .Y(n12626) );
  INVX1 U508 ( .A(n12626), .Y(n386) );
  AND2X1 U509 ( .A(ram[1453]), .B(n10810), .Y(n12613) );
  INVX1 U510 ( .A(n12613), .Y(n387) );
  AND2X1 U511 ( .A(ram[1440]), .B(n10810), .Y(n12600) );
  INVX1 U512 ( .A(n12600), .Y(n388) );
  AND2X1 U513 ( .A(ram[1427]), .B(n10810), .Y(n12587) );
  INVX1 U514 ( .A(n12587), .Y(n389) );
  AND2X1 U515 ( .A(ram[1415]), .B(n10810), .Y(n12575) );
  INVX1 U516 ( .A(n12575), .Y(n390) );
  AND2X1 U517 ( .A(ram[1399]), .B(n10808), .Y(n12557) );
  INVX1 U518 ( .A(n12557), .Y(n391) );
  AND2X1 U519 ( .A(ram[1386]), .B(n10808), .Y(n12544) );
  INVX1 U520 ( .A(n12544), .Y(n392) );
  AND2X1 U521 ( .A(ram[1373]), .B(n10808), .Y(n12531) );
  INVX1 U522 ( .A(n12531), .Y(n393) );
  AND2X1 U523 ( .A(ram[1360]), .B(n10808), .Y(n12518) );
  INVX1 U524 ( .A(n12518), .Y(n394) );
  AND2X1 U525 ( .A(ram[1348]), .B(n10808), .Y(n12506) );
  INVX1 U526 ( .A(n12506), .Y(n395) );
  AND2X1 U527 ( .A(ram[1336]), .B(n10806), .Y(n12492) );
  INVX1 U528 ( .A(n12492), .Y(n396) );
  AND2X1 U529 ( .A(ram[1323]), .B(n10806), .Y(n12479) );
  INVX1 U530 ( .A(n12479), .Y(n397) );
  AND2X1 U531 ( .A(ram[1310]), .B(n10806), .Y(n12466) );
  INVX1 U532 ( .A(n12466), .Y(n398) );
  AND2X1 U533 ( .A(ram[1297]), .B(n10806), .Y(n12453) );
  INVX1 U534 ( .A(n12453), .Y(n399) );
  AND2X1 U535 ( .A(ram[1285]), .B(n10806), .Y(n12441) );
  INVX1 U536 ( .A(n12441), .Y(n400) );
  AND2X1 U537 ( .A(ram[1277]), .B(n10804), .Y(n12431) );
  INVX1 U538 ( .A(n12431), .Y(n401) );
  AND2X1 U539 ( .A(ram[1264]), .B(n10804), .Y(n12418) );
  INVX1 U540 ( .A(n12418), .Y(n402) );
  AND2X1 U541 ( .A(ram[1251]), .B(n10804), .Y(n12405) );
  INVX1 U542 ( .A(n12405), .Y(n403) );
  AND2X1 U543 ( .A(ram[1238]), .B(n10804), .Y(n12392) );
  INVX1 U544 ( .A(n12392), .Y(n404) );
  AND2X1 U545 ( .A(ram[1226]), .B(n10804), .Y(n12380) );
  INVX1 U546 ( .A(n12380), .Y(n405) );
  AND2X1 U547 ( .A(ram[1214]), .B(n10802), .Y(n12366) );
  INVX1 U548 ( .A(n12366), .Y(n406) );
  AND2X1 U549 ( .A(ram[1201]), .B(n10802), .Y(n12353) );
  INVX1 U550 ( .A(n12353), .Y(n407) );
  AND2X1 U551 ( .A(ram[1188]), .B(n10802), .Y(n12340) );
  INVX1 U552 ( .A(n12340), .Y(n408) );
  AND2X1 U553 ( .A(ram[1175]), .B(n10802), .Y(n12327) );
  INVX1 U554 ( .A(n12327), .Y(n409) );
  AND2X1 U555 ( .A(ram[1163]), .B(n10802), .Y(n12315) );
  INVX1 U556 ( .A(n12315), .Y(n410) );
  AND2X1 U557 ( .A(ram[1147]), .B(n10800), .Y(n12297) );
  INVX1 U558 ( .A(n12297), .Y(n411) );
  AND2X1 U559 ( .A(ram[1134]), .B(n10800), .Y(n12284) );
  INVX1 U560 ( .A(n12284), .Y(n412) );
  AND2X1 U561 ( .A(ram[1121]), .B(n10800), .Y(n12271) );
  INVX1 U562 ( .A(n12271), .Y(n413) );
  AND2X1 U563 ( .A(ram[1108]), .B(n10800), .Y(n12258) );
  INVX1 U564 ( .A(n12258), .Y(n414) );
  AND2X1 U565 ( .A(ram[1096]), .B(n10800), .Y(n12246) );
  INVX1 U566 ( .A(n12246), .Y(n415) );
  AND2X1 U567 ( .A(ram[1084]), .B(n10798), .Y(n12232) );
  INVX1 U568 ( .A(n12232), .Y(n416) );
  AND2X1 U569 ( .A(ram[1071]), .B(n10798), .Y(n12219) );
  INVX1 U570 ( .A(n12219), .Y(n417) );
  AND2X1 U571 ( .A(ram[1058]), .B(n10798), .Y(n12206) );
  INVX1 U572 ( .A(n12206), .Y(n418) );
  AND2X1 U573 ( .A(ram[1045]), .B(n10798), .Y(n12193) );
  INVX1 U574 ( .A(n12193), .Y(n419) );
  AND2X1 U575 ( .A(ram[1033]), .B(n10798), .Y(n12181) );
  INVX1 U576 ( .A(n12181), .Y(n420) );
  AND2X1 U577 ( .A(ram[895]), .B(n10792), .Y(n12036) );
  INVX1 U578 ( .A(n12036), .Y(n421) );
  AND2X1 U579 ( .A(ram[882]), .B(n10792), .Y(n12023) );
  INVX1 U580 ( .A(n12023), .Y(n422) );
  AND2X1 U581 ( .A(ram[869]), .B(n10792), .Y(n12010) );
  INVX1 U582 ( .A(n12010), .Y(n423) );
  AND2X1 U583 ( .A(ram[856]), .B(n10792), .Y(n11997) );
  INVX1 U584 ( .A(n11997), .Y(n424) );
  AND2X1 U585 ( .A(ram[761]), .B(n10788), .Y(n11898) );
  INVX1 U586 ( .A(n11898), .Y(n425) );
  AND2X1 U587 ( .A(ram[748]), .B(n10788), .Y(n11885) );
  INVX1 U588 ( .A(n11885), .Y(n426) );
  AND2X1 U589 ( .A(ram[735]), .B(n10788), .Y(n11872) );
  INVX1 U590 ( .A(n11872), .Y(n427) );
  AND2X1 U591 ( .A(ram[722]), .B(n10788), .Y(n11859) );
  INVX1 U592 ( .A(n11859), .Y(n428) );
  AND2X1 U593 ( .A(ram[710]), .B(n10788), .Y(n11847) );
  INVX1 U594 ( .A(n11847), .Y(n429) );
  AND2X1 U595 ( .A(ram[698]), .B(n10786), .Y(n11833) );
  INVX1 U596 ( .A(n11833), .Y(n430) );
  AND2X1 U597 ( .A(ram[685]), .B(n10786), .Y(n11820) );
  INVX1 U598 ( .A(n11820), .Y(n431) );
  AND2X1 U599 ( .A(ram[672]), .B(n10786), .Y(n11807) );
  INVX1 U600 ( .A(n11807), .Y(n432) );
  AND2X1 U601 ( .A(ram[659]), .B(n10786), .Y(n11794) );
  INVX1 U602 ( .A(n11794), .Y(n433) );
  AND2X1 U603 ( .A(ram[647]), .B(n10786), .Y(n11782) );
  INVX1 U604 ( .A(n11782), .Y(n434) );
  AND2X1 U605 ( .A(ram[631]), .B(n10784), .Y(n11764) );
  INVX1 U606 ( .A(n11764), .Y(n435) );
  AND2X1 U607 ( .A(ram[618]), .B(n10784), .Y(n11751) );
  INVX1 U608 ( .A(n11751), .Y(n436) );
  AND2X1 U609 ( .A(ram[605]), .B(n10784), .Y(n11738) );
  INVX1 U610 ( .A(n11738), .Y(n437) );
  AND2X1 U611 ( .A(ram[592]), .B(n10784), .Y(n11725) );
  INVX1 U612 ( .A(n11725), .Y(n438) );
  AND2X1 U613 ( .A(ram[580]), .B(n10784), .Y(n11713) );
  INVX1 U614 ( .A(n11713), .Y(n439) );
  AND2X1 U615 ( .A(ram[568]), .B(n10782), .Y(n11699) );
  INVX1 U616 ( .A(n11699), .Y(n440) );
  AND2X1 U617 ( .A(ram[555]), .B(n10782), .Y(n11686) );
  INVX1 U618 ( .A(n11686), .Y(n441) );
  AND2X1 U619 ( .A(ram[542]), .B(n10782), .Y(n11673) );
  INVX1 U620 ( .A(n11673), .Y(n442) );
  AND2X1 U621 ( .A(ram[529]), .B(n10782), .Y(n11660) );
  INVX1 U622 ( .A(n11660), .Y(n443) );
  AND2X1 U623 ( .A(ram[517]), .B(n10782), .Y(n11648) );
  INVX1 U624 ( .A(n11648), .Y(n444) );
  AND2X1 U625 ( .A(ram[509]), .B(n10780), .Y(n11638) );
  INVX1 U626 ( .A(n11638), .Y(n445) );
  AND2X1 U627 ( .A(ram[496]), .B(n10780), .Y(n11625) );
  INVX1 U628 ( .A(n11625), .Y(n446) );
  AND2X1 U629 ( .A(ram[483]), .B(n10780), .Y(n11612) );
  INVX1 U630 ( .A(n11612), .Y(n447) );
  AND2X1 U631 ( .A(ram[470]), .B(n10780), .Y(n11599) );
  INVX1 U632 ( .A(n11599), .Y(n448) );
  AND2X1 U633 ( .A(ram[458]), .B(n10780), .Y(n11587) );
  INVX1 U634 ( .A(n11587), .Y(n449) );
  AND2X1 U635 ( .A(ram[446]), .B(n10778), .Y(n11572) );
  INVX1 U636 ( .A(n11572), .Y(n450) );
  AND2X1 U637 ( .A(ram[433]), .B(n10778), .Y(n11559) );
  INVX1 U638 ( .A(n11559), .Y(n451) );
  AND2X1 U639 ( .A(ram[420]), .B(n10778), .Y(n11546) );
  INVX1 U640 ( .A(n11546), .Y(n452) );
  AND2X1 U641 ( .A(ram[407]), .B(n10778), .Y(n11533) );
  INVX1 U642 ( .A(n11533), .Y(n453) );
  AND2X1 U643 ( .A(ram[395]), .B(n10778), .Y(n11521) );
  INVX1 U644 ( .A(n11521), .Y(n454) );
  AND2X1 U645 ( .A(ram[379]), .B(n10776), .Y(n11503) );
  INVX1 U646 ( .A(n11503), .Y(n455) );
  AND2X1 U647 ( .A(ram[366]), .B(n10776), .Y(n11490) );
  INVX1 U648 ( .A(n11490), .Y(n456) );
  AND2X1 U649 ( .A(ram[353]), .B(n10776), .Y(n11477) );
  INVX1 U650 ( .A(n11477), .Y(n457) );
  AND2X1 U651 ( .A(ram[340]), .B(n10776), .Y(n11464) );
  INVX1 U652 ( .A(n11464), .Y(n458) );
  AND2X1 U653 ( .A(ram[328]), .B(n10776), .Y(n11452) );
  INVX1 U654 ( .A(n11452), .Y(n459) );
  AND2X1 U655 ( .A(ram[316]), .B(n10774), .Y(n11438) );
  INVX1 U656 ( .A(n11438), .Y(n460) );
  AND2X1 U657 ( .A(ram[303]), .B(n10774), .Y(n11425) );
  INVX1 U658 ( .A(n11425), .Y(n461) );
  AND2X1 U659 ( .A(ram[290]), .B(n10774), .Y(n11412) );
  INVX1 U660 ( .A(n11412), .Y(n462) );
  AND2X1 U661 ( .A(ram[277]), .B(n10774), .Y(n11399) );
  INVX1 U662 ( .A(n11399), .Y(n463) );
  AND2X1 U663 ( .A(ram[265]), .B(n10774), .Y(n11387) );
  INVX1 U664 ( .A(n11387), .Y(n464) );
  AND2X1 U665 ( .A(ram[127]), .B(n10768), .Y(n11243) );
  INVX1 U666 ( .A(n11243), .Y(n465) );
  AND2X1 U667 ( .A(ram[114]), .B(n10768), .Y(n11230) );
  INVX1 U668 ( .A(n11230), .Y(n466) );
  AND2X1 U669 ( .A(ram[101]), .B(n10768), .Y(n11217) );
  INVX1 U670 ( .A(n11217), .Y(n467) );
  AND2X1 U671 ( .A(ram[88]), .B(n10768), .Y(n11204) );
  INVX1 U672 ( .A(n11204), .Y(n468) );
  AND2X1 U673 ( .A(n11112), .B(n11972), .Y(n12037) );
  AND2X1 U674 ( .A(n11112), .B(n11179), .Y(n11244) );
  AND2X1 U675 ( .A(ram[1981]), .B(n10952), .Y(n13220) );
  INVX1 U676 ( .A(n13220), .Y(n469) );
  AND2X1 U677 ( .A(ram[1968]), .B(n10952), .Y(n13194) );
  INVX1 U678 ( .A(n13194), .Y(n470) );
  AND2X1 U679 ( .A(ram[1955]), .B(n10952), .Y(n13168) );
  INVX1 U680 ( .A(n13168), .Y(n471) );
  AND2X1 U681 ( .A(ram[1942]), .B(n10952), .Y(n13142) );
  INVX1 U682 ( .A(n13142), .Y(n472) );
  AND2X1 U683 ( .A(ram[1930]), .B(n10952), .Y(n13118) );
  INVX1 U684 ( .A(n13118), .Y(n473) );
  AND2X1 U685 ( .A(ram[1916]), .B(n10824), .Y(n13091) );
  INVX1 U686 ( .A(n13091), .Y(n474) );
  AND2X1 U687 ( .A(ram[1903]), .B(n10824), .Y(n13078) );
  INVX1 U688 ( .A(n13078), .Y(n475) );
  AND2X1 U689 ( .A(ram[1890]), .B(n10824), .Y(n13065) );
  INVX1 U690 ( .A(n13065), .Y(n476) );
  AND2X1 U691 ( .A(ram[1877]), .B(n10824), .Y(n13052) );
  INVX1 U692 ( .A(n13052), .Y(n477) );
  AND2X1 U693 ( .A(ram[1865]), .B(n10824), .Y(n13040) );
  INVX1 U694 ( .A(n13040), .Y(n478) );
  AND2X1 U695 ( .A(ram[1851]), .B(n10822), .Y(n13024) );
  INVX1 U696 ( .A(n13024), .Y(n479) );
  AND2X1 U697 ( .A(ram[1838]), .B(n10822), .Y(n13011) );
  INVX1 U698 ( .A(n13011), .Y(n480) );
  AND2X1 U699 ( .A(ram[1825]), .B(n10822), .Y(n12998) );
  INVX1 U700 ( .A(n12998), .Y(n481) );
  AND2X1 U701 ( .A(ram[1812]), .B(n10822), .Y(n12985) );
  INVX1 U702 ( .A(n12985), .Y(n482) );
  AND2X1 U703 ( .A(ram[1800]), .B(n10822), .Y(n12973) );
  INVX1 U704 ( .A(n12973), .Y(n483) );
  AND2X1 U705 ( .A(ram[1599]), .B(n10814), .Y(n12764) );
  INVX1 U706 ( .A(n12764), .Y(n484) );
  AND2X1 U707 ( .A(ram[1586]), .B(n10814), .Y(n12751) );
  INVX1 U708 ( .A(n12751), .Y(n485) );
  AND2X1 U709 ( .A(ram[1573]), .B(n10814), .Y(n12738) );
  INVX1 U710 ( .A(n12738), .Y(n486) );
  AND2X1 U711 ( .A(ram[1560]), .B(n10814), .Y(n12725) );
  INVX1 U712 ( .A(n12725), .Y(n487) );
  AND2X1 U713 ( .A(ram[1530]), .B(n10812), .Y(n12693) );
  INVX1 U714 ( .A(n12693), .Y(n488) );
  AND2X1 U715 ( .A(ram[1517]), .B(n10812), .Y(n12680) );
  INVX1 U716 ( .A(n12680), .Y(n489) );
  AND2X1 U717 ( .A(ram[1504]), .B(n10812), .Y(n12667) );
  INVX1 U718 ( .A(n12667), .Y(n490) );
  AND2X1 U719 ( .A(ram[1491]), .B(n10812), .Y(n12654) );
  INVX1 U720 ( .A(n12654), .Y(n491) );
  AND2X1 U721 ( .A(ram[1479]), .B(n10812), .Y(n12642) );
  INVX1 U722 ( .A(n12642), .Y(n492) );
  AND2X1 U723 ( .A(ram[1465]), .B(n10810), .Y(n12625) );
  INVX1 U724 ( .A(n12625), .Y(n493) );
  AND2X1 U725 ( .A(ram[1452]), .B(n10810), .Y(n12612) );
  INVX1 U726 ( .A(n12612), .Y(n494) );
  AND2X1 U727 ( .A(ram[1439]), .B(n10810), .Y(n12599) );
  INVX1 U728 ( .A(n12599), .Y(n495) );
  AND2X1 U729 ( .A(ram[1426]), .B(n10810), .Y(n12586) );
  INVX1 U730 ( .A(n12586), .Y(n496) );
  AND2X1 U731 ( .A(ram[1414]), .B(n10810), .Y(n12574) );
  INVX1 U732 ( .A(n12574), .Y(n497) );
  AND2X1 U733 ( .A(ram[1400]), .B(n10808), .Y(n12558) );
  INVX1 U734 ( .A(n12558), .Y(n498) );
  AND2X1 U735 ( .A(ram[1387]), .B(n10808), .Y(n12545) );
  INVX1 U736 ( .A(n12545), .Y(n499) );
  AND2X1 U737 ( .A(ram[1374]), .B(n10808), .Y(n12532) );
  INVX1 U738 ( .A(n12532), .Y(n500) );
  AND2X1 U739 ( .A(ram[1361]), .B(n10808), .Y(n12519) );
  INVX1 U740 ( .A(n12519), .Y(n501) );
  AND2X1 U741 ( .A(ram[1349]), .B(n10808), .Y(n12507) );
  INVX1 U742 ( .A(n12507), .Y(n502) );
  AND2X1 U743 ( .A(ram[1335]), .B(n10806), .Y(n12491) );
  INVX1 U744 ( .A(n12491), .Y(n503) );
  AND2X1 U745 ( .A(ram[1322]), .B(n10806), .Y(n12478) );
  INVX1 U746 ( .A(n12478), .Y(n504) );
  AND2X1 U747 ( .A(ram[1309]), .B(n10806), .Y(n12465) );
  INVX1 U748 ( .A(n12465), .Y(n505) );
  AND2X1 U749 ( .A(ram[1296]), .B(n10806), .Y(n12452) );
  INVX1 U750 ( .A(n12452), .Y(n506) );
  AND2X1 U751 ( .A(ram[1284]), .B(n10806), .Y(n12440) );
  INVX1 U752 ( .A(n12440), .Y(n507) );
  AND2X1 U753 ( .A(ram[1278]), .B(n10804), .Y(n12432) );
  INVX1 U754 ( .A(n12432), .Y(n508) );
  AND2X1 U755 ( .A(ram[1265]), .B(n10804), .Y(n12419) );
  INVX1 U756 ( .A(n12419), .Y(n509) );
  AND2X1 U757 ( .A(ram[1252]), .B(n10804), .Y(n12406) );
  INVX1 U758 ( .A(n12406), .Y(n510) );
  AND2X1 U759 ( .A(ram[1239]), .B(n10804), .Y(n12393) );
  INVX1 U760 ( .A(n12393), .Y(n511) );
  AND2X1 U761 ( .A(ram[1227]), .B(n10804), .Y(n12381) );
  INVX1 U762 ( .A(n12381), .Y(n512) );
  AND2X1 U763 ( .A(ram[1213]), .B(n10802), .Y(n12365) );
  INVX1 U764 ( .A(n12365), .Y(n513) );
  AND2X1 U765 ( .A(ram[1200]), .B(n10802), .Y(n12352) );
  INVX1 U766 ( .A(n12352), .Y(n514) );
  AND2X1 U767 ( .A(ram[1187]), .B(n10802), .Y(n12339) );
  INVX1 U768 ( .A(n12339), .Y(n515) );
  AND2X1 U769 ( .A(ram[1174]), .B(n10802), .Y(n12326) );
  INVX1 U770 ( .A(n12326), .Y(n516) );
  AND2X1 U771 ( .A(ram[1162]), .B(n10802), .Y(n12314) );
  INVX1 U772 ( .A(n12314), .Y(n517) );
  AND2X1 U773 ( .A(ram[1148]), .B(n10800), .Y(n12298) );
  INVX1 U774 ( .A(n12298), .Y(n518) );
  AND2X1 U775 ( .A(ram[1135]), .B(n10800), .Y(n12285) );
  INVX1 U776 ( .A(n12285), .Y(n519) );
  AND2X1 U777 ( .A(ram[1122]), .B(n10800), .Y(n12272) );
  INVX1 U778 ( .A(n12272), .Y(n520) );
  AND2X1 U779 ( .A(ram[1109]), .B(n10800), .Y(n12259) );
  INVX1 U780 ( .A(n12259), .Y(n521) );
  AND2X1 U781 ( .A(ram[1097]), .B(n10800), .Y(n12247) );
  INVX1 U782 ( .A(n12247), .Y(n522) );
  AND2X1 U783 ( .A(ram[1083]), .B(n10798), .Y(n12231) );
  INVX1 U784 ( .A(n12231), .Y(n523) );
  AND2X1 U785 ( .A(ram[1070]), .B(n10798), .Y(n12218) );
  INVX1 U786 ( .A(n12218), .Y(n524) );
  AND2X1 U787 ( .A(ram[1057]), .B(n10798), .Y(n12205) );
  INVX1 U788 ( .A(n12205), .Y(n525) );
  AND2X1 U789 ( .A(ram[1044]), .B(n10798), .Y(n12192) );
  INVX1 U790 ( .A(n12192), .Y(n526) );
  AND2X1 U791 ( .A(ram[1032]), .B(n10798), .Y(n12180) );
  INVX1 U792 ( .A(n12180), .Y(n527) );
  AND2X1 U793 ( .A(ram[831]), .B(n10790), .Y(n11970) );
  INVX1 U794 ( .A(n11970), .Y(n528) );
  AND2X1 U795 ( .A(ram[818]), .B(n10790), .Y(n11957) );
  INVX1 U796 ( .A(n11957), .Y(n529) );
  AND2X1 U797 ( .A(ram[805]), .B(n10790), .Y(n11944) );
  INVX1 U798 ( .A(n11944), .Y(n530) );
  AND2X1 U799 ( .A(ram[792]), .B(n10790), .Y(n11931) );
  INVX1 U800 ( .A(n11931), .Y(n531) );
  AND2X1 U801 ( .A(ram[762]), .B(n10788), .Y(n11899) );
  INVX1 U802 ( .A(n11899), .Y(n532) );
  AND2X1 U803 ( .A(ram[749]), .B(n10788), .Y(n11886) );
  INVX1 U804 ( .A(n11886), .Y(n533) );
  AND2X1 U805 ( .A(ram[736]), .B(n10788), .Y(n11873) );
  INVX1 U806 ( .A(n11873), .Y(n534) );
  AND2X1 U807 ( .A(ram[723]), .B(n10788), .Y(n11860) );
  INVX1 U808 ( .A(n11860), .Y(n535) );
  AND2X1 U809 ( .A(ram[711]), .B(n10788), .Y(n11848) );
  INVX1 U810 ( .A(n11848), .Y(n536) );
  AND2X1 U811 ( .A(ram[697]), .B(n10786), .Y(n11832) );
  INVX1 U812 ( .A(n11832), .Y(n537) );
  AND2X1 U813 ( .A(ram[684]), .B(n10786), .Y(n11819) );
  INVX1 U814 ( .A(n11819), .Y(n538) );
  AND2X1 U815 ( .A(ram[671]), .B(n10786), .Y(n11806) );
  INVX1 U816 ( .A(n11806), .Y(n539) );
  AND2X1 U817 ( .A(ram[658]), .B(n10786), .Y(n11793) );
  INVX1 U818 ( .A(n11793), .Y(n540) );
  AND2X1 U819 ( .A(ram[646]), .B(n10786), .Y(n11781) );
  INVX1 U820 ( .A(n11781), .Y(n541) );
  AND2X1 U821 ( .A(ram[632]), .B(n10784), .Y(n11765) );
  INVX1 U822 ( .A(n11765), .Y(n542) );
  AND2X1 U823 ( .A(ram[619]), .B(n10784), .Y(n11752) );
  INVX1 U824 ( .A(n11752), .Y(n543) );
  AND2X1 U825 ( .A(ram[606]), .B(n10784), .Y(n11739) );
  INVX1 U826 ( .A(n11739), .Y(n544) );
  AND2X1 U827 ( .A(ram[593]), .B(n10784), .Y(n11726) );
  INVX1 U828 ( .A(n11726), .Y(n545) );
  AND2X1 U829 ( .A(ram[581]), .B(n10784), .Y(n11714) );
  INVX1 U830 ( .A(n11714), .Y(n546) );
  AND2X1 U831 ( .A(ram[567]), .B(n10782), .Y(n11698) );
  INVX1 U832 ( .A(n11698), .Y(n547) );
  AND2X1 U833 ( .A(ram[554]), .B(n10782), .Y(n11685) );
  INVX1 U834 ( .A(n11685), .Y(n548) );
  AND2X1 U835 ( .A(ram[541]), .B(n10782), .Y(n11672) );
  INVX1 U836 ( .A(n11672), .Y(n549) );
  AND2X1 U837 ( .A(ram[528]), .B(n10782), .Y(n11659) );
  INVX1 U838 ( .A(n11659), .Y(n550) );
  AND2X1 U839 ( .A(ram[516]), .B(n10782), .Y(n11647) );
  INVX1 U840 ( .A(n11647), .Y(n551) );
  AND2X1 U841 ( .A(ram[510]), .B(n10780), .Y(n11639) );
  INVX1 U842 ( .A(n11639), .Y(n552) );
  AND2X1 U843 ( .A(ram[497]), .B(n10780), .Y(n11626) );
  INVX1 U844 ( .A(n11626), .Y(n553) );
  AND2X1 U845 ( .A(ram[484]), .B(n10780), .Y(n11613) );
  INVX1 U846 ( .A(n11613), .Y(n554) );
  AND2X1 U847 ( .A(ram[471]), .B(n10780), .Y(n11600) );
  INVX1 U848 ( .A(n11600), .Y(n555) );
  AND2X1 U849 ( .A(ram[459]), .B(n10780), .Y(n11588) );
  INVX1 U850 ( .A(n11588), .Y(n556) );
  AND2X1 U851 ( .A(ram[445]), .B(n10778), .Y(n11571) );
  INVX1 U852 ( .A(n11571), .Y(n557) );
  AND2X1 U853 ( .A(ram[432]), .B(n10778), .Y(n11558) );
  INVX1 U854 ( .A(n11558), .Y(n558) );
  AND2X1 U855 ( .A(ram[419]), .B(n10778), .Y(n11545) );
  INVX1 U856 ( .A(n11545), .Y(n559) );
  AND2X1 U857 ( .A(ram[406]), .B(n10778), .Y(n11532) );
  INVX1 U858 ( .A(n11532), .Y(n560) );
  AND2X1 U859 ( .A(ram[394]), .B(n10778), .Y(n11520) );
  INVX1 U860 ( .A(n11520), .Y(n561) );
  AND2X1 U861 ( .A(ram[380]), .B(n10776), .Y(n11504) );
  INVX1 U862 ( .A(n11504), .Y(n562) );
  AND2X1 U863 ( .A(ram[367]), .B(n10776), .Y(n11491) );
  INVX1 U864 ( .A(n11491), .Y(n563) );
  AND2X1 U865 ( .A(ram[354]), .B(n10776), .Y(n11478) );
  INVX1 U866 ( .A(n11478), .Y(n564) );
  AND2X1 U867 ( .A(ram[341]), .B(n10776), .Y(n11465) );
  INVX1 U868 ( .A(n11465), .Y(n565) );
  AND2X1 U869 ( .A(ram[329]), .B(n10776), .Y(n11453) );
  INVX1 U870 ( .A(n11453), .Y(n566) );
  AND2X1 U871 ( .A(ram[315]), .B(n10774), .Y(n11437) );
  INVX1 U872 ( .A(n11437), .Y(n567) );
  AND2X1 U873 ( .A(ram[302]), .B(n10774), .Y(n11424) );
  INVX1 U874 ( .A(n11424), .Y(n568) );
  AND2X1 U875 ( .A(ram[289]), .B(n10774), .Y(n11411) );
  INVX1 U876 ( .A(n11411), .Y(n569) );
  AND2X1 U877 ( .A(ram[276]), .B(n10774), .Y(n11398) );
  INVX1 U878 ( .A(n11398), .Y(n570) );
  AND2X1 U879 ( .A(ram[264]), .B(n10774), .Y(n11386) );
  INVX1 U880 ( .A(n11386), .Y(n571) );
  AND2X1 U881 ( .A(ram[63]), .B(n10766), .Y(n11177) );
  INVX1 U882 ( .A(n11177), .Y(n572) );
  AND2X1 U883 ( .A(ram[50]), .B(n10766), .Y(n11164) );
  INVX1 U884 ( .A(n11164), .Y(n573) );
  AND2X1 U885 ( .A(ram[37]), .B(n10766), .Y(n11151) );
  INVX1 U886 ( .A(n11151), .Y(n574) );
  AND2X1 U887 ( .A(ram[24]), .B(n10766), .Y(n11138) );
  INVX1 U888 ( .A(n11138), .Y(n575) );
  AND2X1 U889 ( .A(n11112), .B(n12303), .Y(n12368) );
  AND2X1 U890 ( .A(n11112), .B(n11509), .Y(n11574) );
  AND2X1 U891 ( .A(ram[1787]), .B(n10820), .Y(n12958) );
  INVX1 U892 ( .A(n12958), .Y(n576) );
  AND2X1 U893 ( .A(ram[1774]), .B(n10820), .Y(n12945) );
  INVX1 U894 ( .A(n12945), .Y(n577) );
  AND2X1 U895 ( .A(ram[1761]), .B(n10820), .Y(n12932) );
  INVX1 U896 ( .A(n12932), .Y(n578) );
  AND2X1 U897 ( .A(ram[1748]), .B(n10820), .Y(n12919) );
  INVX1 U898 ( .A(n12919), .Y(n579) );
  AND2X1 U899 ( .A(ram[1736]), .B(n10820), .Y(n12907) );
  INVX1 U900 ( .A(n12907), .Y(n580) );
  AND2X1 U901 ( .A(ram[1724]), .B(n10818), .Y(n12893) );
  INVX1 U902 ( .A(n12893), .Y(n581) );
  AND2X1 U903 ( .A(ram[1711]), .B(n10818), .Y(n12880) );
  INVX1 U904 ( .A(n12880), .Y(n582) );
  AND2X1 U905 ( .A(ram[1698]), .B(n10818), .Y(n12867) );
  INVX1 U906 ( .A(n12867), .Y(n583) );
  AND2X1 U907 ( .A(ram[1685]), .B(n10818), .Y(n12854) );
  INVX1 U908 ( .A(n12854), .Y(n584) );
  AND2X1 U909 ( .A(ram[1673]), .B(n10818), .Y(n12842) );
  INVX1 U910 ( .A(n12842), .Y(n585) );
  AND2X1 U911 ( .A(ram[1661]), .B(n10816), .Y(n12828) );
  INVX1 U912 ( .A(n12828), .Y(n586) );
  AND2X1 U913 ( .A(ram[1648]), .B(n10816), .Y(n12815) );
  INVX1 U914 ( .A(n12815), .Y(n587) );
  AND2X1 U915 ( .A(ram[1635]), .B(n10816), .Y(n12802) );
  INVX1 U916 ( .A(n12802), .Y(n588) );
  AND2X1 U917 ( .A(ram[1622]), .B(n10816), .Y(n12789) );
  INVX1 U918 ( .A(n12789), .Y(n589) );
  AND2X1 U919 ( .A(ram[1610]), .B(n10816), .Y(n12777) );
  INVX1 U920 ( .A(n12777), .Y(n590) );
  AND2X1 U921 ( .A(ram[1598]), .B(n10814), .Y(n12763) );
  INVX1 U922 ( .A(n12763), .Y(n591) );
  AND2X1 U923 ( .A(ram[1585]), .B(n10814), .Y(n12750) );
  INVX1 U924 ( .A(n12750), .Y(n592) );
  AND2X1 U925 ( .A(ram[1572]), .B(n10814), .Y(n12737) );
  INVX1 U926 ( .A(n12737), .Y(n593) );
  AND2X1 U927 ( .A(ram[1559]), .B(n10814), .Y(n12724) );
  INVX1 U928 ( .A(n12724), .Y(n594) );
  AND2X1 U929 ( .A(ram[1547]), .B(n10814), .Y(n12712) );
  INVX1 U930 ( .A(n12712), .Y(n595) );
  AND2X1 U931 ( .A(ram[1523]), .B(n10812), .Y(n12686) );
  INVX1 U932 ( .A(n12686), .Y(n596) );
  AND2X1 U933 ( .A(ram[1510]), .B(n10812), .Y(n12673) );
  INVX1 U934 ( .A(n12673), .Y(n597) );
  AND2X1 U935 ( .A(ram[1497]), .B(n10812), .Y(n12660) );
  INVX1 U936 ( .A(n12660), .Y(n598) );
  AND2X1 U937 ( .A(ram[1484]), .B(n10812), .Y(n12647) );
  INVX1 U938 ( .A(n12647), .Y(n599) );
  AND2X1 U939 ( .A(ram[1472]), .B(n10812), .Y(n12635) );
  INVX1 U940 ( .A(n12635), .Y(n600) );
  AND2X1 U941 ( .A(ram[1460]), .B(n10810), .Y(n12620) );
  INVX1 U942 ( .A(n12620), .Y(n601) );
  AND2X1 U943 ( .A(ram[1447]), .B(n10810), .Y(n12607) );
  INVX1 U944 ( .A(n12607), .Y(n602) );
  AND2X1 U945 ( .A(ram[1434]), .B(n10810), .Y(n12594) );
  INVX1 U946 ( .A(n12594), .Y(n603) );
  AND2X1 U947 ( .A(ram[1421]), .B(n10810), .Y(n12581) );
  INVX1 U948 ( .A(n12581), .Y(n604) );
  AND2X1 U949 ( .A(ram[1409]), .B(n10810), .Y(n12569) );
  INVX1 U950 ( .A(n12569), .Y(n605) );
  AND2X1 U951 ( .A(ram[1397]), .B(n10808), .Y(n12555) );
  INVX1 U952 ( .A(n12555), .Y(n606) );
  AND2X1 U953 ( .A(ram[1384]), .B(n10808), .Y(n12542) );
  INVX1 U954 ( .A(n12542), .Y(n607) );
  AND2X1 U955 ( .A(ram[1371]), .B(n10808), .Y(n12529) );
  INVX1 U956 ( .A(n12529), .Y(n608) );
  AND2X1 U957 ( .A(ram[1358]), .B(n10808), .Y(n12516) );
  INVX1 U958 ( .A(n12516), .Y(n609) );
  AND2X1 U959 ( .A(ram[1346]), .B(n10808), .Y(n12504) );
  INVX1 U960 ( .A(n12504), .Y(n610) );
  AND2X1 U961 ( .A(ram[1334]), .B(n10806), .Y(n12490) );
  INVX1 U962 ( .A(n12490), .Y(n611) );
  AND2X1 U963 ( .A(ram[1321]), .B(n10806), .Y(n12477) );
  INVX1 U964 ( .A(n12477), .Y(n612) );
  AND2X1 U965 ( .A(ram[1308]), .B(n10806), .Y(n12464) );
  INVX1 U966 ( .A(n12464), .Y(n613) );
  AND2X1 U967 ( .A(ram[1295]), .B(n10806), .Y(n12451) );
  INVX1 U968 ( .A(n12451), .Y(n614) );
  AND2X1 U969 ( .A(ram[1283]), .B(n10806), .Y(n12439) );
  INVX1 U970 ( .A(n12439), .Y(n615) );
  AND2X1 U971 ( .A(ram[1279]), .B(n10804), .Y(n12433) );
  INVX1 U972 ( .A(n12433), .Y(n616) );
  AND2X1 U973 ( .A(ram[1266]), .B(n10804), .Y(n12420) );
  INVX1 U974 ( .A(n12420), .Y(n617) );
  AND2X1 U975 ( .A(ram[1253]), .B(n10804), .Y(n12407) );
  INVX1 U976 ( .A(n12407), .Y(n618) );
  AND2X1 U977 ( .A(ram[1240]), .B(n10804), .Y(n12394) );
  INVX1 U978 ( .A(n12394), .Y(n619) );
  AND2X1 U979 ( .A(ram[1019]), .B(n10796), .Y(n12165) );
  INVX1 U980 ( .A(n12165), .Y(n620) );
  AND2X1 U981 ( .A(ram[1006]), .B(n10796), .Y(n12152) );
  INVX1 U982 ( .A(n12152), .Y(n621) );
  AND2X1 U983 ( .A(ram[993]), .B(n10796), .Y(n12139) );
  INVX1 U984 ( .A(n12139), .Y(n622) );
  AND2X1 U985 ( .A(ram[980]), .B(n10796), .Y(n12126) );
  INVX1 U986 ( .A(n12126), .Y(n623) );
  AND2X1 U987 ( .A(ram[968]), .B(n10796), .Y(n12114) );
  INVX1 U988 ( .A(n12114), .Y(n624) );
  AND2X1 U989 ( .A(ram[956]), .B(n10794), .Y(n12099) );
  INVX1 U990 ( .A(n12099), .Y(n625) );
  AND2X1 U991 ( .A(ram[943]), .B(n10794), .Y(n12086) );
  INVX1 U992 ( .A(n12086), .Y(n626) );
  AND2X1 U993 ( .A(ram[930]), .B(n10794), .Y(n12073) );
  INVX1 U994 ( .A(n12073), .Y(n627) );
  AND2X1 U995 ( .A(ram[917]), .B(n10794), .Y(n12060) );
  INVX1 U996 ( .A(n12060), .Y(n628) );
  AND2X1 U997 ( .A(ram[905]), .B(n10794), .Y(n12048) );
  INVX1 U998 ( .A(n12048), .Y(n629) );
  AND2X1 U999 ( .A(ram[893]), .B(n10792), .Y(n12034) );
  INVX1 U1000 ( .A(n12034), .Y(n630) );
  AND2X1 U1001 ( .A(ram[880]), .B(n10792), .Y(n12021) );
  INVX1 U1002 ( .A(n12021), .Y(n631) );
  AND2X1 U1003 ( .A(ram[867]), .B(n10792), .Y(n12008) );
  INVX1 U1004 ( .A(n12008), .Y(n632) );
  AND2X1 U1005 ( .A(ram[854]), .B(n10792), .Y(n11995) );
  INVX1 U1006 ( .A(n11995), .Y(n633) );
  AND2X1 U1007 ( .A(ram[842]), .B(n10792), .Y(n11983) );
  INVX1 U1008 ( .A(n11983), .Y(n634) );
  AND2X1 U1009 ( .A(ram[830]), .B(n10790), .Y(n11969) );
  INVX1 U1010 ( .A(n11969), .Y(n635) );
  AND2X1 U1011 ( .A(ram[817]), .B(n10790), .Y(n11956) );
  INVX1 U1012 ( .A(n11956), .Y(n636) );
  AND2X1 U1013 ( .A(ram[804]), .B(n10790), .Y(n11943) );
  INVX1 U1014 ( .A(n11943), .Y(n637) );
  AND2X1 U1015 ( .A(ram[791]), .B(n10790), .Y(n11930) );
  INVX1 U1016 ( .A(n11930), .Y(n638) );
  AND2X1 U1017 ( .A(ram[779]), .B(n10790), .Y(n11918) );
  INVX1 U1018 ( .A(n11918), .Y(n639) );
  AND2X1 U1019 ( .A(ram[755]), .B(n10788), .Y(n11892) );
  INVX1 U1020 ( .A(n11892), .Y(n640) );
  AND2X1 U1021 ( .A(ram[742]), .B(n10788), .Y(n11879) );
  INVX1 U1022 ( .A(n11879), .Y(n641) );
  AND2X1 U1023 ( .A(ram[729]), .B(n10788), .Y(n11866) );
  INVX1 U1024 ( .A(n11866), .Y(n642) );
  AND2X1 U1025 ( .A(ram[716]), .B(n10788), .Y(n11853) );
  INVX1 U1026 ( .A(n11853), .Y(n643) );
  AND2X1 U1027 ( .A(ram[704]), .B(n10788), .Y(n11841) );
  INVX1 U1028 ( .A(n11841), .Y(n644) );
  AND2X1 U1029 ( .A(ram[692]), .B(n10786), .Y(n11827) );
  INVX1 U1030 ( .A(n11827), .Y(n645) );
  AND2X1 U1031 ( .A(ram[679]), .B(n10786), .Y(n11814) );
  INVX1 U1032 ( .A(n11814), .Y(n646) );
  AND2X1 U1033 ( .A(ram[666]), .B(n10786), .Y(n11801) );
  INVX1 U1034 ( .A(n11801), .Y(n647) );
  AND2X1 U1035 ( .A(ram[653]), .B(n10786), .Y(n11788) );
  INVX1 U1036 ( .A(n11788), .Y(n648) );
  AND2X1 U1037 ( .A(ram[641]), .B(n10786), .Y(n11776) );
  INVX1 U1038 ( .A(n11776), .Y(n649) );
  AND2X1 U1039 ( .A(ram[629]), .B(n10784), .Y(n11762) );
  INVX1 U1040 ( .A(n11762), .Y(n650) );
  AND2X1 U1041 ( .A(ram[616]), .B(n10784), .Y(n11749) );
  INVX1 U1042 ( .A(n11749), .Y(n651) );
  AND2X1 U1043 ( .A(ram[603]), .B(n10784), .Y(n11736) );
  INVX1 U1044 ( .A(n11736), .Y(n652) );
  AND2X1 U1045 ( .A(ram[590]), .B(n10784), .Y(n11723) );
  INVX1 U1046 ( .A(n11723), .Y(n653) );
  AND2X1 U1047 ( .A(ram[578]), .B(n10784), .Y(n11711) );
  INVX1 U1048 ( .A(n11711), .Y(n654) );
  AND2X1 U1049 ( .A(ram[566]), .B(n10782), .Y(n11697) );
  INVX1 U1050 ( .A(n11697), .Y(n655) );
  AND2X1 U1051 ( .A(ram[553]), .B(n10782), .Y(n11684) );
  INVX1 U1052 ( .A(n11684), .Y(n656) );
  AND2X1 U1053 ( .A(ram[540]), .B(n10782), .Y(n11671) );
  INVX1 U1054 ( .A(n11671), .Y(n657) );
  AND2X1 U1055 ( .A(ram[527]), .B(n10782), .Y(n11658) );
  INVX1 U1056 ( .A(n11658), .Y(n658) );
  AND2X1 U1057 ( .A(ram[515]), .B(n10782), .Y(n11646) );
  INVX1 U1058 ( .A(n11646), .Y(n659) );
  AND2X1 U1059 ( .A(ram[511]), .B(n10780), .Y(n11640) );
  INVX1 U1060 ( .A(n11640), .Y(n660) );
  AND2X1 U1061 ( .A(ram[498]), .B(n10780), .Y(n11627) );
  INVX1 U1062 ( .A(n11627), .Y(n661) );
  AND2X1 U1063 ( .A(ram[485]), .B(n10780), .Y(n11614) );
  INVX1 U1064 ( .A(n11614), .Y(n662) );
  AND2X1 U1065 ( .A(ram[472]), .B(n10780), .Y(n11601) );
  INVX1 U1066 ( .A(n11601), .Y(n663) );
  AND2X1 U1067 ( .A(ram[251]), .B(n10772), .Y(n11371) );
  INVX1 U1068 ( .A(n11371), .Y(n664) );
  AND2X1 U1069 ( .A(ram[238]), .B(n10772), .Y(n11358) );
  INVX1 U1070 ( .A(n11358), .Y(n665) );
  AND2X1 U1071 ( .A(ram[225]), .B(n10772), .Y(n11345) );
  INVX1 U1072 ( .A(n11345), .Y(n666) );
  AND2X1 U1073 ( .A(ram[212]), .B(n10772), .Y(n11332) );
  INVX1 U1074 ( .A(n11332), .Y(n667) );
  AND2X1 U1075 ( .A(ram[200]), .B(n10772), .Y(n11320) );
  INVX1 U1076 ( .A(n11320), .Y(n668) );
  AND2X1 U1077 ( .A(ram[188]), .B(n10770), .Y(n11306) );
  INVX1 U1078 ( .A(n11306), .Y(n669) );
  AND2X1 U1079 ( .A(ram[175]), .B(n10770), .Y(n11293) );
  INVX1 U1080 ( .A(n11293), .Y(n670) );
  AND2X1 U1081 ( .A(ram[162]), .B(n10770), .Y(n11280) );
  INVX1 U1082 ( .A(n11280), .Y(n671) );
  AND2X1 U1083 ( .A(ram[149]), .B(n10770), .Y(n11267) );
  INVX1 U1084 ( .A(n11267), .Y(n672) );
  AND2X1 U1085 ( .A(ram[137]), .B(n10770), .Y(n11255) );
  INVX1 U1086 ( .A(n11255), .Y(n673) );
  AND2X1 U1087 ( .A(ram[125]), .B(n10768), .Y(n11241) );
  INVX1 U1088 ( .A(n11241), .Y(n674) );
  AND2X1 U1089 ( .A(ram[112]), .B(n10768), .Y(n11228) );
  INVX1 U1090 ( .A(n11228), .Y(n675) );
  AND2X1 U1091 ( .A(ram[99]), .B(n10768), .Y(n11215) );
  INVX1 U1092 ( .A(n11215), .Y(n676) );
  AND2X1 U1093 ( .A(ram[86]), .B(n10768), .Y(n11202) );
  INVX1 U1094 ( .A(n11202), .Y(n677) );
  AND2X1 U1095 ( .A(ram[74]), .B(n10768), .Y(n11190) );
  INVX1 U1096 ( .A(n11190), .Y(n678) );
  AND2X1 U1097 ( .A(ram[62]), .B(n10766), .Y(n11176) );
  INVX1 U1098 ( .A(n11176), .Y(n679) );
  AND2X1 U1099 ( .A(ram[49]), .B(n10766), .Y(n11163) );
  INVX1 U1100 ( .A(n11163), .Y(n680) );
  AND2X1 U1101 ( .A(ram[36]), .B(n10766), .Y(n11150) );
  INVX1 U1102 ( .A(n11150), .Y(n681) );
  AND2X1 U1103 ( .A(ram[23]), .B(n10766), .Y(n11137) );
  INVX1 U1104 ( .A(n11137), .Y(n682) );
  AND2X1 U1105 ( .A(ram[11]), .B(n10766), .Y(n11125) );
  INVX1 U1106 ( .A(n11125), .Y(n683) );
  AND2X1 U1107 ( .A(n11112), .B(n12237), .Y(n12302) );
  AND2X1 U1108 ( .A(ram[1983]), .B(n10952), .Y(n13224) );
  INVX1 U1109 ( .A(n13224), .Y(n684) );
  AND2X1 U1110 ( .A(ram[1970]), .B(n10952), .Y(n13198) );
  INVX1 U1111 ( .A(n13198), .Y(n685) );
  AND2X1 U1112 ( .A(ram[1957]), .B(n10952), .Y(n13172) );
  INVX1 U1113 ( .A(n13172), .Y(n686) );
  AND2X1 U1114 ( .A(ram[1944]), .B(n10952), .Y(n13146) );
  INVX1 U1115 ( .A(n13146), .Y(n687) );
  AND2X1 U1116 ( .A(ram[1788]), .B(n10820), .Y(n12959) );
  INVX1 U1117 ( .A(n12959), .Y(n688) );
  AND2X1 U1118 ( .A(ram[1775]), .B(n10820), .Y(n12946) );
  INVX1 U1119 ( .A(n12946), .Y(n689) );
  AND2X1 U1120 ( .A(ram[1762]), .B(n10820), .Y(n12933) );
  INVX1 U1121 ( .A(n12933), .Y(n690) );
  AND2X1 U1122 ( .A(ram[1749]), .B(n10820), .Y(n12920) );
  INVX1 U1123 ( .A(n12920), .Y(n691) );
  AND2X1 U1124 ( .A(ram[1737]), .B(n10820), .Y(n12908) );
  INVX1 U1125 ( .A(n12908), .Y(n692) );
  AND2X1 U1126 ( .A(ram[1723]), .B(n10818), .Y(n12892) );
  INVX1 U1127 ( .A(n12892), .Y(n693) );
  AND2X1 U1128 ( .A(ram[1710]), .B(n10818), .Y(n12879) );
  INVX1 U1129 ( .A(n12879), .Y(n694) );
  AND2X1 U1130 ( .A(ram[1697]), .B(n10818), .Y(n12866) );
  INVX1 U1131 ( .A(n12866), .Y(n695) );
  AND2X1 U1132 ( .A(ram[1684]), .B(n10818), .Y(n12853) );
  INVX1 U1133 ( .A(n12853), .Y(n696) );
  AND2X1 U1134 ( .A(ram[1672]), .B(n10818), .Y(n12841) );
  INVX1 U1135 ( .A(n12841), .Y(n697) );
  AND2X1 U1136 ( .A(ram[1662]), .B(n10816), .Y(n12829) );
  INVX1 U1137 ( .A(n12829), .Y(n698) );
  AND2X1 U1138 ( .A(ram[1649]), .B(n10816), .Y(n12816) );
  INVX1 U1139 ( .A(n12816), .Y(n699) );
  AND2X1 U1140 ( .A(ram[1636]), .B(n10816), .Y(n12803) );
  INVX1 U1141 ( .A(n12803), .Y(n700) );
  AND2X1 U1142 ( .A(ram[1623]), .B(n10816), .Y(n12790) );
  INVX1 U1143 ( .A(n12790), .Y(n701) );
  AND2X1 U1144 ( .A(ram[1611]), .B(n10816), .Y(n12778) );
  INVX1 U1145 ( .A(n12778), .Y(n702) );
  AND2X1 U1146 ( .A(ram[1597]), .B(n10814), .Y(n12762) );
  INVX1 U1147 ( .A(n12762), .Y(n703) );
  AND2X1 U1148 ( .A(ram[1584]), .B(n10814), .Y(n12749) );
  INVX1 U1149 ( .A(n12749), .Y(n704) );
  AND2X1 U1150 ( .A(ram[1571]), .B(n10814), .Y(n12736) );
  INVX1 U1151 ( .A(n12736), .Y(n705) );
  AND2X1 U1152 ( .A(ram[1558]), .B(n10814), .Y(n12723) );
  INVX1 U1153 ( .A(n12723), .Y(n706) );
  AND2X1 U1154 ( .A(ram[1546]), .B(n10814), .Y(n12711) );
  INVX1 U1155 ( .A(n12711), .Y(n707) );
  AND2X1 U1156 ( .A(ram[1524]), .B(n10812), .Y(n12687) );
  INVX1 U1157 ( .A(n12687), .Y(n708) );
  AND2X1 U1158 ( .A(ram[1511]), .B(n10812), .Y(n12674) );
  INVX1 U1159 ( .A(n12674), .Y(n709) );
  AND2X1 U1160 ( .A(ram[1498]), .B(n10812), .Y(n12661) );
  INVX1 U1161 ( .A(n12661), .Y(n710) );
  AND2X1 U1162 ( .A(ram[1485]), .B(n10812), .Y(n12648) );
  INVX1 U1163 ( .A(n12648), .Y(n711) );
  AND2X1 U1164 ( .A(ram[1473]), .B(n10812), .Y(n12636) );
  INVX1 U1165 ( .A(n12636), .Y(n712) );
  AND2X1 U1166 ( .A(ram[1459]), .B(n10810), .Y(n12619) );
  INVX1 U1167 ( .A(n12619), .Y(n713) );
  AND2X1 U1168 ( .A(ram[1446]), .B(n10810), .Y(n12606) );
  INVX1 U1169 ( .A(n12606), .Y(n714) );
  AND2X1 U1170 ( .A(ram[1433]), .B(n10810), .Y(n12593) );
  INVX1 U1171 ( .A(n12593), .Y(n715) );
  AND2X1 U1172 ( .A(ram[1420]), .B(n10810), .Y(n12580) );
  INVX1 U1173 ( .A(n12580), .Y(n716) );
  AND2X1 U1174 ( .A(ram[1408]), .B(n10810), .Y(n12568) );
  INVX1 U1175 ( .A(n12568), .Y(n717) );
  AND2X1 U1176 ( .A(ram[1398]), .B(n10808), .Y(n12556) );
  INVX1 U1177 ( .A(n12556), .Y(n718) );
  AND2X1 U1178 ( .A(ram[1385]), .B(n10808), .Y(n12543) );
  INVX1 U1179 ( .A(n12543), .Y(n719) );
  AND2X1 U1180 ( .A(ram[1372]), .B(n10808), .Y(n12530) );
  INVX1 U1181 ( .A(n12530), .Y(n720) );
  AND2X1 U1182 ( .A(ram[1359]), .B(n10808), .Y(n12517) );
  INVX1 U1183 ( .A(n12517), .Y(n721) );
  AND2X1 U1184 ( .A(ram[1347]), .B(n10808), .Y(n12505) );
  INVX1 U1185 ( .A(n12505), .Y(n722) );
  AND2X1 U1186 ( .A(ram[1333]), .B(n10806), .Y(n12489) );
  INVX1 U1187 ( .A(n12489), .Y(n723) );
  AND2X1 U1188 ( .A(ram[1320]), .B(n10806), .Y(n12476) );
  INVX1 U1189 ( .A(n12476), .Y(n724) );
  AND2X1 U1190 ( .A(ram[1307]), .B(n10806), .Y(n12463) );
  INVX1 U1191 ( .A(n12463), .Y(n725) );
  AND2X1 U1192 ( .A(ram[1294]), .B(n10806), .Y(n12450) );
  INVX1 U1193 ( .A(n12450), .Y(n726) );
  AND2X1 U1194 ( .A(ram[1282]), .B(n10806), .Y(n12438) );
  INVX1 U1195 ( .A(n12438), .Y(n727) );
  AND2X1 U1196 ( .A(ram[1215]), .B(n10802), .Y(n12367) );
  INVX1 U1197 ( .A(n12367), .Y(n728) );
  AND2X1 U1198 ( .A(ram[1202]), .B(n10802), .Y(n12354) );
  INVX1 U1199 ( .A(n12354), .Y(n729) );
  AND2X1 U1200 ( .A(ram[1189]), .B(n10802), .Y(n12341) );
  INVX1 U1201 ( .A(n12341), .Y(n730) );
  AND2X1 U1202 ( .A(ram[1176]), .B(n10802), .Y(n12328) );
  INVX1 U1203 ( .A(n12328), .Y(n731) );
  AND2X1 U1204 ( .A(ram[1020]), .B(n10796), .Y(n12166) );
  INVX1 U1205 ( .A(n12166), .Y(n732) );
  AND2X1 U1206 ( .A(ram[1007]), .B(n10796), .Y(n12153) );
  INVX1 U1207 ( .A(n12153), .Y(n733) );
  AND2X1 U1208 ( .A(ram[994]), .B(n10796), .Y(n12140) );
  INVX1 U1209 ( .A(n12140), .Y(n734) );
  AND2X1 U1210 ( .A(ram[981]), .B(n10796), .Y(n12127) );
  INVX1 U1211 ( .A(n12127), .Y(n735) );
  AND2X1 U1212 ( .A(ram[969]), .B(n10796), .Y(n12115) );
  INVX1 U1213 ( .A(n12115), .Y(n736) );
  AND2X1 U1214 ( .A(ram[955]), .B(n10794), .Y(n12098) );
  INVX1 U1215 ( .A(n12098), .Y(n737) );
  AND2X1 U1216 ( .A(ram[942]), .B(n10794), .Y(n12085) );
  INVX1 U1217 ( .A(n12085), .Y(n738) );
  AND2X1 U1218 ( .A(ram[929]), .B(n10794), .Y(n12072) );
  INVX1 U1219 ( .A(n12072), .Y(n739) );
  AND2X1 U1220 ( .A(ram[916]), .B(n10794), .Y(n12059) );
  INVX1 U1221 ( .A(n12059), .Y(n740) );
  AND2X1 U1222 ( .A(ram[904]), .B(n10794), .Y(n12047) );
  INVX1 U1223 ( .A(n12047), .Y(n741) );
  AND2X1 U1224 ( .A(ram[894]), .B(n10792), .Y(n12035) );
  INVX1 U1225 ( .A(n12035), .Y(n742) );
  AND2X1 U1226 ( .A(ram[881]), .B(n10792), .Y(n12022) );
  INVX1 U1227 ( .A(n12022), .Y(n743) );
  AND2X1 U1228 ( .A(ram[868]), .B(n10792), .Y(n12009) );
  INVX1 U1229 ( .A(n12009), .Y(n744) );
  AND2X1 U1230 ( .A(ram[855]), .B(n10792), .Y(n11996) );
  INVX1 U1231 ( .A(n11996), .Y(n745) );
  AND2X1 U1232 ( .A(ram[843]), .B(n10792), .Y(n11984) );
  INVX1 U1233 ( .A(n11984), .Y(n746) );
  AND2X1 U1234 ( .A(ram[829]), .B(n10790), .Y(n11968) );
  INVX1 U1235 ( .A(n11968), .Y(n747) );
  AND2X1 U1236 ( .A(ram[816]), .B(n10790), .Y(n11955) );
  INVX1 U1237 ( .A(n11955), .Y(n748) );
  AND2X1 U1238 ( .A(ram[803]), .B(n10790), .Y(n11942) );
  INVX1 U1239 ( .A(n11942), .Y(n749) );
  AND2X1 U1240 ( .A(ram[790]), .B(n10790), .Y(n11929) );
  INVX1 U1241 ( .A(n11929), .Y(n750) );
  AND2X1 U1242 ( .A(ram[778]), .B(n10790), .Y(n11917) );
  INVX1 U1243 ( .A(n11917), .Y(n751) );
  AND2X1 U1244 ( .A(ram[756]), .B(n10788), .Y(n11893) );
  INVX1 U1245 ( .A(n11893), .Y(n752) );
  AND2X1 U1246 ( .A(ram[743]), .B(n10788), .Y(n11880) );
  INVX1 U1247 ( .A(n11880), .Y(n753) );
  AND2X1 U1248 ( .A(ram[730]), .B(n10788), .Y(n11867) );
  INVX1 U1249 ( .A(n11867), .Y(n754) );
  AND2X1 U1250 ( .A(ram[717]), .B(n10788), .Y(n11854) );
  INVX1 U1251 ( .A(n11854), .Y(n755) );
  AND2X1 U1252 ( .A(ram[705]), .B(n10788), .Y(n11842) );
  INVX1 U1253 ( .A(n11842), .Y(n756) );
  AND2X1 U1254 ( .A(ram[691]), .B(n10786), .Y(n11826) );
  INVX1 U1255 ( .A(n11826), .Y(n757) );
  AND2X1 U1256 ( .A(ram[678]), .B(n10786), .Y(n11813) );
  INVX1 U1257 ( .A(n11813), .Y(n758) );
  AND2X1 U1258 ( .A(ram[665]), .B(n10786), .Y(n11800) );
  INVX1 U1259 ( .A(n11800), .Y(n759) );
  AND2X1 U1260 ( .A(ram[652]), .B(n10786), .Y(n11787) );
  INVX1 U1261 ( .A(n11787), .Y(n760) );
  AND2X1 U1262 ( .A(ram[640]), .B(n10786), .Y(n11775) );
  INVX1 U1263 ( .A(n11775), .Y(n761) );
  AND2X1 U1264 ( .A(ram[630]), .B(n10784), .Y(n11763) );
  INVX1 U1265 ( .A(n11763), .Y(n762) );
  AND2X1 U1266 ( .A(ram[617]), .B(n10784), .Y(n11750) );
  INVX1 U1267 ( .A(n11750), .Y(n763) );
  AND2X1 U1268 ( .A(ram[604]), .B(n10784), .Y(n11737) );
  INVX1 U1269 ( .A(n11737), .Y(n764) );
  AND2X1 U1270 ( .A(ram[591]), .B(n10784), .Y(n11724) );
  INVX1 U1271 ( .A(n11724), .Y(n765) );
  AND2X1 U1272 ( .A(ram[579]), .B(n10784), .Y(n11712) );
  INVX1 U1273 ( .A(n11712), .Y(n766) );
  AND2X1 U1274 ( .A(ram[565]), .B(n10782), .Y(n11696) );
  INVX1 U1275 ( .A(n11696), .Y(n767) );
  AND2X1 U1276 ( .A(ram[552]), .B(n10782), .Y(n11683) );
  INVX1 U1277 ( .A(n11683), .Y(n768) );
  AND2X1 U1278 ( .A(ram[539]), .B(n10782), .Y(n11670) );
  INVX1 U1279 ( .A(n11670), .Y(n769) );
  AND2X1 U1280 ( .A(ram[526]), .B(n10782), .Y(n11657) );
  INVX1 U1281 ( .A(n11657), .Y(n770) );
  AND2X1 U1282 ( .A(ram[514]), .B(n10782), .Y(n11645) );
  INVX1 U1283 ( .A(n11645), .Y(n771) );
  AND2X1 U1284 ( .A(ram[447]), .B(n10778), .Y(n11573) );
  INVX1 U1285 ( .A(n11573), .Y(n772) );
  AND2X1 U1286 ( .A(ram[434]), .B(n10778), .Y(n11560) );
  INVX1 U1287 ( .A(n11560), .Y(n773) );
  AND2X1 U1288 ( .A(ram[421]), .B(n10778), .Y(n11547) );
  INVX1 U1289 ( .A(n11547), .Y(n774) );
  AND2X1 U1290 ( .A(ram[408]), .B(n10778), .Y(n11534) );
  INVX1 U1291 ( .A(n11534), .Y(n775) );
  AND2X1 U1292 ( .A(ram[252]), .B(n10772), .Y(n11372) );
  INVX1 U1293 ( .A(n11372), .Y(n776) );
  AND2X1 U1294 ( .A(ram[239]), .B(n10772), .Y(n11359) );
  INVX1 U1295 ( .A(n11359), .Y(n777) );
  AND2X1 U1296 ( .A(ram[226]), .B(n10772), .Y(n11346) );
  INVX1 U1297 ( .A(n11346), .Y(n778) );
  AND2X1 U1298 ( .A(ram[213]), .B(n10772), .Y(n11333) );
  INVX1 U1299 ( .A(n11333), .Y(n779) );
  AND2X1 U1300 ( .A(ram[201]), .B(n10772), .Y(n11321) );
  INVX1 U1301 ( .A(n11321), .Y(n780) );
  AND2X1 U1302 ( .A(ram[187]), .B(n10770), .Y(n11305) );
  INVX1 U1303 ( .A(n11305), .Y(n781) );
  AND2X1 U1304 ( .A(ram[174]), .B(n10770), .Y(n11292) );
  INVX1 U1305 ( .A(n11292), .Y(n782) );
  AND2X1 U1306 ( .A(ram[161]), .B(n10770), .Y(n11279) );
  INVX1 U1307 ( .A(n11279), .Y(n783) );
  AND2X1 U1308 ( .A(ram[148]), .B(n10770), .Y(n11266) );
  INVX1 U1309 ( .A(n11266), .Y(n784) );
  AND2X1 U1310 ( .A(ram[136]), .B(n10770), .Y(n11254) );
  INVX1 U1311 ( .A(n11254), .Y(n785) );
  AND2X1 U1312 ( .A(ram[126]), .B(n10768), .Y(n11242) );
  INVX1 U1313 ( .A(n11242), .Y(n786) );
  AND2X1 U1314 ( .A(ram[113]), .B(n10768), .Y(n11229) );
  INVX1 U1315 ( .A(n11229), .Y(n787) );
  AND2X1 U1316 ( .A(ram[100]), .B(n10768), .Y(n11216) );
  INVX1 U1317 ( .A(n11216), .Y(n788) );
  AND2X1 U1318 ( .A(ram[87]), .B(n10768), .Y(n11203) );
  INVX1 U1319 ( .A(n11203), .Y(n789) );
  AND2X1 U1320 ( .A(ram[75]), .B(n10768), .Y(n11191) );
  INVX1 U1321 ( .A(n11191), .Y(n790) );
  AND2X1 U1322 ( .A(ram[61]), .B(n10766), .Y(n11175) );
  INVX1 U1323 ( .A(n11175), .Y(n791) );
  AND2X1 U1324 ( .A(ram[48]), .B(n10766), .Y(n11162) );
  INVX1 U1325 ( .A(n11162), .Y(n792) );
  AND2X1 U1326 ( .A(ram[35]), .B(n10766), .Y(n11149) );
  INVX1 U1327 ( .A(n11149), .Y(n793) );
  AND2X1 U1328 ( .A(ram[22]), .B(n10766), .Y(n11136) );
  INVX1 U1329 ( .A(n11136), .Y(n794) );
  AND2X1 U1330 ( .A(ram[10]), .B(n10766), .Y(n11124) );
  INVX1 U1331 ( .A(n11124), .Y(n795) );
  AND2X1 U1332 ( .A(n11112), .B(n12964), .Y(n13029) );
  AND2X1 U1333 ( .A(n11112), .B(n12171), .Y(n12236) );
  AND2X1 U1334 ( .A(n11112), .B(n11377), .Y(n11442) );
  AND2X1 U1335 ( .A(ram[1919]), .B(n10824), .Y(n13094) );
  INVX1 U1336 ( .A(n13094), .Y(n796) );
  AND2X1 U1337 ( .A(ram[1906]), .B(n10824), .Y(n13081) );
  INVX1 U1338 ( .A(n13081), .Y(n797) );
  AND2X1 U1339 ( .A(ram[1893]), .B(n10824), .Y(n13068) );
  INVX1 U1340 ( .A(n13068), .Y(n798) );
  AND2X1 U1341 ( .A(ram[1880]), .B(n10824), .Y(n13055) );
  INVX1 U1342 ( .A(n13055), .Y(n799) );
  AND2X1 U1343 ( .A(ram[1789]), .B(n10820), .Y(n12960) );
  INVX1 U1344 ( .A(n12960), .Y(n800) );
  AND2X1 U1345 ( .A(ram[1776]), .B(n10820), .Y(n12947) );
  INVX1 U1346 ( .A(n12947), .Y(n801) );
  AND2X1 U1347 ( .A(ram[1763]), .B(n10820), .Y(n12934) );
  INVX1 U1348 ( .A(n12934), .Y(n802) );
  AND2X1 U1349 ( .A(ram[1750]), .B(n10820), .Y(n12921) );
  INVX1 U1350 ( .A(n12921), .Y(n803) );
  AND2X1 U1351 ( .A(ram[1738]), .B(n10820), .Y(n12909) );
  INVX1 U1352 ( .A(n12909), .Y(n804) );
  AND2X1 U1353 ( .A(ram[1726]), .B(n10818), .Y(n12895) );
  INVX1 U1354 ( .A(n12895), .Y(n805) );
  AND2X1 U1355 ( .A(ram[1713]), .B(n10818), .Y(n12882) );
  INVX1 U1356 ( .A(n12882), .Y(n806) );
  AND2X1 U1357 ( .A(ram[1700]), .B(n10818), .Y(n12869) );
  INVX1 U1358 ( .A(n12869), .Y(n807) );
  AND2X1 U1359 ( .A(ram[1687]), .B(n10818), .Y(n12856) );
  INVX1 U1360 ( .A(n12856), .Y(n808) );
  AND2X1 U1361 ( .A(ram[1675]), .B(n10818), .Y(n12844) );
  INVX1 U1362 ( .A(n12844), .Y(n809) );
  AND2X1 U1363 ( .A(ram[1659]), .B(n10816), .Y(n12826) );
  INVX1 U1364 ( .A(n12826), .Y(n810) );
  AND2X1 U1365 ( .A(ram[1646]), .B(n10816), .Y(n12813) );
  INVX1 U1366 ( .A(n12813), .Y(n811) );
  AND2X1 U1367 ( .A(ram[1633]), .B(n10816), .Y(n12800) );
  INVX1 U1368 ( .A(n12800), .Y(n812) );
  AND2X1 U1369 ( .A(ram[1620]), .B(n10816), .Y(n12787) );
  INVX1 U1370 ( .A(n12787), .Y(n813) );
  AND2X1 U1371 ( .A(ram[1608]), .B(n10816), .Y(n12775) );
  INVX1 U1372 ( .A(n12775), .Y(n814) );
  AND2X1 U1373 ( .A(ram[1596]), .B(n10814), .Y(n12761) );
  INVX1 U1374 ( .A(n12761), .Y(n815) );
  AND2X1 U1375 ( .A(ram[1583]), .B(n10814), .Y(n12748) );
  INVX1 U1376 ( .A(n12748), .Y(n816) );
  AND2X1 U1377 ( .A(ram[1570]), .B(n10814), .Y(n12735) );
  INVX1 U1378 ( .A(n12735), .Y(n817) );
  AND2X1 U1379 ( .A(ram[1557]), .B(n10814), .Y(n12722) );
  INVX1 U1380 ( .A(n12722), .Y(n818) );
  AND2X1 U1381 ( .A(ram[1545]), .B(n10814), .Y(n12710) );
  INVX1 U1382 ( .A(n12710), .Y(n819) );
  AND2X1 U1383 ( .A(ram[1525]), .B(n10812), .Y(n12688) );
  INVX1 U1384 ( .A(n12688), .Y(n820) );
  AND2X1 U1385 ( .A(ram[1512]), .B(n10812), .Y(n12675) );
  INVX1 U1386 ( .A(n12675), .Y(n821) );
  AND2X1 U1387 ( .A(ram[1499]), .B(n10812), .Y(n12662) );
  INVX1 U1388 ( .A(n12662), .Y(n822) );
  AND2X1 U1389 ( .A(ram[1486]), .B(n10812), .Y(n12649) );
  INVX1 U1390 ( .A(n12649), .Y(n823) );
  AND2X1 U1391 ( .A(ram[1474]), .B(n10812), .Y(n12637) );
  INVX1 U1392 ( .A(n12637), .Y(n824) );
  AND2X1 U1393 ( .A(ram[1462]), .B(n10810), .Y(n12622) );
  INVX1 U1394 ( .A(n12622), .Y(n825) );
  AND2X1 U1395 ( .A(ram[1449]), .B(n10810), .Y(n12609) );
  INVX1 U1396 ( .A(n12609), .Y(n826) );
  AND2X1 U1397 ( .A(ram[1436]), .B(n10810), .Y(n12596) );
  INVX1 U1398 ( .A(n12596), .Y(n827) );
  AND2X1 U1399 ( .A(ram[1423]), .B(n10810), .Y(n12583) );
  INVX1 U1400 ( .A(n12583), .Y(n828) );
  AND2X1 U1401 ( .A(ram[1411]), .B(n10810), .Y(n12571) );
  INVX1 U1402 ( .A(n12571), .Y(n829) );
  AND2X1 U1403 ( .A(ram[1395]), .B(n10808), .Y(n12553) );
  INVX1 U1404 ( .A(n12553), .Y(n830) );
  AND2X1 U1405 ( .A(ram[1382]), .B(n10808), .Y(n12540) );
  INVX1 U1406 ( .A(n12540), .Y(n831) );
  AND2X1 U1407 ( .A(ram[1369]), .B(n10808), .Y(n12527) );
  INVX1 U1408 ( .A(n12527), .Y(n832) );
  AND2X1 U1409 ( .A(ram[1356]), .B(n10808), .Y(n12514) );
  INVX1 U1410 ( .A(n12514), .Y(n833) );
  AND2X1 U1411 ( .A(ram[1344]), .B(n10808), .Y(n12502) );
  INVX1 U1412 ( .A(n12502), .Y(n834) );
  AND2X1 U1413 ( .A(ram[1332]), .B(n10806), .Y(n12488) );
  INVX1 U1414 ( .A(n12488), .Y(n835) );
  AND2X1 U1415 ( .A(ram[1319]), .B(n10806), .Y(n12475) );
  INVX1 U1416 ( .A(n12475), .Y(n836) );
  AND2X1 U1417 ( .A(ram[1306]), .B(n10806), .Y(n12462) );
  INVX1 U1418 ( .A(n12462), .Y(n837) );
  AND2X1 U1419 ( .A(ram[1293]), .B(n10806), .Y(n12449) );
  INVX1 U1420 ( .A(n12449), .Y(n838) );
  AND2X1 U1421 ( .A(ram[1281]), .B(n10806), .Y(n12437) );
  INVX1 U1422 ( .A(n12437), .Y(n839) );
  AND2X1 U1423 ( .A(ram[1151]), .B(n10800), .Y(n12301) );
  INVX1 U1424 ( .A(n12301), .Y(n840) );
  AND2X1 U1425 ( .A(ram[1138]), .B(n10800), .Y(n12288) );
  INVX1 U1426 ( .A(n12288), .Y(n841) );
  AND2X1 U1427 ( .A(ram[1125]), .B(n10800), .Y(n12275) );
  INVX1 U1428 ( .A(n12275), .Y(n842) );
  AND2X1 U1429 ( .A(ram[1112]), .B(n10800), .Y(n12262) );
  INVX1 U1430 ( .A(n12262), .Y(n843) );
  AND2X1 U1431 ( .A(ram[1021]), .B(n10796), .Y(n12167) );
  INVX1 U1432 ( .A(n12167), .Y(n844) );
  AND2X1 U1433 ( .A(ram[1008]), .B(n10796), .Y(n12154) );
  INVX1 U1434 ( .A(n12154), .Y(n845) );
  AND2X1 U1435 ( .A(ram[995]), .B(n10796), .Y(n12141) );
  INVX1 U1436 ( .A(n12141), .Y(n846) );
  AND2X1 U1437 ( .A(ram[982]), .B(n10796), .Y(n12128) );
  INVX1 U1438 ( .A(n12128), .Y(n847) );
  AND2X1 U1439 ( .A(ram[970]), .B(n10796), .Y(n12116) );
  INVX1 U1440 ( .A(n12116), .Y(n848) );
  AND2X1 U1441 ( .A(ram[958]), .B(n10794), .Y(n12101) );
  INVX1 U1442 ( .A(n12101), .Y(n849) );
  AND2X1 U1443 ( .A(ram[945]), .B(n10794), .Y(n12088) );
  INVX1 U1444 ( .A(n12088), .Y(n850) );
  AND2X1 U1445 ( .A(ram[932]), .B(n10794), .Y(n12075) );
  INVX1 U1446 ( .A(n12075), .Y(n851) );
  AND2X1 U1447 ( .A(ram[919]), .B(n10794), .Y(n12062) );
  INVX1 U1448 ( .A(n12062), .Y(n852) );
  AND2X1 U1449 ( .A(ram[907]), .B(n10794), .Y(n12050) );
  INVX1 U1450 ( .A(n12050), .Y(n853) );
  AND2X1 U1451 ( .A(ram[891]), .B(n10792), .Y(n12032) );
  INVX1 U1452 ( .A(n12032), .Y(n854) );
  AND2X1 U1453 ( .A(ram[878]), .B(n10792), .Y(n12019) );
  INVX1 U1454 ( .A(n12019), .Y(n855) );
  AND2X1 U1455 ( .A(ram[865]), .B(n10792), .Y(n12006) );
  INVX1 U1456 ( .A(n12006), .Y(n856) );
  AND2X1 U1457 ( .A(ram[852]), .B(n10792), .Y(n11993) );
  INVX1 U1458 ( .A(n11993), .Y(n857) );
  AND2X1 U1459 ( .A(ram[840]), .B(n10792), .Y(n11981) );
  INVX1 U1460 ( .A(n11981), .Y(n858) );
  AND2X1 U1461 ( .A(ram[828]), .B(n10790), .Y(n11967) );
  INVX1 U1462 ( .A(n11967), .Y(n859) );
  AND2X1 U1463 ( .A(ram[815]), .B(n10790), .Y(n11954) );
  INVX1 U1464 ( .A(n11954), .Y(n860) );
  AND2X1 U1465 ( .A(ram[802]), .B(n10790), .Y(n11941) );
  INVX1 U1466 ( .A(n11941), .Y(n861) );
  AND2X1 U1467 ( .A(ram[789]), .B(n10790), .Y(n11928) );
  INVX1 U1468 ( .A(n11928), .Y(n862) );
  AND2X1 U1469 ( .A(ram[777]), .B(n10790), .Y(n11916) );
  INVX1 U1470 ( .A(n11916), .Y(n863) );
  AND2X1 U1471 ( .A(ram[757]), .B(n10788), .Y(n11894) );
  INVX1 U1472 ( .A(n11894), .Y(n864) );
  AND2X1 U1473 ( .A(ram[744]), .B(n10788), .Y(n11881) );
  INVX1 U1474 ( .A(n11881), .Y(n865) );
  AND2X1 U1475 ( .A(ram[731]), .B(n10788), .Y(n11868) );
  INVX1 U1476 ( .A(n11868), .Y(n866) );
  AND2X1 U1477 ( .A(ram[718]), .B(n10788), .Y(n11855) );
  INVX1 U1478 ( .A(n11855), .Y(n867) );
  AND2X1 U1479 ( .A(ram[706]), .B(n10788), .Y(n11843) );
  INVX1 U1480 ( .A(n11843), .Y(n868) );
  AND2X1 U1481 ( .A(ram[694]), .B(n10786), .Y(n11829) );
  INVX1 U1482 ( .A(n11829), .Y(n869) );
  AND2X1 U1483 ( .A(ram[681]), .B(n10786), .Y(n11816) );
  INVX1 U1484 ( .A(n11816), .Y(n870) );
  AND2X1 U1485 ( .A(ram[668]), .B(n10786), .Y(n11803) );
  INVX1 U1486 ( .A(n11803), .Y(n871) );
  AND2X1 U1487 ( .A(ram[655]), .B(n10786), .Y(n11790) );
  INVX1 U1488 ( .A(n11790), .Y(n872) );
  AND2X1 U1489 ( .A(ram[643]), .B(n10786), .Y(n11778) );
  INVX1 U1490 ( .A(n11778), .Y(n873) );
  AND2X1 U1491 ( .A(ram[627]), .B(n10784), .Y(n11760) );
  INVX1 U1492 ( .A(n11760), .Y(n874) );
  AND2X1 U1493 ( .A(ram[614]), .B(n10784), .Y(n11747) );
  INVX1 U1494 ( .A(n11747), .Y(n875) );
  AND2X1 U1495 ( .A(ram[601]), .B(n10784), .Y(n11734) );
  INVX1 U1496 ( .A(n11734), .Y(n876) );
  AND2X1 U1497 ( .A(ram[588]), .B(n10784), .Y(n11721) );
  INVX1 U1498 ( .A(n11721), .Y(n877) );
  AND2X1 U1499 ( .A(ram[576]), .B(n10784), .Y(n11709) );
  INVX1 U1500 ( .A(n11709), .Y(n878) );
  AND2X1 U1501 ( .A(ram[564]), .B(n10782), .Y(n11695) );
  INVX1 U1502 ( .A(n11695), .Y(n879) );
  AND2X1 U1503 ( .A(ram[551]), .B(n10782), .Y(n11682) );
  INVX1 U1504 ( .A(n11682), .Y(n880) );
  AND2X1 U1505 ( .A(ram[538]), .B(n10782), .Y(n11669) );
  INVX1 U1506 ( .A(n11669), .Y(n881) );
  AND2X1 U1507 ( .A(ram[525]), .B(n10782), .Y(n11656) );
  INVX1 U1508 ( .A(n11656), .Y(n882) );
  AND2X1 U1509 ( .A(ram[513]), .B(n10782), .Y(n11644) );
  INVX1 U1510 ( .A(n11644), .Y(n883) );
  AND2X1 U1511 ( .A(ram[383]), .B(n10776), .Y(n11507) );
  INVX1 U1512 ( .A(n11507), .Y(n884) );
  AND2X1 U1513 ( .A(ram[370]), .B(n10776), .Y(n11494) );
  INVX1 U1514 ( .A(n11494), .Y(n885) );
  AND2X1 U1515 ( .A(ram[357]), .B(n10776), .Y(n11481) );
  INVX1 U1516 ( .A(n11481), .Y(n886) );
  AND2X1 U1517 ( .A(ram[344]), .B(n10776), .Y(n11468) );
  INVX1 U1518 ( .A(n11468), .Y(n887) );
  AND2X1 U1519 ( .A(ram[253]), .B(n10772), .Y(n11373) );
  INVX1 U1520 ( .A(n11373), .Y(n888) );
  AND2X1 U1521 ( .A(ram[240]), .B(n10772), .Y(n11360) );
  INVX1 U1522 ( .A(n11360), .Y(n889) );
  AND2X1 U1523 ( .A(ram[227]), .B(n10772), .Y(n11347) );
  INVX1 U1524 ( .A(n11347), .Y(n890) );
  AND2X1 U1525 ( .A(ram[214]), .B(n10772), .Y(n11334) );
  INVX1 U1526 ( .A(n11334), .Y(n891) );
  AND2X1 U1527 ( .A(ram[202]), .B(n10772), .Y(n11322) );
  INVX1 U1528 ( .A(n11322), .Y(n892) );
  AND2X1 U1529 ( .A(ram[190]), .B(n10770), .Y(n11308) );
  INVX1 U1530 ( .A(n11308), .Y(n893) );
  AND2X1 U1531 ( .A(ram[177]), .B(n10770), .Y(n11295) );
  INVX1 U1532 ( .A(n11295), .Y(n894) );
  AND2X1 U1533 ( .A(ram[164]), .B(n10770), .Y(n11282) );
  INVX1 U1534 ( .A(n11282), .Y(n895) );
  AND2X1 U1535 ( .A(ram[151]), .B(n10770), .Y(n11269) );
  INVX1 U1536 ( .A(n11269), .Y(n896) );
  AND2X1 U1537 ( .A(ram[139]), .B(n10770), .Y(n11257) );
  INVX1 U1538 ( .A(n11257), .Y(n897) );
  AND2X1 U1539 ( .A(ram[123]), .B(n10768), .Y(n11239) );
  INVX1 U1540 ( .A(n11239), .Y(n898) );
  AND2X1 U1541 ( .A(ram[110]), .B(n10768), .Y(n11226) );
  INVX1 U1542 ( .A(n11226), .Y(n899) );
  AND2X1 U1543 ( .A(ram[97]), .B(n10768), .Y(n11213) );
  INVX1 U1544 ( .A(n11213), .Y(n900) );
  AND2X1 U1545 ( .A(ram[84]), .B(n10768), .Y(n11200) );
  INVX1 U1546 ( .A(n11200), .Y(n901) );
  AND2X1 U1547 ( .A(ram[72]), .B(n10768), .Y(n11188) );
  INVX1 U1548 ( .A(n11188), .Y(n902) );
  AND2X1 U1549 ( .A(ram[60]), .B(n10766), .Y(n11174) );
  INVX1 U1550 ( .A(n11174), .Y(n903) );
  AND2X1 U1551 ( .A(ram[47]), .B(n10766), .Y(n11161) );
  INVX1 U1552 ( .A(n11161), .Y(n904) );
  AND2X1 U1553 ( .A(ram[34]), .B(n10766), .Y(n11148) );
  INVX1 U1554 ( .A(n11148), .Y(n905) );
  AND2X1 U1555 ( .A(ram[21]), .B(n10766), .Y(n11135) );
  INVX1 U1556 ( .A(n11135), .Y(n906) );
  AND2X1 U1557 ( .A(ram[9]), .B(n10766), .Y(n11123) );
  INVX1 U1558 ( .A(n11123), .Y(n907) );
  AND2X1 U1559 ( .A(n11112), .B(n13030), .Y(n13095) );
  AND2X1 U1560 ( .A(n11112), .B(n11576), .Y(n11641) );
  AND2X1 U1561 ( .A(n11112), .B(n11443), .Y(n11508) );
  AND2X1 U1562 ( .A(ram[1855]), .B(n10822), .Y(n13028) );
  INVX1 U1563 ( .A(n13028), .Y(n908) );
  AND2X1 U1564 ( .A(ram[1842]), .B(n10822), .Y(n13015) );
  INVX1 U1565 ( .A(n13015), .Y(n909) );
  AND2X1 U1566 ( .A(ram[1829]), .B(n10822), .Y(n13002) );
  INVX1 U1567 ( .A(n13002), .Y(n910) );
  AND2X1 U1568 ( .A(ram[1816]), .B(n10822), .Y(n12989) );
  INVX1 U1569 ( .A(n12989), .Y(n911) );
  AND2X1 U1570 ( .A(ram[1790]), .B(n10820), .Y(n12961) );
  INVX1 U1571 ( .A(n12961), .Y(n912) );
  AND2X1 U1572 ( .A(ram[1777]), .B(n10820), .Y(n12948) );
  INVX1 U1573 ( .A(n12948), .Y(n913) );
  AND2X1 U1574 ( .A(ram[1764]), .B(n10820), .Y(n12935) );
  INVX1 U1575 ( .A(n12935), .Y(n914) );
  AND2X1 U1576 ( .A(ram[1751]), .B(n10820), .Y(n12922) );
  INVX1 U1577 ( .A(n12922), .Y(n915) );
  AND2X1 U1578 ( .A(ram[1739]), .B(n10820), .Y(n12910) );
  INVX1 U1579 ( .A(n12910), .Y(n916) );
  AND2X1 U1580 ( .A(ram[1725]), .B(n10818), .Y(n12894) );
  INVX1 U1581 ( .A(n12894), .Y(n917) );
  AND2X1 U1582 ( .A(ram[1712]), .B(n10818), .Y(n12881) );
  INVX1 U1583 ( .A(n12881), .Y(n918) );
  AND2X1 U1584 ( .A(ram[1699]), .B(n10818), .Y(n12868) );
  INVX1 U1585 ( .A(n12868), .Y(n919) );
  AND2X1 U1586 ( .A(ram[1686]), .B(n10818), .Y(n12855) );
  INVX1 U1587 ( .A(n12855), .Y(n920) );
  AND2X1 U1588 ( .A(ram[1674]), .B(n10818), .Y(n12843) );
  INVX1 U1589 ( .A(n12843), .Y(n921) );
  AND2X1 U1590 ( .A(ram[1660]), .B(n10816), .Y(n12827) );
  INVX1 U1591 ( .A(n12827), .Y(n922) );
  AND2X1 U1592 ( .A(ram[1647]), .B(n10816), .Y(n12814) );
  INVX1 U1593 ( .A(n12814), .Y(n923) );
  AND2X1 U1594 ( .A(ram[1634]), .B(n10816), .Y(n12801) );
  INVX1 U1595 ( .A(n12801), .Y(n924) );
  AND2X1 U1596 ( .A(ram[1621]), .B(n10816), .Y(n12788) );
  INVX1 U1597 ( .A(n12788), .Y(n925) );
  AND2X1 U1598 ( .A(ram[1609]), .B(n10816), .Y(n12776) );
  INVX1 U1599 ( .A(n12776), .Y(n926) );
  AND2X1 U1600 ( .A(ram[1595]), .B(n10814), .Y(n12760) );
  INVX1 U1601 ( .A(n12760), .Y(n927) );
  AND2X1 U1602 ( .A(ram[1582]), .B(n10814), .Y(n12747) );
  INVX1 U1603 ( .A(n12747), .Y(n928) );
  AND2X1 U1604 ( .A(ram[1569]), .B(n10814), .Y(n12734) );
  INVX1 U1605 ( .A(n12734), .Y(n929) );
  AND2X1 U1606 ( .A(ram[1556]), .B(n10814), .Y(n12721) );
  INVX1 U1607 ( .A(n12721), .Y(n930) );
  AND2X1 U1608 ( .A(ram[1544]), .B(n10814), .Y(n12709) );
  INVX1 U1609 ( .A(n12709), .Y(n931) );
  AND2X1 U1610 ( .A(ram[1526]), .B(n10812), .Y(n12689) );
  INVX1 U1611 ( .A(n12689), .Y(n932) );
  AND2X1 U1612 ( .A(ram[1513]), .B(n10812), .Y(n12676) );
  INVX1 U1613 ( .A(n12676), .Y(n933) );
  AND2X1 U1614 ( .A(ram[1500]), .B(n10812), .Y(n12663) );
  INVX1 U1615 ( .A(n12663), .Y(n934) );
  AND2X1 U1616 ( .A(ram[1487]), .B(n10812), .Y(n12650) );
  INVX1 U1617 ( .A(n12650), .Y(n935) );
  AND2X1 U1618 ( .A(ram[1475]), .B(n10812), .Y(n12638) );
  INVX1 U1619 ( .A(n12638), .Y(n936) );
  AND2X1 U1620 ( .A(ram[1461]), .B(n10810), .Y(n12621) );
  INVX1 U1621 ( .A(n12621), .Y(n937) );
  AND2X1 U1622 ( .A(ram[1448]), .B(n10810), .Y(n12608) );
  INVX1 U1623 ( .A(n12608), .Y(n938) );
  AND2X1 U1624 ( .A(ram[1435]), .B(n10810), .Y(n12595) );
  INVX1 U1625 ( .A(n12595), .Y(n939) );
  AND2X1 U1626 ( .A(ram[1422]), .B(n10810), .Y(n12582) );
  INVX1 U1627 ( .A(n12582), .Y(n940) );
  AND2X1 U1628 ( .A(ram[1410]), .B(n10810), .Y(n12570) );
  INVX1 U1629 ( .A(n12570), .Y(n941) );
  AND2X1 U1630 ( .A(ram[1396]), .B(n10808), .Y(n12554) );
  INVX1 U1631 ( .A(n12554), .Y(n942) );
  AND2X1 U1632 ( .A(ram[1383]), .B(n10808), .Y(n12541) );
  INVX1 U1633 ( .A(n12541), .Y(n943) );
  AND2X1 U1634 ( .A(ram[1370]), .B(n10808), .Y(n12528) );
  INVX1 U1635 ( .A(n12528), .Y(n944) );
  AND2X1 U1636 ( .A(ram[1357]), .B(n10808), .Y(n12515) );
  INVX1 U1637 ( .A(n12515), .Y(n945) );
  AND2X1 U1638 ( .A(ram[1345]), .B(n10808), .Y(n12503) );
  INVX1 U1639 ( .A(n12503), .Y(n946) );
  AND2X1 U1640 ( .A(ram[1331]), .B(n10806), .Y(n12487) );
  INVX1 U1641 ( .A(n12487), .Y(n947) );
  AND2X1 U1642 ( .A(ram[1318]), .B(n10806), .Y(n12474) );
  INVX1 U1643 ( .A(n12474), .Y(n948) );
  AND2X1 U1644 ( .A(ram[1305]), .B(n10806), .Y(n12461) );
  INVX1 U1645 ( .A(n12461), .Y(n949) );
  AND2X1 U1646 ( .A(ram[1292]), .B(n10806), .Y(n12448) );
  INVX1 U1647 ( .A(n12448), .Y(n950) );
  AND2X1 U1648 ( .A(ram[1280]), .B(n10806), .Y(n12436) );
  INVX1 U1649 ( .A(n12436), .Y(n951) );
  AND2X1 U1650 ( .A(ram[1087]), .B(n10798), .Y(n12235) );
  INVX1 U1651 ( .A(n12235), .Y(n952) );
  AND2X1 U1652 ( .A(ram[1074]), .B(n10798), .Y(n12222) );
  INVX1 U1653 ( .A(n12222), .Y(n953) );
  AND2X1 U1654 ( .A(ram[1061]), .B(n10798), .Y(n12209) );
  INVX1 U1655 ( .A(n12209), .Y(n954) );
  AND2X1 U1656 ( .A(ram[1048]), .B(n10798), .Y(n12196) );
  INVX1 U1657 ( .A(n12196), .Y(n955) );
  AND2X1 U1658 ( .A(ram[1022]), .B(n10796), .Y(n12168) );
  INVX1 U1659 ( .A(n12168), .Y(n956) );
  AND2X1 U1660 ( .A(ram[1009]), .B(n10796), .Y(n12155) );
  INVX1 U1661 ( .A(n12155), .Y(n957) );
  AND2X1 U1662 ( .A(ram[996]), .B(n10796), .Y(n12142) );
  INVX1 U1663 ( .A(n12142), .Y(n958) );
  AND2X1 U1664 ( .A(ram[983]), .B(n10796), .Y(n12129) );
  INVX1 U1665 ( .A(n12129), .Y(n959) );
  AND2X1 U1666 ( .A(ram[971]), .B(n10796), .Y(n12117) );
  INVX1 U1667 ( .A(n12117), .Y(n960) );
  AND2X1 U1668 ( .A(ram[957]), .B(n10794), .Y(n12100) );
  INVX1 U1669 ( .A(n12100), .Y(n961) );
  AND2X1 U1670 ( .A(ram[944]), .B(n10794), .Y(n12087) );
  INVX1 U1671 ( .A(n12087), .Y(n962) );
  AND2X1 U1672 ( .A(ram[931]), .B(n10794), .Y(n12074) );
  INVX1 U1673 ( .A(n12074), .Y(n963) );
  AND2X1 U1674 ( .A(ram[918]), .B(n10794), .Y(n12061) );
  INVX1 U1675 ( .A(n12061), .Y(n964) );
  AND2X1 U1676 ( .A(ram[906]), .B(n10794), .Y(n12049) );
  INVX1 U1677 ( .A(n12049), .Y(n965) );
  AND2X1 U1678 ( .A(ram[892]), .B(n10792), .Y(n12033) );
  INVX1 U1679 ( .A(n12033), .Y(n966) );
  AND2X1 U1680 ( .A(ram[879]), .B(n10792), .Y(n12020) );
  INVX1 U1681 ( .A(n12020), .Y(n967) );
  AND2X1 U1682 ( .A(ram[866]), .B(n10792), .Y(n12007) );
  INVX1 U1683 ( .A(n12007), .Y(n968) );
  AND2X1 U1684 ( .A(ram[853]), .B(n10792), .Y(n11994) );
  INVX1 U1685 ( .A(n11994), .Y(n969) );
  AND2X1 U1686 ( .A(ram[841]), .B(n10792), .Y(n11982) );
  INVX1 U1687 ( .A(n11982), .Y(n970) );
  AND2X1 U1688 ( .A(ram[827]), .B(n10790), .Y(n11966) );
  INVX1 U1689 ( .A(n11966), .Y(n971) );
  AND2X1 U1690 ( .A(ram[814]), .B(n10790), .Y(n11953) );
  INVX1 U1691 ( .A(n11953), .Y(n972) );
  AND2X1 U1692 ( .A(ram[801]), .B(n10790), .Y(n11940) );
  INVX1 U1693 ( .A(n11940), .Y(n973) );
  AND2X1 U1694 ( .A(ram[788]), .B(n10790), .Y(n11927) );
  INVX1 U1695 ( .A(n11927), .Y(n974) );
  AND2X1 U1696 ( .A(ram[776]), .B(n10790), .Y(n11915) );
  INVX1 U1697 ( .A(n11915), .Y(n975) );
  AND2X1 U1698 ( .A(ram[758]), .B(n10788), .Y(n11895) );
  INVX1 U1699 ( .A(n11895), .Y(n976) );
  AND2X1 U1700 ( .A(ram[745]), .B(n10788), .Y(n11882) );
  INVX1 U1701 ( .A(n11882), .Y(n977) );
  AND2X1 U1702 ( .A(ram[732]), .B(n10788), .Y(n11869) );
  INVX1 U1703 ( .A(n11869), .Y(n978) );
  AND2X1 U1704 ( .A(ram[719]), .B(n10788), .Y(n11856) );
  INVX1 U1705 ( .A(n11856), .Y(n979) );
  AND2X1 U1706 ( .A(ram[707]), .B(n10788), .Y(n11844) );
  INVX1 U1707 ( .A(n11844), .Y(n980) );
  AND2X1 U1708 ( .A(ram[693]), .B(n10786), .Y(n11828) );
  INVX1 U1709 ( .A(n11828), .Y(n981) );
  AND2X1 U1710 ( .A(ram[680]), .B(n10786), .Y(n11815) );
  INVX1 U1711 ( .A(n11815), .Y(n982) );
  AND2X1 U1712 ( .A(ram[667]), .B(n10786), .Y(n11802) );
  INVX1 U1713 ( .A(n11802), .Y(n983) );
  AND2X1 U1714 ( .A(ram[654]), .B(n10786), .Y(n11789) );
  INVX1 U1715 ( .A(n11789), .Y(n984) );
  AND2X1 U1716 ( .A(ram[642]), .B(n10786), .Y(n11777) );
  INVX1 U1717 ( .A(n11777), .Y(n985) );
  AND2X1 U1718 ( .A(ram[628]), .B(n10784), .Y(n11761) );
  INVX1 U1719 ( .A(n11761), .Y(n986) );
  AND2X1 U1720 ( .A(ram[615]), .B(n10784), .Y(n11748) );
  INVX1 U1721 ( .A(n11748), .Y(n987) );
  AND2X1 U1722 ( .A(ram[602]), .B(n10784), .Y(n11735) );
  INVX1 U1723 ( .A(n11735), .Y(n988) );
  AND2X1 U1724 ( .A(ram[589]), .B(n10784), .Y(n11722) );
  INVX1 U1725 ( .A(n11722), .Y(n989) );
  AND2X1 U1726 ( .A(ram[577]), .B(n10784), .Y(n11710) );
  INVX1 U1727 ( .A(n11710), .Y(n990) );
  AND2X1 U1728 ( .A(ram[563]), .B(n10782), .Y(n11694) );
  INVX1 U1729 ( .A(n11694), .Y(n991) );
  AND2X1 U1730 ( .A(ram[550]), .B(n10782), .Y(n11681) );
  INVX1 U1731 ( .A(n11681), .Y(n992) );
  AND2X1 U1732 ( .A(ram[537]), .B(n10782), .Y(n11668) );
  INVX1 U1733 ( .A(n11668), .Y(n993) );
  AND2X1 U1734 ( .A(ram[524]), .B(n10782), .Y(n11655) );
  INVX1 U1735 ( .A(n11655), .Y(n994) );
  AND2X1 U1736 ( .A(ram[512]), .B(n10782), .Y(n11643) );
  INVX1 U1737 ( .A(n11643), .Y(n995) );
  AND2X1 U1738 ( .A(ram[319]), .B(n10774), .Y(n11441) );
  INVX1 U1739 ( .A(n11441), .Y(n996) );
  AND2X1 U1740 ( .A(ram[306]), .B(n10774), .Y(n11428) );
  INVX1 U1741 ( .A(n11428), .Y(n997) );
  AND2X1 U1742 ( .A(ram[293]), .B(n10774), .Y(n11415) );
  INVX1 U1743 ( .A(n11415), .Y(n998) );
  AND2X1 U1744 ( .A(ram[280]), .B(n10774), .Y(n11402) );
  INVX1 U1745 ( .A(n11402), .Y(n999) );
  AND2X1 U1746 ( .A(ram[254]), .B(n10772), .Y(n11374) );
  INVX1 U1747 ( .A(n11374), .Y(n1000) );
  AND2X1 U1748 ( .A(ram[241]), .B(n10772), .Y(n11361) );
  INVX1 U1749 ( .A(n11361), .Y(n1001) );
  AND2X1 U1750 ( .A(ram[228]), .B(n10772), .Y(n11348) );
  INVX1 U1751 ( .A(n11348), .Y(n1002) );
  AND2X1 U1752 ( .A(ram[215]), .B(n10772), .Y(n11335) );
  INVX1 U1753 ( .A(n11335), .Y(n1003) );
  AND2X1 U1754 ( .A(ram[203]), .B(n10772), .Y(n11323) );
  INVX1 U1755 ( .A(n11323), .Y(n1004) );
  AND2X1 U1756 ( .A(ram[189]), .B(n10770), .Y(n11307) );
  INVX1 U1757 ( .A(n11307), .Y(n1005) );
  AND2X1 U1758 ( .A(ram[176]), .B(n10770), .Y(n11294) );
  INVX1 U1759 ( .A(n11294), .Y(n1006) );
  AND2X1 U1760 ( .A(ram[163]), .B(n10770), .Y(n11281) );
  INVX1 U1761 ( .A(n11281), .Y(n1007) );
  AND2X1 U1762 ( .A(ram[150]), .B(n10770), .Y(n11268) );
  INVX1 U1763 ( .A(n11268), .Y(n1008) );
  AND2X1 U1764 ( .A(ram[138]), .B(n10770), .Y(n11256) );
  INVX1 U1765 ( .A(n11256), .Y(n1009) );
  AND2X1 U1766 ( .A(ram[124]), .B(n10768), .Y(n11240) );
  INVX1 U1767 ( .A(n11240), .Y(n1010) );
  AND2X1 U1768 ( .A(ram[111]), .B(n10768), .Y(n11227) );
  INVX1 U1769 ( .A(n11227), .Y(n1011) );
  AND2X1 U1770 ( .A(ram[98]), .B(n10768), .Y(n11214) );
  INVX1 U1771 ( .A(n11214), .Y(n1012) );
  AND2X1 U1772 ( .A(ram[85]), .B(n10768), .Y(n11201) );
  INVX1 U1773 ( .A(n11201), .Y(n1013) );
  AND2X1 U1774 ( .A(ram[73]), .B(n10768), .Y(n11189) );
  INVX1 U1775 ( .A(n11189), .Y(n1014) );
  AND2X1 U1776 ( .A(ram[59]), .B(n10766), .Y(n11173) );
  INVX1 U1777 ( .A(n11173), .Y(n1015) );
  AND2X1 U1778 ( .A(ram[46]), .B(n10766), .Y(n11160) );
  INVX1 U1779 ( .A(n11160), .Y(n1016) );
  AND2X1 U1780 ( .A(ram[33]), .B(n10766), .Y(n11147) );
  INVX1 U1781 ( .A(n11147), .Y(n1017) );
  AND2X1 U1782 ( .A(ram[20]), .B(n10766), .Y(n11134) );
  INVX1 U1783 ( .A(n11134), .Y(n1018) );
  AND2X1 U1784 ( .A(ram[8]), .B(n10766), .Y(n11122) );
  INVX1 U1785 ( .A(n11122), .Y(n1019) );
  AND2X1 U1786 ( .A(n11112), .B(n12501), .Y(n12566) );
  AND2X1 U1787 ( .A(n11112), .B(n11774), .Y(n11839) );
  AND2X1 U1788 ( .A(ram[1972]), .B(n10952), .Y(n13202) );
  INVX1 U1789 ( .A(n13202), .Y(n1020) );
  AND2X1 U1790 ( .A(ram[1959]), .B(n10952), .Y(n13176) );
  INVX1 U1791 ( .A(n13176), .Y(n1021) );
  AND2X1 U1792 ( .A(ram[1946]), .B(n10952), .Y(n13150) );
  INVX1 U1793 ( .A(n13150), .Y(n1022) );
  AND2X1 U1794 ( .A(ram[1933]), .B(n10952), .Y(n13124) );
  INVX1 U1795 ( .A(n13124), .Y(n1023) );
  AND2X1 U1796 ( .A(ram[1921]), .B(n10952), .Y(n13100) );
  INVX1 U1797 ( .A(n13100), .Y(n1024) );
  AND2X1 U1798 ( .A(ram[1909]), .B(n10824), .Y(n13084) );
  INVX1 U1799 ( .A(n13084), .Y(n1025) );
  AND2X1 U1800 ( .A(ram[1896]), .B(n10824), .Y(n13071) );
  INVX1 U1801 ( .A(n13071), .Y(n1026) );
  AND2X1 U1802 ( .A(ram[1883]), .B(n10824), .Y(n13058) );
  INVX1 U1803 ( .A(n13058), .Y(n1027) );
  AND2X1 U1804 ( .A(ram[1870]), .B(n10824), .Y(n13045) );
  INVX1 U1805 ( .A(n13045), .Y(n1028) );
  AND2X1 U1806 ( .A(ram[1858]), .B(n10824), .Y(n13033) );
  INVX1 U1807 ( .A(n13033), .Y(n1029) );
  AND2X1 U1808 ( .A(ram[1846]), .B(n10822), .Y(n13019) );
  INVX1 U1809 ( .A(n13019), .Y(n1030) );
  AND2X1 U1810 ( .A(ram[1833]), .B(n10822), .Y(n13006) );
  INVX1 U1811 ( .A(n13006), .Y(n1031) );
  AND2X1 U1812 ( .A(ram[1820]), .B(n10822), .Y(n12993) );
  INVX1 U1813 ( .A(n12993), .Y(n1032) );
  AND2X1 U1814 ( .A(ram[1807]), .B(n10822), .Y(n12980) );
  INVX1 U1815 ( .A(n12980), .Y(n1033) );
  AND2X1 U1816 ( .A(ram[1795]), .B(n10822), .Y(n12968) );
  INVX1 U1817 ( .A(n12968), .Y(n1034) );
  AND2X1 U1818 ( .A(ram[1783]), .B(n10820), .Y(n12954) );
  INVX1 U1819 ( .A(n12954), .Y(n1035) );
  AND2X1 U1820 ( .A(ram[1770]), .B(n10820), .Y(n12941) );
  INVX1 U1821 ( .A(n12941), .Y(n1036) );
  AND2X1 U1822 ( .A(ram[1757]), .B(n10820), .Y(n12928) );
  INVX1 U1823 ( .A(n12928), .Y(n1037) );
  AND2X1 U1824 ( .A(ram[1744]), .B(n10820), .Y(n12915) );
  INVX1 U1825 ( .A(n12915), .Y(n1038) );
  AND2X1 U1826 ( .A(ram[1732]), .B(n10820), .Y(n12903) );
  INVX1 U1827 ( .A(n12903), .Y(n1039) );
  AND2X1 U1828 ( .A(ram[1720]), .B(n10818), .Y(n12889) );
  INVX1 U1829 ( .A(n12889), .Y(n1040) );
  AND2X1 U1830 ( .A(ram[1707]), .B(n10818), .Y(n12876) );
  INVX1 U1831 ( .A(n12876), .Y(n1041) );
  AND2X1 U1832 ( .A(ram[1694]), .B(n10818), .Y(n12863) );
  INVX1 U1833 ( .A(n12863), .Y(n1042) );
  AND2X1 U1834 ( .A(ram[1681]), .B(n10818), .Y(n12850) );
  INVX1 U1835 ( .A(n12850), .Y(n1043) );
  AND2X1 U1836 ( .A(ram[1669]), .B(n10818), .Y(n12838) );
  INVX1 U1837 ( .A(n12838), .Y(n1044) );
  AND2X1 U1838 ( .A(ram[1657]), .B(n10816), .Y(n12824) );
  INVX1 U1839 ( .A(n12824), .Y(n1045) );
  AND2X1 U1840 ( .A(ram[1644]), .B(n10816), .Y(n12811) );
  INVX1 U1841 ( .A(n12811), .Y(n1046) );
  AND2X1 U1842 ( .A(ram[1631]), .B(n10816), .Y(n12798) );
  INVX1 U1843 ( .A(n12798), .Y(n1047) );
  AND2X1 U1844 ( .A(ram[1618]), .B(n10816), .Y(n12785) );
  INVX1 U1845 ( .A(n12785), .Y(n1048) );
  AND2X1 U1846 ( .A(ram[1606]), .B(n10816), .Y(n12773) );
  INVX1 U1847 ( .A(n12773), .Y(n1049) );
  AND2X1 U1848 ( .A(ram[1594]), .B(n10814), .Y(n12759) );
  INVX1 U1849 ( .A(n12759), .Y(n1050) );
  AND2X1 U1850 ( .A(ram[1581]), .B(n10814), .Y(n12746) );
  INVX1 U1851 ( .A(n12746), .Y(n1051) );
  AND2X1 U1852 ( .A(ram[1568]), .B(n10814), .Y(n12733) );
  INVX1 U1853 ( .A(n12733), .Y(n1052) );
  AND2X1 U1854 ( .A(ram[1555]), .B(n10814), .Y(n12720) );
  INVX1 U1855 ( .A(n12720), .Y(n1053) );
  AND2X1 U1856 ( .A(ram[1543]), .B(n10814), .Y(n12708) );
  INVX1 U1857 ( .A(n12708), .Y(n1054) );
  AND2X1 U1858 ( .A(ram[1535]), .B(n10812), .Y(n12698) );
  INVX1 U1859 ( .A(n12698), .Y(n1055) );
  AND2X1 U1860 ( .A(ram[1522]), .B(n10812), .Y(n12685) );
  INVX1 U1861 ( .A(n12685), .Y(n1056) );
  AND2X1 U1862 ( .A(ram[1509]), .B(n10812), .Y(n12672) );
  INVX1 U1863 ( .A(n12672), .Y(n1057) );
  AND2X1 U1864 ( .A(ram[1496]), .B(n10812), .Y(n12659) );
  INVX1 U1865 ( .A(n12659), .Y(n1058) );
  AND2X1 U1866 ( .A(ram[1267]), .B(n10804), .Y(n12421) );
  INVX1 U1867 ( .A(n12421), .Y(n1059) );
  AND2X1 U1868 ( .A(ram[1254]), .B(n10804), .Y(n12408) );
  INVX1 U1869 ( .A(n12408), .Y(n1060) );
  AND2X1 U1870 ( .A(ram[1241]), .B(n10804), .Y(n12395) );
  INVX1 U1871 ( .A(n12395), .Y(n1061) );
  AND2X1 U1872 ( .A(ram[1228]), .B(n10804), .Y(n12382) );
  INVX1 U1873 ( .A(n12382), .Y(n1062) );
  AND2X1 U1874 ( .A(ram[1216]), .B(n10804), .Y(n12370) );
  INVX1 U1875 ( .A(n12370), .Y(n1063) );
  AND2X1 U1876 ( .A(ram[1204]), .B(n10802), .Y(n12356) );
  INVX1 U1877 ( .A(n12356), .Y(n1064) );
  AND2X1 U1878 ( .A(ram[1191]), .B(n10802), .Y(n12343) );
  INVX1 U1879 ( .A(n12343), .Y(n1065) );
  AND2X1 U1880 ( .A(ram[1178]), .B(n10802), .Y(n12330) );
  INVX1 U1881 ( .A(n12330), .Y(n1066) );
  AND2X1 U1882 ( .A(ram[1165]), .B(n10802), .Y(n12317) );
  INVX1 U1883 ( .A(n12317), .Y(n1067) );
  AND2X1 U1884 ( .A(ram[1153]), .B(n10802), .Y(n12305) );
  INVX1 U1885 ( .A(n12305), .Y(n1068) );
  AND2X1 U1886 ( .A(ram[1141]), .B(n10800), .Y(n12291) );
  INVX1 U1887 ( .A(n12291), .Y(n1069) );
  AND2X1 U1888 ( .A(ram[1128]), .B(n10800), .Y(n12278) );
  INVX1 U1889 ( .A(n12278), .Y(n1070) );
  AND2X1 U1890 ( .A(ram[1115]), .B(n10800), .Y(n12265) );
  INVX1 U1891 ( .A(n12265), .Y(n1071) );
  AND2X1 U1892 ( .A(ram[1102]), .B(n10800), .Y(n12252) );
  INVX1 U1893 ( .A(n12252), .Y(n1072) );
  AND2X1 U1894 ( .A(ram[1090]), .B(n10800), .Y(n12240) );
  INVX1 U1895 ( .A(n12240), .Y(n1073) );
  AND2X1 U1896 ( .A(ram[1078]), .B(n10798), .Y(n12226) );
  INVX1 U1897 ( .A(n12226), .Y(n1074) );
  AND2X1 U1898 ( .A(ram[1065]), .B(n10798), .Y(n12213) );
  INVX1 U1899 ( .A(n12213), .Y(n1075) );
  AND2X1 U1900 ( .A(ram[1052]), .B(n10798), .Y(n12200) );
  INVX1 U1901 ( .A(n12200), .Y(n1076) );
  AND2X1 U1902 ( .A(ram[1039]), .B(n10798), .Y(n12187) );
  INVX1 U1903 ( .A(n12187), .Y(n1077) );
  AND2X1 U1904 ( .A(ram[1027]), .B(n10798), .Y(n12175) );
  INVX1 U1905 ( .A(n12175), .Y(n1078) );
  AND2X1 U1906 ( .A(ram[1015]), .B(n10796), .Y(n12161) );
  INVX1 U1907 ( .A(n12161), .Y(n1079) );
  AND2X1 U1908 ( .A(ram[1002]), .B(n10796), .Y(n12148) );
  INVX1 U1909 ( .A(n12148), .Y(n1080) );
  AND2X1 U1910 ( .A(ram[989]), .B(n10796), .Y(n12135) );
  INVX1 U1911 ( .A(n12135), .Y(n1081) );
  AND2X1 U1912 ( .A(ram[976]), .B(n10796), .Y(n12122) );
  INVX1 U1913 ( .A(n12122), .Y(n1082) );
  AND2X1 U1914 ( .A(ram[964]), .B(n10796), .Y(n12110) );
  INVX1 U1915 ( .A(n12110), .Y(n1083) );
  AND2X1 U1916 ( .A(ram[952]), .B(n10794), .Y(n12095) );
  INVX1 U1917 ( .A(n12095), .Y(n1084) );
  AND2X1 U1918 ( .A(ram[939]), .B(n10794), .Y(n12082) );
  INVX1 U1919 ( .A(n12082), .Y(n1085) );
  AND2X1 U1920 ( .A(ram[926]), .B(n10794), .Y(n12069) );
  INVX1 U1921 ( .A(n12069), .Y(n1086) );
  AND2X1 U1922 ( .A(ram[913]), .B(n10794), .Y(n12056) );
  INVX1 U1923 ( .A(n12056), .Y(n1087) );
  AND2X1 U1924 ( .A(ram[901]), .B(n10794), .Y(n12044) );
  INVX1 U1925 ( .A(n12044), .Y(n1088) );
  AND2X1 U1926 ( .A(ram[889]), .B(n10792), .Y(n12030) );
  INVX1 U1927 ( .A(n12030), .Y(n1089) );
  AND2X1 U1928 ( .A(ram[876]), .B(n10792), .Y(n12017) );
  INVX1 U1929 ( .A(n12017), .Y(n1090) );
  AND2X1 U1930 ( .A(ram[863]), .B(n10792), .Y(n12004) );
  INVX1 U1931 ( .A(n12004), .Y(n1091) );
  AND2X1 U1932 ( .A(ram[850]), .B(n10792), .Y(n11991) );
  INVX1 U1933 ( .A(n11991), .Y(n1092) );
  AND2X1 U1934 ( .A(ram[838]), .B(n10792), .Y(n11979) );
  INVX1 U1935 ( .A(n11979), .Y(n1093) );
  AND2X1 U1936 ( .A(ram[826]), .B(n10790), .Y(n11965) );
  INVX1 U1937 ( .A(n11965), .Y(n1094) );
  AND2X1 U1938 ( .A(ram[813]), .B(n10790), .Y(n11952) );
  INVX1 U1939 ( .A(n11952), .Y(n1095) );
  AND2X1 U1940 ( .A(ram[800]), .B(n10790), .Y(n11939) );
  INVX1 U1941 ( .A(n11939), .Y(n1096) );
  AND2X1 U1942 ( .A(ram[787]), .B(n10790), .Y(n11926) );
  INVX1 U1943 ( .A(n11926), .Y(n1097) );
  AND2X1 U1944 ( .A(ram[775]), .B(n10790), .Y(n11914) );
  INVX1 U1945 ( .A(n11914), .Y(n1098) );
  AND2X1 U1946 ( .A(ram[767]), .B(n10788), .Y(n11904) );
  INVX1 U1947 ( .A(n11904), .Y(n1099) );
  AND2X1 U1948 ( .A(ram[754]), .B(n10788), .Y(n11891) );
  INVX1 U1949 ( .A(n11891), .Y(n1100) );
  AND2X1 U1950 ( .A(ram[741]), .B(n10788), .Y(n11878) );
  INVX1 U1951 ( .A(n11878), .Y(n1101) );
  AND2X1 U1952 ( .A(ram[728]), .B(n10788), .Y(n11865) );
  INVX1 U1953 ( .A(n11865), .Y(n1102) );
  AND2X1 U1954 ( .A(ram[499]), .B(n10780), .Y(n11628) );
  INVX1 U1955 ( .A(n11628), .Y(n1103) );
  AND2X1 U1956 ( .A(ram[486]), .B(n10780), .Y(n11615) );
  INVX1 U1957 ( .A(n11615), .Y(n1104) );
  AND2X1 U1958 ( .A(ram[473]), .B(n10780), .Y(n11602) );
  INVX1 U1959 ( .A(n11602), .Y(n1105) );
  AND2X1 U1960 ( .A(ram[460]), .B(n10780), .Y(n11589) );
  INVX1 U1961 ( .A(n11589), .Y(n1106) );
  AND2X1 U1962 ( .A(ram[448]), .B(n10780), .Y(n11577) );
  INVX1 U1963 ( .A(n11577), .Y(n1107) );
  AND2X1 U1964 ( .A(ram[436]), .B(n10778), .Y(n11562) );
  INVX1 U1965 ( .A(n11562), .Y(n1108) );
  AND2X1 U1966 ( .A(ram[423]), .B(n10778), .Y(n11549) );
  INVX1 U1967 ( .A(n11549), .Y(n1109) );
  AND2X1 U1968 ( .A(ram[410]), .B(n10778), .Y(n11536) );
  INVX1 U1969 ( .A(n11536), .Y(n1110) );
  AND2X1 U1970 ( .A(ram[397]), .B(n10778), .Y(n11523) );
  INVX1 U1971 ( .A(n11523), .Y(n1111) );
  AND2X1 U1972 ( .A(ram[385]), .B(n10778), .Y(n11511) );
  INVX1 U1973 ( .A(n11511), .Y(n1112) );
  AND2X1 U1974 ( .A(ram[373]), .B(n10776), .Y(n11497) );
  INVX1 U1975 ( .A(n11497), .Y(n1113) );
  AND2X1 U1976 ( .A(ram[360]), .B(n10776), .Y(n11484) );
  INVX1 U1977 ( .A(n11484), .Y(n1114) );
  AND2X1 U1978 ( .A(ram[347]), .B(n10776), .Y(n11471) );
  INVX1 U1979 ( .A(n11471), .Y(n1115) );
  AND2X1 U1980 ( .A(ram[334]), .B(n10776), .Y(n11458) );
  INVX1 U1981 ( .A(n11458), .Y(n1116) );
  AND2X1 U1982 ( .A(ram[322]), .B(n10776), .Y(n11446) );
  INVX1 U1983 ( .A(n11446), .Y(n1117) );
  AND2X1 U1984 ( .A(ram[310]), .B(n10774), .Y(n11432) );
  INVX1 U1985 ( .A(n11432), .Y(n1118) );
  AND2X1 U1986 ( .A(ram[297]), .B(n10774), .Y(n11419) );
  INVX1 U1987 ( .A(n11419), .Y(n1119) );
  AND2X1 U1988 ( .A(ram[284]), .B(n10774), .Y(n11406) );
  INVX1 U1989 ( .A(n11406), .Y(n1120) );
  AND2X1 U1990 ( .A(ram[271]), .B(n10774), .Y(n11393) );
  INVX1 U1991 ( .A(n11393), .Y(n1121) );
  AND2X1 U1992 ( .A(ram[259]), .B(n10774), .Y(n11381) );
  INVX1 U1993 ( .A(n11381), .Y(n1122) );
  AND2X1 U1994 ( .A(ram[247]), .B(n10772), .Y(n11367) );
  INVX1 U1995 ( .A(n11367), .Y(n1123) );
  AND2X1 U1996 ( .A(ram[234]), .B(n10772), .Y(n11354) );
  INVX1 U1997 ( .A(n11354), .Y(n1124) );
  AND2X1 U1998 ( .A(ram[221]), .B(n10772), .Y(n11341) );
  INVX1 U1999 ( .A(n11341), .Y(n1125) );
  AND2X1 U2000 ( .A(ram[208]), .B(n10772), .Y(n11328) );
  INVX1 U2001 ( .A(n11328), .Y(n1126) );
  AND2X1 U2002 ( .A(ram[196]), .B(n10772), .Y(n11316) );
  INVX1 U2003 ( .A(n11316), .Y(n1127) );
  AND2X1 U2004 ( .A(ram[184]), .B(n10770), .Y(n11302) );
  INVX1 U2005 ( .A(n11302), .Y(n1128) );
  AND2X1 U2006 ( .A(ram[171]), .B(n10770), .Y(n11289) );
  INVX1 U2007 ( .A(n11289), .Y(n1129) );
  AND2X1 U2008 ( .A(ram[158]), .B(n10770), .Y(n11276) );
  INVX1 U2009 ( .A(n11276), .Y(n1130) );
  AND2X1 U2010 ( .A(ram[145]), .B(n10770), .Y(n11263) );
  INVX1 U2011 ( .A(n11263), .Y(n1131) );
  AND2X1 U2012 ( .A(ram[133]), .B(n10770), .Y(n11251) );
  INVX1 U2013 ( .A(n11251), .Y(n1132) );
  AND2X1 U2014 ( .A(ram[121]), .B(n10768), .Y(n11237) );
  INVX1 U2015 ( .A(n11237), .Y(n1133) );
  AND2X1 U2016 ( .A(ram[108]), .B(n10768), .Y(n11224) );
  INVX1 U2017 ( .A(n11224), .Y(n1134) );
  AND2X1 U2018 ( .A(ram[95]), .B(n10768), .Y(n11211) );
  INVX1 U2019 ( .A(n11211), .Y(n1135) );
  AND2X1 U2020 ( .A(ram[82]), .B(n10768), .Y(n11198) );
  INVX1 U2021 ( .A(n11198), .Y(n1136) );
  AND2X1 U2022 ( .A(ram[70]), .B(n10768), .Y(n11186) );
  INVX1 U2023 ( .A(n11186), .Y(n1137) );
  AND2X1 U2024 ( .A(ram[58]), .B(n10766), .Y(n11172) );
  INVX1 U2025 ( .A(n11172), .Y(n1138) );
  AND2X1 U2026 ( .A(ram[45]), .B(n10766), .Y(n11159) );
  INVX1 U2027 ( .A(n11159), .Y(n1139) );
  AND2X1 U2028 ( .A(ram[32]), .B(n10766), .Y(n11146) );
  INVX1 U2029 ( .A(n11146), .Y(n1140) );
  AND2X1 U2030 ( .A(ram[19]), .B(n10766), .Y(n11133) );
  INVX1 U2031 ( .A(n11133), .Y(n1141) );
  AND2X1 U2032 ( .A(ram[7]), .B(n10766), .Y(n11121) );
  INVX1 U2033 ( .A(n11121), .Y(n1142) );
  BUFX2 U2034 ( .A(n2785), .Y(n1143) );
  BUFX2 U2035 ( .A(n2718), .Y(n1144) );
  AND2X1 U2036 ( .A(n11112), .B(n11708), .Y(n11773) );
  AND2X1 U2037 ( .A(ram[1971]), .B(n10952), .Y(n13200) );
  INVX1 U2038 ( .A(n13200), .Y(n1145) );
  AND2X1 U2039 ( .A(ram[1958]), .B(n10952), .Y(n13174) );
  INVX1 U2040 ( .A(n13174), .Y(n1146) );
  AND2X1 U2041 ( .A(ram[1945]), .B(n10952), .Y(n13148) );
  INVX1 U2042 ( .A(n13148), .Y(n1147) );
  AND2X1 U2043 ( .A(ram[1932]), .B(n10952), .Y(n13122) );
  INVX1 U2044 ( .A(n13122), .Y(n1148) );
  AND2X1 U2045 ( .A(ram[1920]), .B(n10952), .Y(n13098) );
  INVX1 U2046 ( .A(n13098), .Y(n1149) );
  AND2X1 U2047 ( .A(ram[1910]), .B(n10824), .Y(n13085) );
  INVX1 U2048 ( .A(n13085), .Y(n1150) );
  AND2X1 U2049 ( .A(ram[1897]), .B(n10824), .Y(n13072) );
  INVX1 U2050 ( .A(n13072), .Y(n1151) );
  AND2X1 U2051 ( .A(ram[1884]), .B(n10824), .Y(n13059) );
  INVX1 U2052 ( .A(n13059), .Y(n1152) );
  AND2X1 U2053 ( .A(ram[1871]), .B(n10824), .Y(n13046) );
  INVX1 U2054 ( .A(n13046), .Y(n1153) );
  AND2X1 U2055 ( .A(ram[1859]), .B(n10824), .Y(n13034) );
  INVX1 U2056 ( .A(n13034), .Y(n1154) );
  AND2X1 U2057 ( .A(ram[1845]), .B(n10822), .Y(n13018) );
  INVX1 U2058 ( .A(n13018), .Y(n1155) );
  AND2X1 U2059 ( .A(ram[1832]), .B(n10822), .Y(n13005) );
  INVX1 U2060 ( .A(n13005), .Y(n1156) );
  AND2X1 U2061 ( .A(ram[1819]), .B(n10822), .Y(n12992) );
  INVX1 U2062 ( .A(n12992), .Y(n1157) );
  AND2X1 U2063 ( .A(ram[1806]), .B(n10822), .Y(n12979) );
  INVX1 U2064 ( .A(n12979), .Y(n1158) );
  AND2X1 U2065 ( .A(ram[1794]), .B(n10822), .Y(n12967) );
  INVX1 U2066 ( .A(n12967), .Y(n1159) );
  AND2X1 U2067 ( .A(ram[1784]), .B(n10820), .Y(n12955) );
  INVX1 U2068 ( .A(n12955), .Y(n1160) );
  AND2X1 U2069 ( .A(ram[1771]), .B(n10820), .Y(n12942) );
  INVX1 U2070 ( .A(n12942), .Y(n1161) );
  AND2X1 U2071 ( .A(ram[1758]), .B(n10820), .Y(n12929) );
  INVX1 U2072 ( .A(n12929), .Y(n1162) );
  AND2X1 U2073 ( .A(ram[1745]), .B(n10820), .Y(n12916) );
  INVX1 U2074 ( .A(n12916), .Y(n1163) );
  AND2X1 U2075 ( .A(ram[1733]), .B(n10820), .Y(n12904) );
  INVX1 U2076 ( .A(n12904), .Y(n1164) );
  AND2X1 U2077 ( .A(ram[1719]), .B(n10818), .Y(n12888) );
  INVX1 U2078 ( .A(n12888), .Y(n1165) );
  AND2X1 U2079 ( .A(ram[1706]), .B(n10818), .Y(n12875) );
  INVX1 U2080 ( .A(n12875), .Y(n1166) );
  AND2X1 U2081 ( .A(ram[1693]), .B(n10818), .Y(n12862) );
  INVX1 U2082 ( .A(n12862), .Y(n1167) );
  AND2X1 U2083 ( .A(ram[1680]), .B(n10818), .Y(n12849) );
  INVX1 U2084 ( .A(n12849), .Y(n1168) );
  AND2X1 U2085 ( .A(ram[1668]), .B(n10818), .Y(n12837) );
  INVX1 U2086 ( .A(n12837), .Y(n1169) );
  AND2X1 U2087 ( .A(ram[1658]), .B(n10816), .Y(n12825) );
  INVX1 U2088 ( .A(n12825), .Y(n1170) );
  AND2X1 U2089 ( .A(ram[1645]), .B(n10816), .Y(n12812) );
  INVX1 U2090 ( .A(n12812), .Y(n1171) );
  AND2X1 U2091 ( .A(ram[1632]), .B(n10816), .Y(n12799) );
  INVX1 U2092 ( .A(n12799), .Y(n1172) );
  AND2X1 U2093 ( .A(ram[1619]), .B(n10816), .Y(n12786) );
  INVX1 U2094 ( .A(n12786), .Y(n1173) );
  AND2X1 U2095 ( .A(ram[1607]), .B(n10816), .Y(n12774) );
  INVX1 U2096 ( .A(n12774), .Y(n1174) );
  AND2X1 U2097 ( .A(ram[1593]), .B(n10814), .Y(n12758) );
  INVX1 U2098 ( .A(n12758), .Y(n1175) );
  AND2X1 U2099 ( .A(ram[1580]), .B(n10814), .Y(n12745) );
  INVX1 U2100 ( .A(n12745), .Y(n1176) );
  AND2X1 U2101 ( .A(ram[1567]), .B(n10814), .Y(n12732) );
  INVX1 U2102 ( .A(n12732), .Y(n1177) );
  AND2X1 U2103 ( .A(ram[1554]), .B(n10814), .Y(n12719) );
  INVX1 U2104 ( .A(n12719), .Y(n1178) );
  AND2X1 U2105 ( .A(ram[1542]), .B(n10814), .Y(n12707) );
  INVX1 U2106 ( .A(n12707), .Y(n1179) );
  AND2X1 U2107 ( .A(ram[1471]), .B(n10810), .Y(n12631) );
  INVX1 U2108 ( .A(n12631), .Y(n1180) );
  AND2X1 U2109 ( .A(ram[1458]), .B(n10810), .Y(n12618) );
  INVX1 U2110 ( .A(n12618), .Y(n1181) );
  AND2X1 U2111 ( .A(ram[1445]), .B(n10810), .Y(n12605) );
  INVX1 U2112 ( .A(n12605), .Y(n1182) );
  AND2X1 U2113 ( .A(ram[1432]), .B(n10810), .Y(n12592) );
  INVX1 U2114 ( .A(n12592), .Y(n1183) );
  AND2X1 U2115 ( .A(ram[1268]), .B(n10804), .Y(n12422) );
  INVX1 U2116 ( .A(n12422), .Y(n1184) );
  AND2X1 U2117 ( .A(ram[1255]), .B(n10804), .Y(n12409) );
  INVX1 U2118 ( .A(n12409), .Y(n1185) );
  AND2X1 U2119 ( .A(ram[1242]), .B(n10804), .Y(n12396) );
  INVX1 U2120 ( .A(n12396), .Y(n1186) );
  AND2X1 U2121 ( .A(ram[1229]), .B(n10804), .Y(n12383) );
  INVX1 U2122 ( .A(n12383), .Y(n1187) );
  AND2X1 U2123 ( .A(ram[1217]), .B(n10804), .Y(n12371) );
  INVX1 U2124 ( .A(n12371), .Y(n1188) );
  AND2X1 U2125 ( .A(ram[1203]), .B(n10802), .Y(n12355) );
  INVX1 U2126 ( .A(n12355), .Y(n1189) );
  AND2X1 U2127 ( .A(ram[1190]), .B(n10802), .Y(n12342) );
  INVX1 U2128 ( .A(n12342), .Y(n1190) );
  AND2X1 U2129 ( .A(ram[1177]), .B(n10802), .Y(n12329) );
  INVX1 U2130 ( .A(n12329), .Y(n1191) );
  AND2X1 U2131 ( .A(ram[1164]), .B(n10802), .Y(n12316) );
  INVX1 U2132 ( .A(n12316), .Y(n1192) );
  AND2X1 U2133 ( .A(ram[1152]), .B(n10802), .Y(n12304) );
  INVX1 U2134 ( .A(n12304), .Y(n1193) );
  AND2X1 U2135 ( .A(ram[1142]), .B(n10800), .Y(n12292) );
  INVX1 U2136 ( .A(n12292), .Y(n1194) );
  AND2X1 U2137 ( .A(ram[1129]), .B(n10800), .Y(n12279) );
  INVX1 U2138 ( .A(n12279), .Y(n1195) );
  AND2X1 U2139 ( .A(ram[1116]), .B(n10800), .Y(n12266) );
  INVX1 U2140 ( .A(n12266), .Y(n1196) );
  AND2X1 U2141 ( .A(ram[1103]), .B(n10800), .Y(n12253) );
  INVX1 U2142 ( .A(n12253), .Y(n1197) );
  AND2X1 U2143 ( .A(ram[1091]), .B(n10800), .Y(n12241) );
  INVX1 U2144 ( .A(n12241), .Y(n1198) );
  AND2X1 U2145 ( .A(ram[1077]), .B(n10798), .Y(n12225) );
  INVX1 U2146 ( .A(n12225), .Y(n1199) );
  AND2X1 U2147 ( .A(ram[1064]), .B(n10798), .Y(n12212) );
  INVX1 U2148 ( .A(n12212), .Y(n1200) );
  AND2X1 U2149 ( .A(ram[1051]), .B(n10798), .Y(n12199) );
  INVX1 U2150 ( .A(n12199), .Y(n1201) );
  AND2X1 U2151 ( .A(ram[1038]), .B(n10798), .Y(n12186) );
  INVX1 U2152 ( .A(n12186), .Y(n1202) );
  AND2X1 U2153 ( .A(ram[1026]), .B(n10798), .Y(n12174) );
  INVX1 U2154 ( .A(n12174), .Y(n1203) );
  AND2X1 U2155 ( .A(ram[1016]), .B(n10796), .Y(n12162) );
  INVX1 U2156 ( .A(n12162), .Y(n1204) );
  AND2X1 U2157 ( .A(ram[1003]), .B(n10796), .Y(n12149) );
  INVX1 U2158 ( .A(n12149), .Y(n1205) );
  AND2X1 U2159 ( .A(ram[990]), .B(n10796), .Y(n12136) );
  INVX1 U2160 ( .A(n12136), .Y(n1206) );
  AND2X1 U2161 ( .A(ram[977]), .B(n10796), .Y(n12123) );
  INVX1 U2162 ( .A(n12123), .Y(n1207) );
  AND2X1 U2163 ( .A(ram[965]), .B(n10796), .Y(n12111) );
  INVX1 U2164 ( .A(n12111), .Y(n1208) );
  AND2X1 U2165 ( .A(ram[951]), .B(n10794), .Y(n12094) );
  INVX1 U2166 ( .A(n12094), .Y(n1209) );
  AND2X1 U2167 ( .A(ram[938]), .B(n10794), .Y(n12081) );
  INVX1 U2168 ( .A(n12081), .Y(n1210) );
  AND2X1 U2169 ( .A(ram[925]), .B(n10794), .Y(n12068) );
  INVX1 U2170 ( .A(n12068), .Y(n1211) );
  AND2X1 U2171 ( .A(ram[912]), .B(n10794), .Y(n12055) );
  INVX1 U2172 ( .A(n12055), .Y(n1212) );
  AND2X1 U2173 ( .A(ram[900]), .B(n10794), .Y(n12043) );
  INVX1 U2174 ( .A(n12043), .Y(n1213) );
  AND2X1 U2175 ( .A(ram[890]), .B(n10792), .Y(n12031) );
  INVX1 U2176 ( .A(n12031), .Y(n1214) );
  AND2X1 U2177 ( .A(ram[877]), .B(n10792), .Y(n12018) );
  INVX1 U2178 ( .A(n12018), .Y(n1215) );
  AND2X1 U2179 ( .A(ram[864]), .B(n10792), .Y(n12005) );
  INVX1 U2180 ( .A(n12005), .Y(n1216) );
  AND2X1 U2181 ( .A(ram[851]), .B(n10792), .Y(n11992) );
  INVX1 U2182 ( .A(n11992), .Y(n1217) );
  AND2X1 U2183 ( .A(ram[839]), .B(n10792), .Y(n11980) );
  INVX1 U2184 ( .A(n11980), .Y(n1218) );
  AND2X1 U2185 ( .A(ram[825]), .B(n10790), .Y(n11964) );
  INVX1 U2186 ( .A(n11964), .Y(n1219) );
  AND2X1 U2187 ( .A(ram[812]), .B(n10790), .Y(n11951) );
  INVX1 U2188 ( .A(n11951), .Y(n1220) );
  AND2X1 U2189 ( .A(ram[799]), .B(n10790), .Y(n11938) );
  INVX1 U2190 ( .A(n11938), .Y(n1221) );
  AND2X1 U2191 ( .A(ram[786]), .B(n10790), .Y(n11925) );
  INVX1 U2192 ( .A(n11925), .Y(n1222) );
  AND2X1 U2193 ( .A(ram[774]), .B(n10790), .Y(n11913) );
  INVX1 U2194 ( .A(n11913), .Y(n1223) );
  AND2X1 U2195 ( .A(ram[703]), .B(n10786), .Y(n11838) );
  INVX1 U2196 ( .A(n11838), .Y(n1224) );
  AND2X1 U2197 ( .A(ram[690]), .B(n10786), .Y(n11825) );
  INVX1 U2198 ( .A(n11825), .Y(n1225) );
  AND2X1 U2199 ( .A(ram[677]), .B(n10786), .Y(n11812) );
  INVX1 U2200 ( .A(n11812), .Y(n1226) );
  AND2X1 U2201 ( .A(ram[664]), .B(n10786), .Y(n11799) );
  INVX1 U2202 ( .A(n11799), .Y(n1227) );
  AND2X1 U2203 ( .A(ram[500]), .B(n10780), .Y(n11629) );
  INVX1 U2204 ( .A(n11629), .Y(n1228) );
  AND2X1 U2205 ( .A(ram[487]), .B(n10780), .Y(n11616) );
  INVX1 U2206 ( .A(n11616), .Y(n1229) );
  AND2X1 U2207 ( .A(ram[474]), .B(n10780), .Y(n11603) );
  INVX1 U2208 ( .A(n11603), .Y(n1230) );
  AND2X1 U2209 ( .A(ram[461]), .B(n10780), .Y(n11590) );
  INVX1 U2210 ( .A(n11590), .Y(n1231) );
  AND2X1 U2211 ( .A(ram[449]), .B(n10780), .Y(n11578) );
  INVX1 U2212 ( .A(n11578), .Y(n1232) );
  AND2X1 U2213 ( .A(ram[435]), .B(n10778), .Y(n11561) );
  INVX1 U2214 ( .A(n11561), .Y(n1233) );
  AND2X1 U2215 ( .A(ram[422]), .B(n10778), .Y(n11548) );
  INVX1 U2216 ( .A(n11548), .Y(n1234) );
  AND2X1 U2217 ( .A(ram[409]), .B(n10778), .Y(n11535) );
  INVX1 U2218 ( .A(n11535), .Y(n1235) );
  AND2X1 U2219 ( .A(ram[396]), .B(n10778), .Y(n11522) );
  INVX1 U2220 ( .A(n11522), .Y(n1236) );
  AND2X1 U2221 ( .A(ram[384]), .B(n10778), .Y(n11510) );
  INVX1 U2222 ( .A(n11510), .Y(n1237) );
  AND2X1 U2223 ( .A(ram[374]), .B(n10776), .Y(n11498) );
  INVX1 U2224 ( .A(n11498), .Y(n1238) );
  AND2X1 U2225 ( .A(ram[361]), .B(n10776), .Y(n11485) );
  INVX1 U2226 ( .A(n11485), .Y(n1239) );
  AND2X1 U2227 ( .A(ram[348]), .B(n10776), .Y(n11472) );
  INVX1 U2228 ( .A(n11472), .Y(n1240) );
  AND2X1 U2229 ( .A(ram[335]), .B(n10776), .Y(n11459) );
  INVX1 U2230 ( .A(n11459), .Y(n1241) );
  AND2X1 U2231 ( .A(ram[323]), .B(n10776), .Y(n11447) );
  INVX1 U2232 ( .A(n11447), .Y(n1242) );
  AND2X1 U2233 ( .A(ram[309]), .B(n10774), .Y(n11431) );
  INVX1 U2234 ( .A(n11431), .Y(n1243) );
  AND2X1 U2235 ( .A(ram[296]), .B(n10774), .Y(n11418) );
  INVX1 U2236 ( .A(n11418), .Y(n1244) );
  AND2X1 U2237 ( .A(ram[283]), .B(n10774), .Y(n11405) );
  INVX1 U2238 ( .A(n11405), .Y(n1245) );
  AND2X1 U2239 ( .A(ram[270]), .B(n10774), .Y(n11392) );
  INVX1 U2240 ( .A(n11392), .Y(n1246) );
  AND2X1 U2241 ( .A(ram[258]), .B(n10774), .Y(n11380) );
  INVX1 U2242 ( .A(n11380), .Y(n1247) );
  AND2X1 U2243 ( .A(ram[248]), .B(n10772), .Y(n11368) );
  INVX1 U2244 ( .A(n11368), .Y(n1248) );
  AND2X1 U2245 ( .A(ram[235]), .B(n10772), .Y(n11355) );
  INVX1 U2246 ( .A(n11355), .Y(n1249) );
  AND2X1 U2247 ( .A(ram[222]), .B(n10772), .Y(n11342) );
  INVX1 U2248 ( .A(n11342), .Y(n1250) );
  AND2X1 U2249 ( .A(ram[209]), .B(n10772), .Y(n11329) );
  INVX1 U2250 ( .A(n11329), .Y(n1251) );
  AND2X1 U2251 ( .A(ram[197]), .B(n10772), .Y(n11317) );
  INVX1 U2252 ( .A(n11317), .Y(n1252) );
  AND2X1 U2253 ( .A(ram[183]), .B(n10770), .Y(n11301) );
  INVX1 U2254 ( .A(n11301), .Y(n1253) );
  AND2X1 U2255 ( .A(ram[170]), .B(n10770), .Y(n11288) );
  INVX1 U2256 ( .A(n11288), .Y(n1254) );
  AND2X1 U2257 ( .A(ram[157]), .B(n10770), .Y(n11275) );
  INVX1 U2258 ( .A(n11275), .Y(n1255) );
  AND2X1 U2259 ( .A(ram[144]), .B(n10770), .Y(n11262) );
  INVX1 U2260 ( .A(n11262), .Y(n1256) );
  AND2X1 U2261 ( .A(ram[132]), .B(n10770), .Y(n11250) );
  INVX1 U2262 ( .A(n11250), .Y(n1257) );
  AND2X1 U2263 ( .A(ram[122]), .B(n10768), .Y(n11238) );
  INVX1 U2264 ( .A(n11238), .Y(n1258) );
  AND2X1 U2265 ( .A(ram[109]), .B(n10768), .Y(n11225) );
  INVX1 U2266 ( .A(n11225), .Y(n1259) );
  AND2X1 U2267 ( .A(ram[96]), .B(n10768), .Y(n11212) );
  INVX1 U2268 ( .A(n11212), .Y(n1260) );
  AND2X1 U2269 ( .A(ram[83]), .B(n10768), .Y(n11199) );
  INVX1 U2270 ( .A(n11199), .Y(n1261) );
  AND2X1 U2271 ( .A(ram[71]), .B(n10768), .Y(n11187) );
  INVX1 U2272 ( .A(n11187), .Y(n1262) );
  AND2X1 U2273 ( .A(ram[57]), .B(n10766), .Y(n11171) );
  INVX1 U2274 ( .A(n11171), .Y(n1263) );
  AND2X1 U2275 ( .A(ram[44]), .B(n10766), .Y(n11158) );
  INVX1 U2276 ( .A(n11158), .Y(n1264) );
  AND2X1 U2277 ( .A(ram[31]), .B(n10766), .Y(n11145) );
  INVX1 U2278 ( .A(n11145), .Y(n1265) );
  AND2X1 U2279 ( .A(ram[18]), .B(n10766), .Y(n11132) );
  INVX1 U2280 ( .A(n11132), .Y(n1266) );
  AND2X1 U2281 ( .A(ram[6]), .B(n10766), .Y(n11120) );
  INVX1 U2282 ( .A(n11120), .Y(n1267) );
  BUFX2 U2283 ( .A(n2852), .Y(n1268) );
  BUFX2 U2284 ( .A(n2651), .Y(n1269) );
  AND2X1 U2285 ( .A(n11112), .B(n12634), .Y(n12699) );
  AND2X1 U2286 ( .A(n11112), .B(n11642), .Y(n11707) );
  AND2X1 U2287 ( .A(ram[1974]), .B(n10952), .Y(n13206) );
  INVX1 U2288 ( .A(n13206), .Y(n1270) );
  AND2X1 U2289 ( .A(ram[1961]), .B(n10952), .Y(n13180) );
  INVX1 U2290 ( .A(n13180), .Y(n1271) );
  AND2X1 U2291 ( .A(ram[1948]), .B(n10952), .Y(n13154) );
  INVX1 U2292 ( .A(n13154), .Y(n1272) );
  AND2X1 U2293 ( .A(ram[1935]), .B(n10952), .Y(n13128) );
  INVX1 U2294 ( .A(n13128), .Y(n1273) );
  AND2X1 U2295 ( .A(ram[1923]), .B(n10952), .Y(n13104) );
  INVX1 U2296 ( .A(n13104), .Y(n1274) );
  AND2X1 U2297 ( .A(ram[1907]), .B(n10824), .Y(n13082) );
  INVX1 U2298 ( .A(n13082), .Y(n1275) );
  AND2X1 U2299 ( .A(ram[1894]), .B(n10824), .Y(n13069) );
  INVX1 U2300 ( .A(n13069), .Y(n1276) );
  AND2X1 U2301 ( .A(ram[1881]), .B(n10824), .Y(n13056) );
  INVX1 U2302 ( .A(n13056), .Y(n1277) );
  AND2X1 U2303 ( .A(ram[1868]), .B(n10824), .Y(n13043) );
  INVX1 U2304 ( .A(n13043), .Y(n1278) );
  AND2X1 U2305 ( .A(ram[1856]), .B(n10824), .Y(n13031) );
  INVX1 U2306 ( .A(n13031), .Y(n1279) );
  AND2X1 U2307 ( .A(ram[1844]), .B(n10822), .Y(n13017) );
  INVX1 U2308 ( .A(n13017), .Y(n1280) );
  AND2X1 U2309 ( .A(ram[1831]), .B(n10822), .Y(n13004) );
  INVX1 U2310 ( .A(n13004), .Y(n1281) );
  AND2X1 U2311 ( .A(ram[1818]), .B(n10822), .Y(n12991) );
  INVX1 U2312 ( .A(n12991), .Y(n1282) );
  AND2X1 U2313 ( .A(ram[1805]), .B(n10822), .Y(n12978) );
  INVX1 U2314 ( .A(n12978), .Y(n1283) );
  AND2X1 U2315 ( .A(ram[1793]), .B(n10822), .Y(n12966) );
  INVX1 U2316 ( .A(n12966), .Y(n1284) );
  AND2X1 U2317 ( .A(ram[1785]), .B(n10820), .Y(n12956) );
  INVX1 U2318 ( .A(n12956), .Y(n1285) );
  AND2X1 U2319 ( .A(ram[1772]), .B(n10820), .Y(n12943) );
  INVX1 U2320 ( .A(n12943), .Y(n1286) );
  AND2X1 U2321 ( .A(ram[1759]), .B(n10820), .Y(n12930) );
  INVX1 U2322 ( .A(n12930), .Y(n1287) );
  AND2X1 U2323 ( .A(ram[1746]), .B(n10820), .Y(n12917) );
  INVX1 U2324 ( .A(n12917), .Y(n1288) );
  AND2X1 U2325 ( .A(ram[1734]), .B(n10820), .Y(n12905) );
  INVX1 U2326 ( .A(n12905), .Y(n1289) );
  AND2X1 U2327 ( .A(ram[1722]), .B(n10818), .Y(n12891) );
  INVX1 U2328 ( .A(n12891), .Y(n1290) );
  AND2X1 U2329 ( .A(ram[1709]), .B(n10818), .Y(n12878) );
  INVX1 U2330 ( .A(n12878), .Y(n1291) );
  AND2X1 U2331 ( .A(ram[1696]), .B(n10818), .Y(n12865) );
  INVX1 U2332 ( .A(n12865), .Y(n1292) );
  AND2X1 U2333 ( .A(ram[1683]), .B(n10818), .Y(n12852) );
  INVX1 U2334 ( .A(n12852), .Y(n1293) );
  AND2X1 U2335 ( .A(ram[1671]), .B(n10818), .Y(n12840) );
  INVX1 U2336 ( .A(n12840), .Y(n1294) );
  AND2X1 U2337 ( .A(ram[1655]), .B(n10816), .Y(n12822) );
  INVX1 U2338 ( .A(n12822), .Y(n1295) );
  AND2X1 U2339 ( .A(ram[1642]), .B(n10816), .Y(n12809) );
  INVX1 U2340 ( .A(n12809), .Y(n1296) );
  AND2X1 U2341 ( .A(ram[1629]), .B(n10816), .Y(n12796) );
  INVX1 U2342 ( .A(n12796), .Y(n1297) );
  AND2X1 U2343 ( .A(ram[1616]), .B(n10816), .Y(n12783) );
  INVX1 U2344 ( .A(n12783), .Y(n1298) );
  AND2X1 U2345 ( .A(ram[1604]), .B(n10816), .Y(n12771) );
  INVX1 U2346 ( .A(n12771), .Y(n1299) );
  AND2X1 U2347 ( .A(ram[1592]), .B(n10814), .Y(n12757) );
  INVX1 U2348 ( .A(n12757), .Y(n1300) );
  AND2X1 U2349 ( .A(ram[1579]), .B(n10814), .Y(n12744) );
  INVX1 U2350 ( .A(n12744), .Y(n1301) );
  AND2X1 U2351 ( .A(ram[1566]), .B(n10814), .Y(n12731) );
  INVX1 U2352 ( .A(n12731), .Y(n1302) );
  AND2X1 U2353 ( .A(ram[1553]), .B(n10814), .Y(n12718) );
  INVX1 U2354 ( .A(n12718), .Y(n1303) );
  AND2X1 U2355 ( .A(ram[1541]), .B(n10814), .Y(n12706) );
  INVX1 U2356 ( .A(n12706), .Y(n1304) );
  AND2X1 U2357 ( .A(ram[1407]), .B(n10808), .Y(n12565) );
  INVX1 U2358 ( .A(n12565), .Y(n1305) );
  AND2X1 U2359 ( .A(ram[1394]), .B(n10808), .Y(n12552) );
  INVX1 U2360 ( .A(n12552), .Y(n1306) );
  AND2X1 U2361 ( .A(ram[1381]), .B(n10808), .Y(n12539) );
  INVX1 U2362 ( .A(n12539), .Y(n1307) );
  AND2X1 U2363 ( .A(ram[1368]), .B(n10808), .Y(n12526) );
  INVX1 U2364 ( .A(n12526), .Y(n1308) );
  AND2X1 U2365 ( .A(ram[1269]), .B(n10804), .Y(n12423) );
  INVX1 U2366 ( .A(n12423), .Y(n1309) );
  AND2X1 U2367 ( .A(ram[1256]), .B(n10804), .Y(n12410) );
  INVX1 U2368 ( .A(n12410), .Y(n1310) );
  AND2X1 U2369 ( .A(ram[1243]), .B(n10804), .Y(n12397) );
  INVX1 U2370 ( .A(n12397), .Y(n1311) );
  AND2X1 U2371 ( .A(ram[1230]), .B(n10804), .Y(n12384) );
  INVX1 U2372 ( .A(n12384), .Y(n1312) );
  AND2X1 U2373 ( .A(ram[1218]), .B(n10804), .Y(n12372) );
  INVX1 U2374 ( .A(n12372), .Y(n1313) );
  AND2X1 U2375 ( .A(ram[1206]), .B(n10802), .Y(n12358) );
  INVX1 U2376 ( .A(n12358), .Y(n1314) );
  AND2X1 U2377 ( .A(ram[1193]), .B(n10802), .Y(n12345) );
  INVX1 U2378 ( .A(n12345), .Y(n1315) );
  AND2X1 U2379 ( .A(ram[1180]), .B(n10802), .Y(n12332) );
  INVX1 U2380 ( .A(n12332), .Y(n1316) );
  AND2X1 U2381 ( .A(ram[1167]), .B(n10802), .Y(n12319) );
  INVX1 U2382 ( .A(n12319), .Y(n1317) );
  AND2X1 U2383 ( .A(ram[1155]), .B(n10802), .Y(n12307) );
  INVX1 U2384 ( .A(n12307), .Y(n1318) );
  AND2X1 U2385 ( .A(ram[1139]), .B(n10800), .Y(n12289) );
  INVX1 U2386 ( .A(n12289), .Y(n1319) );
  AND2X1 U2387 ( .A(ram[1126]), .B(n10800), .Y(n12276) );
  INVX1 U2388 ( .A(n12276), .Y(n1320) );
  AND2X1 U2389 ( .A(ram[1113]), .B(n10800), .Y(n12263) );
  INVX1 U2390 ( .A(n12263), .Y(n1321) );
  AND2X1 U2391 ( .A(ram[1100]), .B(n10800), .Y(n12250) );
  INVX1 U2392 ( .A(n12250), .Y(n1322) );
  AND2X1 U2393 ( .A(ram[1088]), .B(n10800), .Y(n12238) );
  INVX1 U2394 ( .A(n12238), .Y(n1323) );
  AND2X1 U2395 ( .A(ram[1076]), .B(n10798), .Y(n12224) );
  INVX1 U2396 ( .A(n12224), .Y(n1324) );
  AND2X1 U2397 ( .A(ram[1063]), .B(n10798), .Y(n12211) );
  INVX1 U2398 ( .A(n12211), .Y(n1325) );
  AND2X1 U2399 ( .A(ram[1050]), .B(n10798), .Y(n12198) );
  INVX1 U2400 ( .A(n12198), .Y(n1326) );
  AND2X1 U2401 ( .A(ram[1037]), .B(n10798), .Y(n12185) );
  INVX1 U2402 ( .A(n12185), .Y(n1327) );
  AND2X1 U2403 ( .A(ram[1025]), .B(n10798), .Y(n12173) );
  INVX1 U2404 ( .A(n12173), .Y(n1328) );
  AND2X1 U2405 ( .A(ram[1017]), .B(n10796), .Y(n12163) );
  INVX1 U2406 ( .A(n12163), .Y(n1329) );
  AND2X1 U2407 ( .A(ram[1004]), .B(n10796), .Y(n12150) );
  INVX1 U2408 ( .A(n12150), .Y(n1330) );
  AND2X1 U2409 ( .A(ram[991]), .B(n10796), .Y(n12137) );
  INVX1 U2410 ( .A(n12137), .Y(n1331) );
  AND2X1 U2411 ( .A(ram[978]), .B(n10796), .Y(n12124) );
  INVX1 U2412 ( .A(n12124), .Y(n1332) );
  AND2X1 U2413 ( .A(ram[966]), .B(n10796), .Y(n12112) );
  INVX1 U2414 ( .A(n12112), .Y(n1333) );
  AND2X1 U2415 ( .A(ram[954]), .B(n10794), .Y(n12097) );
  INVX1 U2416 ( .A(n12097), .Y(n1334) );
  AND2X1 U2417 ( .A(ram[941]), .B(n10794), .Y(n12084) );
  INVX1 U2418 ( .A(n12084), .Y(n1335) );
  AND2X1 U2419 ( .A(ram[928]), .B(n10794), .Y(n12071) );
  INVX1 U2420 ( .A(n12071), .Y(n1336) );
  AND2X1 U2421 ( .A(ram[915]), .B(n10794), .Y(n12058) );
  INVX1 U2422 ( .A(n12058), .Y(n1337) );
  AND2X1 U2423 ( .A(ram[903]), .B(n10794), .Y(n12046) );
  INVX1 U2424 ( .A(n12046), .Y(n1338) );
  AND2X1 U2425 ( .A(ram[887]), .B(n10792), .Y(n12028) );
  INVX1 U2426 ( .A(n12028), .Y(n1339) );
  AND2X1 U2427 ( .A(ram[874]), .B(n10792), .Y(n12015) );
  INVX1 U2428 ( .A(n12015), .Y(n1340) );
  AND2X1 U2429 ( .A(ram[861]), .B(n10792), .Y(n12002) );
  INVX1 U2430 ( .A(n12002), .Y(n1341) );
  AND2X1 U2431 ( .A(ram[848]), .B(n10792), .Y(n11989) );
  INVX1 U2432 ( .A(n11989), .Y(n1342) );
  AND2X1 U2433 ( .A(ram[836]), .B(n10792), .Y(n11977) );
  INVX1 U2434 ( .A(n11977), .Y(n1343) );
  AND2X1 U2435 ( .A(ram[824]), .B(n10790), .Y(n11963) );
  INVX1 U2436 ( .A(n11963), .Y(n1344) );
  AND2X1 U2437 ( .A(ram[811]), .B(n10790), .Y(n11950) );
  INVX1 U2438 ( .A(n11950), .Y(n1345) );
  AND2X1 U2439 ( .A(ram[798]), .B(n10790), .Y(n11937) );
  INVX1 U2440 ( .A(n11937), .Y(n1346) );
  AND2X1 U2441 ( .A(ram[785]), .B(n10790), .Y(n11924) );
  INVX1 U2442 ( .A(n11924), .Y(n1347) );
  AND2X1 U2443 ( .A(ram[773]), .B(n10790), .Y(n11912) );
  INVX1 U2444 ( .A(n11912), .Y(n1348) );
  AND2X1 U2445 ( .A(ram[639]), .B(n10784), .Y(n11772) );
  INVX1 U2446 ( .A(n11772), .Y(n1349) );
  AND2X1 U2447 ( .A(ram[626]), .B(n10784), .Y(n11759) );
  INVX1 U2448 ( .A(n11759), .Y(n1350) );
  AND2X1 U2449 ( .A(ram[613]), .B(n10784), .Y(n11746) );
  INVX1 U2450 ( .A(n11746), .Y(n1351) );
  AND2X1 U2451 ( .A(ram[600]), .B(n10784), .Y(n11733) );
  INVX1 U2452 ( .A(n11733), .Y(n1352) );
  AND2X1 U2453 ( .A(ram[501]), .B(n10780), .Y(n11630) );
  INVX1 U2454 ( .A(n11630), .Y(n1353) );
  AND2X1 U2455 ( .A(ram[488]), .B(n10780), .Y(n11617) );
  INVX1 U2456 ( .A(n11617), .Y(n1354) );
  AND2X1 U2457 ( .A(ram[475]), .B(n10780), .Y(n11604) );
  INVX1 U2458 ( .A(n11604), .Y(n1355) );
  AND2X1 U2459 ( .A(ram[462]), .B(n10780), .Y(n11591) );
  INVX1 U2460 ( .A(n11591), .Y(n1356) );
  AND2X1 U2461 ( .A(ram[450]), .B(n10780), .Y(n11579) );
  INVX1 U2462 ( .A(n11579), .Y(n1357) );
  AND2X1 U2463 ( .A(ram[438]), .B(n10778), .Y(n11564) );
  INVX1 U2464 ( .A(n11564), .Y(n1358) );
  AND2X1 U2465 ( .A(ram[425]), .B(n10778), .Y(n11551) );
  INVX1 U2466 ( .A(n11551), .Y(n1359) );
  AND2X1 U2467 ( .A(ram[412]), .B(n10778), .Y(n11538) );
  INVX1 U2468 ( .A(n11538), .Y(n1360) );
  AND2X1 U2469 ( .A(ram[399]), .B(n10778), .Y(n11525) );
  INVX1 U2470 ( .A(n11525), .Y(n1361) );
  AND2X1 U2471 ( .A(ram[387]), .B(n10778), .Y(n11513) );
  INVX1 U2472 ( .A(n11513), .Y(n1362) );
  AND2X1 U2473 ( .A(ram[371]), .B(n10776), .Y(n11495) );
  INVX1 U2474 ( .A(n11495), .Y(n1363) );
  AND2X1 U2475 ( .A(ram[358]), .B(n10776), .Y(n11482) );
  INVX1 U2476 ( .A(n11482), .Y(n1364) );
  AND2X1 U2477 ( .A(ram[345]), .B(n10776), .Y(n11469) );
  INVX1 U2478 ( .A(n11469), .Y(n1365) );
  AND2X1 U2479 ( .A(ram[332]), .B(n10776), .Y(n11456) );
  INVX1 U2480 ( .A(n11456), .Y(n1366) );
  AND2X1 U2481 ( .A(ram[320]), .B(n10776), .Y(n11444) );
  INVX1 U2482 ( .A(n11444), .Y(n1367) );
  AND2X1 U2483 ( .A(ram[308]), .B(n10774), .Y(n11430) );
  INVX1 U2484 ( .A(n11430), .Y(n1368) );
  AND2X1 U2485 ( .A(ram[295]), .B(n10774), .Y(n11417) );
  INVX1 U2486 ( .A(n11417), .Y(n1369) );
  AND2X1 U2487 ( .A(ram[282]), .B(n10774), .Y(n11404) );
  INVX1 U2488 ( .A(n11404), .Y(n1370) );
  AND2X1 U2489 ( .A(ram[269]), .B(n10774), .Y(n11391) );
  INVX1 U2490 ( .A(n11391), .Y(n1371) );
  AND2X1 U2491 ( .A(ram[257]), .B(n10774), .Y(n11379) );
  INVX1 U2492 ( .A(n11379), .Y(n1372) );
  AND2X1 U2493 ( .A(ram[249]), .B(n10772), .Y(n11369) );
  INVX1 U2494 ( .A(n11369), .Y(n1373) );
  AND2X1 U2495 ( .A(ram[236]), .B(n10772), .Y(n11356) );
  INVX1 U2496 ( .A(n11356), .Y(n1374) );
  AND2X1 U2497 ( .A(ram[223]), .B(n10772), .Y(n11343) );
  INVX1 U2498 ( .A(n11343), .Y(n1375) );
  AND2X1 U2499 ( .A(ram[210]), .B(n10772), .Y(n11330) );
  INVX1 U2500 ( .A(n11330), .Y(n1376) );
  AND2X1 U2501 ( .A(ram[198]), .B(n10772), .Y(n11318) );
  INVX1 U2502 ( .A(n11318), .Y(n1377) );
  AND2X1 U2503 ( .A(ram[186]), .B(n10770), .Y(n11304) );
  INVX1 U2504 ( .A(n11304), .Y(n1378) );
  AND2X1 U2505 ( .A(ram[173]), .B(n10770), .Y(n11291) );
  INVX1 U2506 ( .A(n11291), .Y(n1379) );
  AND2X1 U2507 ( .A(ram[160]), .B(n10770), .Y(n11278) );
  INVX1 U2508 ( .A(n11278), .Y(n1380) );
  AND2X1 U2509 ( .A(ram[147]), .B(n10770), .Y(n11265) );
  INVX1 U2510 ( .A(n11265), .Y(n1381) );
  AND2X1 U2511 ( .A(ram[135]), .B(n10770), .Y(n11253) );
  INVX1 U2512 ( .A(n11253), .Y(n1382) );
  AND2X1 U2513 ( .A(ram[119]), .B(n10768), .Y(n11235) );
  INVX1 U2514 ( .A(n11235), .Y(n1383) );
  AND2X1 U2515 ( .A(ram[106]), .B(n10768), .Y(n11222) );
  INVX1 U2516 ( .A(n11222), .Y(n1384) );
  AND2X1 U2517 ( .A(ram[93]), .B(n10768), .Y(n11209) );
  INVX1 U2518 ( .A(n11209), .Y(n1385) );
  AND2X1 U2519 ( .A(ram[80]), .B(n10768), .Y(n11196) );
  INVX1 U2520 ( .A(n11196), .Y(n1386) );
  AND2X1 U2521 ( .A(ram[68]), .B(n10768), .Y(n11184) );
  INVX1 U2522 ( .A(n11184), .Y(n1387) );
  AND2X1 U2523 ( .A(ram[56]), .B(n10766), .Y(n11170) );
  INVX1 U2524 ( .A(n11170), .Y(n1388) );
  AND2X1 U2525 ( .A(ram[43]), .B(n10766), .Y(n11157) );
  INVX1 U2526 ( .A(n11157), .Y(n1389) );
  AND2X1 U2527 ( .A(ram[30]), .B(n10766), .Y(n11144) );
  INVX1 U2528 ( .A(n11144), .Y(n1390) );
  AND2X1 U2529 ( .A(ram[17]), .B(n10766), .Y(n11131) );
  INVX1 U2530 ( .A(n11131), .Y(n1391) );
  AND2X1 U2531 ( .A(ram[5]), .B(n10766), .Y(n11119) );
  INVX1 U2532 ( .A(n11119), .Y(n1392) );
  AND2X1 U2533 ( .A(n11015), .B(n1836), .Y(n11042) );
  INVX1 U2534 ( .A(n11042), .Y(n1393) );
  BUFX2 U2535 ( .A(n2919), .Y(n1394) );
  BUFX2 U2536 ( .A(n2584), .Y(n1395) );
  AND2X1 U2537 ( .A(n4508), .B(n10956), .Y(n11112) );
  AND2X1 U2538 ( .A(ram[1973]), .B(n10952), .Y(n13204) );
  INVX1 U2539 ( .A(n13204), .Y(n1396) );
  AND2X1 U2540 ( .A(ram[1960]), .B(n10952), .Y(n13178) );
  INVX1 U2541 ( .A(n13178), .Y(n1397) );
  AND2X1 U2542 ( .A(ram[1947]), .B(n10952), .Y(n13152) );
  INVX1 U2543 ( .A(n13152), .Y(n1398) );
  AND2X1 U2544 ( .A(ram[1934]), .B(n10952), .Y(n13126) );
  INVX1 U2545 ( .A(n13126), .Y(n1399) );
  AND2X1 U2546 ( .A(ram[1922]), .B(n10952), .Y(n13102) );
  INVX1 U2547 ( .A(n13102), .Y(n1400) );
  AND2X1 U2548 ( .A(ram[1908]), .B(n10824), .Y(n13083) );
  INVX1 U2549 ( .A(n13083), .Y(n1401) );
  AND2X1 U2550 ( .A(ram[1895]), .B(n10824), .Y(n13070) );
  INVX1 U2551 ( .A(n13070), .Y(n1402) );
  AND2X1 U2552 ( .A(ram[1882]), .B(n10824), .Y(n13057) );
  INVX1 U2553 ( .A(n13057), .Y(n1403) );
  AND2X1 U2554 ( .A(ram[1869]), .B(n10824), .Y(n13044) );
  INVX1 U2555 ( .A(n13044), .Y(n1404) );
  AND2X1 U2556 ( .A(ram[1857]), .B(n10824), .Y(n13032) );
  INVX1 U2557 ( .A(n13032), .Y(n1405) );
  AND2X1 U2558 ( .A(ram[1843]), .B(n10822), .Y(n13016) );
  INVX1 U2559 ( .A(n13016), .Y(n1406) );
  AND2X1 U2560 ( .A(ram[1830]), .B(n10822), .Y(n13003) );
  INVX1 U2561 ( .A(n13003), .Y(n1407) );
  AND2X1 U2562 ( .A(ram[1817]), .B(n10822), .Y(n12990) );
  INVX1 U2563 ( .A(n12990), .Y(n1408) );
  AND2X1 U2564 ( .A(ram[1804]), .B(n10822), .Y(n12977) );
  INVX1 U2565 ( .A(n12977), .Y(n1409) );
  AND2X1 U2566 ( .A(ram[1792]), .B(n10822), .Y(n12965) );
  INVX1 U2567 ( .A(n12965), .Y(n1410) );
  AND2X1 U2568 ( .A(ram[1786]), .B(n10820), .Y(n12957) );
  INVX1 U2569 ( .A(n12957), .Y(n1411) );
  AND2X1 U2570 ( .A(ram[1773]), .B(n10820), .Y(n12944) );
  INVX1 U2571 ( .A(n12944), .Y(n1412) );
  AND2X1 U2572 ( .A(ram[1760]), .B(n10820), .Y(n12931) );
  INVX1 U2573 ( .A(n12931), .Y(n1413) );
  AND2X1 U2574 ( .A(ram[1747]), .B(n10820), .Y(n12918) );
  INVX1 U2575 ( .A(n12918), .Y(n1414) );
  AND2X1 U2576 ( .A(ram[1735]), .B(n10820), .Y(n12906) );
  INVX1 U2577 ( .A(n12906), .Y(n1415) );
  AND2X1 U2578 ( .A(ram[1721]), .B(n10818), .Y(n12890) );
  INVX1 U2579 ( .A(n12890), .Y(n1416) );
  AND2X1 U2580 ( .A(ram[1708]), .B(n10818), .Y(n12877) );
  INVX1 U2581 ( .A(n12877), .Y(n1417) );
  AND2X1 U2582 ( .A(ram[1695]), .B(n10818), .Y(n12864) );
  INVX1 U2583 ( .A(n12864), .Y(n1418) );
  AND2X1 U2584 ( .A(ram[1682]), .B(n10818), .Y(n12851) );
  INVX1 U2585 ( .A(n12851), .Y(n1419) );
  AND2X1 U2586 ( .A(ram[1670]), .B(n10818), .Y(n12839) );
  INVX1 U2587 ( .A(n12839), .Y(n1420) );
  AND2X1 U2588 ( .A(ram[1656]), .B(n10816), .Y(n12823) );
  INVX1 U2589 ( .A(n12823), .Y(n1421) );
  AND2X1 U2590 ( .A(ram[1643]), .B(n10816), .Y(n12810) );
  INVX1 U2591 ( .A(n12810), .Y(n1422) );
  AND2X1 U2592 ( .A(ram[1630]), .B(n10816), .Y(n12797) );
  INVX1 U2593 ( .A(n12797), .Y(n1423) );
  AND2X1 U2594 ( .A(ram[1617]), .B(n10816), .Y(n12784) );
  INVX1 U2595 ( .A(n12784), .Y(n1424) );
  AND2X1 U2596 ( .A(ram[1605]), .B(n10816), .Y(n12772) );
  INVX1 U2597 ( .A(n12772), .Y(n1425) );
  AND2X1 U2598 ( .A(ram[1591]), .B(n10814), .Y(n12756) );
  INVX1 U2599 ( .A(n12756), .Y(n1426) );
  AND2X1 U2600 ( .A(ram[1578]), .B(n10814), .Y(n12743) );
  INVX1 U2601 ( .A(n12743), .Y(n1427) );
  AND2X1 U2602 ( .A(ram[1565]), .B(n10814), .Y(n12730) );
  INVX1 U2603 ( .A(n12730), .Y(n1428) );
  AND2X1 U2604 ( .A(ram[1552]), .B(n10814), .Y(n12717) );
  INVX1 U2605 ( .A(n12717), .Y(n1429) );
  AND2X1 U2606 ( .A(ram[1540]), .B(n10814), .Y(n12705) );
  INVX1 U2607 ( .A(n12705), .Y(n1430) );
  AND2X1 U2608 ( .A(ram[1343]), .B(n10806), .Y(n12499) );
  INVX1 U2609 ( .A(n12499), .Y(n1431) );
  AND2X1 U2610 ( .A(ram[1330]), .B(n10806), .Y(n12486) );
  INVX1 U2611 ( .A(n12486), .Y(n1432) );
  AND2X1 U2612 ( .A(ram[1317]), .B(n10806), .Y(n12473) );
  INVX1 U2613 ( .A(n12473), .Y(n1433) );
  AND2X1 U2614 ( .A(ram[1304]), .B(n10806), .Y(n12460) );
  INVX1 U2615 ( .A(n12460), .Y(n1434) );
  AND2X1 U2616 ( .A(ram[1270]), .B(n10804), .Y(n12424) );
  INVX1 U2617 ( .A(n12424), .Y(n1435) );
  AND2X1 U2618 ( .A(ram[1257]), .B(n10804), .Y(n12411) );
  INVX1 U2619 ( .A(n12411), .Y(n1436) );
  AND2X1 U2620 ( .A(ram[1244]), .B(n10804), .Y(n12398) );
  INVX1 U2621 ( .A(n12398), .Y(n1437) );
  AND2X1 U2622 ( .A(ram[1231]), .B(n10804), .Y(n12385) );
  INVX1 U2623 ( .A(n12385), .Y(n1438) );
  AND2X1 U2624 ( .A(ram[1219]), .B(n10804), .Y(n12373) );
  INVX1 U2625 ( .A(n12373), .Y(n1439) );
  AND2X1 U2626 ( .A(ram[1205]), .B(n10802), .Y(n12357) );
  INVX1 U2627 ( .A(n12357), .Y(n1440) );
  AND2X1 U2628 ( .A(ram[1192]), .B(n10802), .Y(n12344) );
  INVX1 U2629 ( .A(n12344), .Y(n1441) );
  AND2X1 U2630 ( .A(ram[1179]), .B(n10802), .Y(n12331) );
  INVX1 U2631 ( .A(n12331), .Y(n1442) );
  AND2X1 U2632 ( .A(ram[1166]), .B(n10802), .Y(n12318) );
  INVX1 U2633 ( .A(n12318), .Y(n1443) );
  AND2X1 U2634 ( .A(ram[1154]), .B(n10802), .Y(n12306) );
  INVX1 U2635 ( .A(n12306), .Y(n1444) );
  AND2X1 U2636 ( .A(ram[1140]), .B(n10800), .Y(n12290) );
  INVX1 U2637 ( .A(n12290), .Y(n1445) );
  AND2X1 U2638 ( .A(ram[1127]), .B(n10800), .Y(n12277) );
  INVX1 U2639 ( .A(n12277), .Y(n1446) );
  AND2X1 U2640 ( .A(ram[1114]), .B(n10800), .Y(n12264) );
  INVX1 U2641 ( .A(n12264), .Y(n1447) );
  AND2X1 U2642 ( .A(ram[1101]), .B(n10800), .Y(n12251) );
  INVX1 U2643 ( .A(n12251), .Y(n1448) );
  AND2X1 U2644 ( .A(ram[1089]), .B(n10800), .Y(n12239) );
  INVX1 U2645 ( .A(n12239), .Y(n1449) );
  AND2X1 U2646 ( .A(ram[1075]), .B(n10798), .Y(n12223) );
  INVX1 U2647 ( .A(n12223), .Y(n1450) );
  AND2X1 U2648 ( .A(ram[1062]), .B(n10798), .Y(n12210) );
  INVX1 U2649 ( .A(n12210), .Y(n1451) );
  AND2X1 U2650 ( .A(ram[1049]), .B(n10798), .Y(n12197) );
  INVX1 U2651 ( .A(n12197), .Y(n1452) );
  AND2X1 U2652 ( .A(ram[1036]), .B(n10798), .Y(n12184) );
  INVX1 U2653 ( .A(n12184), .Y(n1453) );
  AND2X1 U2654 ( .A(ram[1024]), .B(n10798), .Y(n12172) );
  INVX1 U2655 ( .A(n12172), .Y(n1454) );
  AND2X1 U2656 ( .A(ram[1018]), .B(n10796), .Y(n12164) );
  INVX1 U2657 ( .A(n12164), .Y(n1455) );
  AND2X1 U2658 ( .A(ram[1005]), .B(n10796), .Y(n12151) );
  INVX1 U2659 ( .A(n12151), .Y(n1456) );
  AND2X1 U2660 ( .A(ram[992]), .B(n10796), .Y(n12138) );
  INVX1 U2661 ( .A(n12138), .Y(n1457) );
  AND2X1 U2662 ( .A(ram[979]), .B(n10796), .Y(n12125) );
  INVX1 U2663 ( .A(n12125), .Y(n1458) );
  AND2X1 U2664 ( .A(ram[967]), .B(n10796), .Y(n12113) );
  INVX1 U2665 ( .A(n12113), .Y(n1459) );
  AND2X1 U2666 ( .A(ram[953]), .B(n10794), .Y(n12096) );
  INVX1 U2667 ( .A(n12096), .Y(n1460) );
  AND2X1 U2668 ( .A(ram[940]), .B(n10794), .Y(n12083) );
  INVX1 U2669 ( .A(n12083), .Y(n1461) );
  AND2X1 U2670 ( .A(ram[927]), .B(n10794), .Y(n12070) );
  INVX1 U2671 ( .A(n12070), .Y(n1462) );
  AND2X1 U2672 ( .A(ram[914]), .B(n10794), .Y(n12057) );
  INVX1 U2673 ( .A(n12057), .Y(n1463) );
  AND2X1 U2674 ( .A(ram[902]), .B(n10794), .Y(n12045) );
  INVX1 U2675 ( .A(n12045), .Y(n1464) );
  AND2X1 U2676 ( .A(ram[888]), .B(n10792), .Y(n12029) );
  INVX1 U2677 ( .A(n12029), .Y(n1465) );
  AND2X1 U2678 ( .A(ram[875]), .B(n10792), .Y(n12016) );
  INVX1 U2679 ( .A(n12016), .Y(n1466) );
  AND2X1 U2680 ( .A(ram[862]), .B(n10792), .Y(n12003) );
  INVX1 U2681 ( .A(n12003), .Y(n1467) );
  AND2X1 U2682 ( .A(ram[849]), .B(n10792), .Y(n11990) );
  INVX1 U2683 ( .A(n11990), .Y(n1468) );
  AND2X1 U2684 ( .A(ram[837]), .B(n10792), .Y(n11978) );
  INVX1 U2685 ( .A(n11978), .Y(n1469) );
  AND2X1 U2686 ( .A(ram[823]), .B(n10790), .Y(n11962) );
  INVX1 U2687 ( .A(n11962), .Y(n1470) );
  AND2X1 U2688 ( .A(ram[810]), .B(n10790), .Y(n11949) );
  INVX1 U2689 ( .A(n11949), .Y(n1471) );
  AND2X1 U2690 ( .A(ram[797]), .B(n10790), .Y(n11936) );
  INVX1 U2691 ( .A(n11936), .Y(n1472) );
  AND2X1 U2692 ( .A(ram[784]), .B(n10790), .Y(n11923) );
  INVX1 U2693 ( .A(n11923), .Y(n1473) );
  AND2X1 U2694 ( .A(ram[772]), .B(n10790), .Y(n11911) );
  INVX1 U2695 ( .A(n11911), .Y(n1474) );
  AND2X1 U2696 ( .A(ram[575]), .B(n10782), .Y(n11706) );
  INVX1 U2697 ( .A(n11706), .Y(n1475) );
  AND2X1 U2698 ( .A(ram[562]), .B(n10782), .Y(n11693) );
  INVX1 U2699 ( .A(n11693), .Y(n1476) );
  AND2X1 U2700 ( .A(ram[549]), .B(n10782), .Y(n11680) );
  INVX1 U2701 ( .A(n11680), .Y(n1477) );
  AND2X1 U2702 ( .A(ram[536]), .B(n10782), .Y(n11667) );
  INVX1 U2703 ( .A(n11667), .Y(n1478) );
  AND2X1 U2704 ( .A(ram[502]), .B(n10780), .Y(n11631) );
  INVX1 U2705 ( .A(n11631), .Y(n1479) );
  AND2X1 U2706 ( .A(ram[489]), .B(n10780), .Y(n11618) );
  INVX1 U2707 ( .A(n11618), .Y(n1480) );
  AND2X1 U2708 ( .A(ram[476]), .B(n10780), .Y(n11605) );
  INVX1 U2709 ( .A(n11605), .Y(n1481) );
  AND2X1 U2710 ( .A(ram[463]), .B(n10780), .Y(n11592) );
  INVX1 U2711 ( .A(n11592), .Y(n1482) );
  AND2X1 U2712 ( .A(ram[451]), .B(n10780), .Y(n11580) );
  INVX1 U2713 ( .A(n11580), .Y(n1483) );
  AND2X1 U2714 ( .A(ram[437]), .B(n10778), .Y(n11563) );
  INVX1 U2715 ( .A(n11563), .Y(n1484) );
  AND2X1 U2716 ( .A(ram[424]), .B(n10778), .Y(n11550) );
  INVX1 U2717 ( .A(n11550), .Y(n1485) );
  AND2X1 U2718 ( .A(ram[411]), .B(n10778), .Y(n11537) );
  INVX1 U2719 ( .A(n11537), .Y(n1486) );
  AND2X1 U2720 ( .A(ram[398]), .B(n10778), .Y(n11524) );
  INVX1 U2721 ( .A(n11524), .Y(n1487) );
  AND2X1 U2722 ( .A(ram[386]), .B(n10778), .Y(n11512) );
  INVX1 U2723 ( .A(n11512), .Y(n1488) );
  AND2X1 U2724 ( .A(ram[372]), .B(n10776), .Y(n11496) );
  INVX1 U2725 ( .A(n11496), .Y(n1489) );
  AND2X1 U2726 ( .A(ram[359]), .B(n10776), .Y(n11483) );
  INVX1 U2727 ( .A(n11483), .Y(n1490) );
  AND2X1 U2728 ( .A(ram[346]), .B(n10776), .Y(n11470) );
  INVX1 U2729 ( .A(n11470), .Y(n1491) );
  AND2X1 U2730 ( .A(ram[333]), .B(n10776), .Y(n11457) );
  INVX1 U2731 ( .A(n11457), .Y(n1492) );
  AND2X1 U2732 ( .A(ram[321]), .B(n10776), .Y(n11445) );
  INVX1 U2733 ( .A(n11445), .Y(n1493) );
  AND2X1 U2734 ( .A(ram[307]), .B(n10774), .Y(n11429) );
  INVX1 U2735 ( .A(n11429), .Y(n1494) );
  AND2X1 U2736 ( .A(ram[294]), .B(n10774), .Y(n11416) );
  INVX1 U2737 ( .A(n11416), .Y(n1495) );
  AND2X1 U2738 ( .A(ram[281]), .B(n10774), .Y(n11403) );
  INVX1 U2739 ( .A(n11403), .Y(n1496) );
  AND2X1 U2740 ( .A(ram[268]), .B(n10774), .Y(n11390) );
  INVX1 U2741 ( .A(n11390), .Y(n1497) );
  AND2X1 U2742 ( .A(ram[256]), .B(n10774), .Y(n11378) );
  INVX1 U2743 ( .A(n11378), .Y(n1498) );
  AND2X1 U2744 ( .A(ram[250]), .B(n10772), .Y(n11370) );
  INVX1 U2745 ( .A(n11370), .Y(n1499) );
  AND2X1 U2746 ( .A(ram[237]), .B(n10772), .Y(n11357) );
  INVX1 U2747 ( .A(n11357), .Y(n1500) );
  AND2X1 U2748 ( .A(ram[224]), .B(n10772), .Y(n11344) );
  INVX1 U2749 ( .A(n11344), .Y(n1501) );
  AND2X1 U2750 ( .A(ram[211]), .B(n10772), .Y(n11331) );
  INVX1 U2751 ( .A(n11331), .Y(n1502) );
  AND2X1 U2752 ( .A(ram[199]), .B(n10772), .Y(n11319) );
  INVX1 U2753 ( .A(n11319), .Y(n1503) );
  AND2X1 U2754 ( .A(ram[185]), .B(n10770), .Y(n11303) );
  INVX1 U2755 ( .A(n11303), .Y(n1504) );
  AND2X1 U2756 ( .A(ram[172]), .B(n10770), .Y(n11290) );
  INVX1 U2757 ( .A(n11290), .Y(n1505) );
  AND2X1 U2758 ( .A(ram[159]), .B(n10770), .Y(n11277) );
  INVX1 U2759 ( .A(n11277), .Y(n1506) );
  AND2X1 U2760 ( .A(ram[146]), .B(n10770), .Y(n11264) );
  INVX1 U2761 ( .A(n11264), .Y(n1507) );
  AND2X1 U2762 ( .A(ram[134]), .B(n10770), .Y(n11252) );
  INVX1 U2763 ( .A(n11252), .Y(n1508) );
  AND2X1 U2764 ( .A(ram[120]), .B(n10768), .Y(n11236) );
  INVX1 U2765 ( .A(n11236), .Y(n1509) );
  AND2X1 U2766 ( .A(ram[107]), .B(n10768), .Y(n11223) );
  INVX1 U2767 ( .A(n11223), .Y(n1510) );
  AND2X1 U2768 ( .A(ram[94]), .B(n10768), .Y(n11210) );
  INVX1 U2769 ( .A(n11210), .Y(n1511) );
  AND2X1 U2770 ( .A(ram[81]), .B(n10768), .Y(n11197) );
  INVX1 U2771 ( .A(n11197), .Y(n1512) );
  AND2X1 U2772 ( .A(ram[69]), .B(n10768), .Y(n11185) );
  INVX1 U2773 ( .A(n11185), .Y(n1513) );
  AND2X1 U2774 ( .A(ram[55]), .B(n10766), .Y(n11169) );
  INVX1 U2775 ( .A(n11169), .Y(n1514) );
  AND2X1 U2776 ( .A(ram[42]), .B(n10766), .Y(n11156) );
  INVX1 U2777 ( .A(n11156), .Y(n1515) );
  AND2X1 U2778 ( .A(ram[29]), .B(n10766), .Y(n11143) );
  INVX1 U2779 ( .A(n11143), .Y(n1516) );
  AND2X1 U2780 ( .A(ram[16]), .B(n10766), .Y(n11130) );
  INVX1 U2781 ( .A(n11130), .Y(n1517) );
  AND2X1 U2782 ( .A(ram[4]), .B(n10766), .Y(n11118) );
  INVX1 U2783 ( .A(n11118), .Y(n1518) );
  AND2X1 U2784 ( .A(n11015), .B(n2152), .Y(n11003) );
  INVX1 U2785 ( .A(n11003), .Y(n1519) );
  BUFX2 U2786 ( .A(n2517), .Y(n1520) );
  AND2X1 U2787 ( .A(ram[1976]), .B(n10952), .Y(n13210) );
  INVX1 U2788 ( .A(n13210), .Y(n1521) );
  AND2X1 U2789 ( .A(ram[1963]), .B(n10952), .Y(n13184) );
  INVX1 U2790 ( .A(n13184), .Y(n1522) );
  AND2X1 U2791 ( .A(ram[1950]), .B(n10952), .Y(n13158) );
  INVX1 U2792 ( .A(n13158), .Y(n1523) );
  AND2X1 U2793 ( .A(ram[1937]), .B(n10952), .Y(n13132) );
  INVX1 U2794 ( .A(n13132), .Y(n1524) );
  AND2X1 U2795 ( .A(ram[1925]), .B(n10952), .Y(n13108) );
  INVX1 U2796 ( .A(n13108), .Y(n1525) );
  AND2X1 U2797 ( .A(ram[1913]), .B(n10824), .Y(n13088) );
  INVX1 U2798 ( .A(n13088), .Y(n1526) );
  AND2X1 U2799 ( .A(ram[1900]), .B(n10824), .Y(n13075) );
  INVX1 U2800 ( .A(n13075), .Y(n1527) );
  AND2X1 U2801 ( .A(ram[1887]), .B(n10824), .Y(n13062) );
  INVX1 U2802 ( .A(n13062), .Y(n1528) );
  AND2X1 U2803 ( .A(ram[1874]), .B(n10824), .Y(n13049) );
  INVX1 U2804 ( .A(n13049), .Y(n1529) );
  AND2X1 U2805 ( .A(ram[1862]), .B(n10824), .Y(n13037) );
  INVX1 U2806 ( .A(n13037), .Y(n1530) );
  AND2X1 U2807 ( .A(ram[1850]), .B(n10822), .Y(n13023) );
  INVX1 U2808 ( .A(n13023), .Y(n1531) );
  AND2X1 U2809 ( .A(ram[1837]), .B(n10822), .Y(n13010) );
  INVX1 U2810 ( .A(n13010), .Y(n1532) );
  AND2X1 U2811 ( .A(ram[1824]), .B(n10822), .Y(n12997) );
  INVX1 U2812 ( .A(n12997), .Y(n1533) );
  AND2X1 U2813 ( .A(ram[1811]), .B(n10822), .Y(n12984) );
  INVX1 U2814 ( .A(n12984), .Y(n1534) );
  AND2X1 U2815 ( .A(ram[1799]), .B(n10822), .Y(n12972) );
  INVX1 U2816 ( .A(n12972), .Y(n1535) );
  AND2X1 U2817 ( .A(ram[1779]), .B(n10820), .Y(n12950) );
  INVX1 U2818 ( .A(n12950), .Y(n1536) );
  AND2X1 U2819 ( .A(ram[1766]), .B(n10820), .Y(n12937) );
  INVX1 U2820 ( .A(n12937), .Y(n1537) );
  AND2X1 U2821 ( .A(ram[1753]), .B(n10820), .Y(n12924) );
  INVX1 U2822 ( .A(n12924), .Y(n1538) );
  AND2X1 U2823 ( .A(ram[1740]), .B(n10820), .Y(n12911) );
  INVX1 U2824 ( .A(n12911), .Y(n1539) );
  AND2X1 U2825 ( .A(ram[1728]), .B(n10820), .Y(n12899) );
  INVX1 U2826 ( .A(n12899), .Y(n1540) );
  AND2X1 U2827 ( .A(ram[1716]), .B(n10818), .Y(n12885) );
  INVX1 U2828 ( .A(n12885), .Y(n1541) );
  AND2X1 U2829 ( .A(ram[1703]), .B(n10818), .Y(n12872) );
  INVX1 U2830 ( .A(n12872), .Y(n1542) );
  AND2X1 U2831 ( .A(ram[1690]), .B(n10818), .Y(n12859) );
  INVX1 U2832 ( .A(n12859), .Y(n1543) );
  AND2X1 U2833 ( .A(ram[1677]), .B(n10818), .Y(n12846) );
  INVX1 U2834 ( .A(n12846), .Y(n1544) );
  AND2X1 U2835 ( .A(ram[1665]), .B(n10818), .Y(n12834) );
  INVX1 U2836 ( .A(n12834), .Y(n1545) );
  AND2X1 U2837 ( .A(ram[1653]), .B(n10816), .Y(n12820) );
  INVX1 U2838 ( .A(n12820), .Y(n1546) );
  AND2X1 U2839 ( .A(ram[1640]), .B(n10816), .Y(n12807) );
  INVX1 U2840 ( .A(n12807), .Y(n1547) );
  AND2X1 U2841 ( .A(ram[1627]), .B(n10816), .Y(n12794) );
  INVX1 U2842 ( .A(n12794), .Y(n1548) );
  AND2X1 U2843 ( .A(ram[1614]), .B(n10816), .Y(n12781) );
  INVX1 U2844 ( .A(n12781), .Y(n1549) );
  AND2X1 U2845 ( .A(ram[1602]), .B(n10816), .Y(n12769) );
  INVX1 U2846 ( .A(n12769), .Y(n1550) );
  AND2X1 U2847 ( .A(ram[1590]), .B(n10814), .Y(n12755) );
  INVX1 U2848 ( .A(n12755), .Y(n1551) );
  AND2X1 U2849 ( .A(ram[1577]), .B(n10814), .Y(n12742) );
  INVX1 U2850 ( .A(n12742), .Y(n1552) );
  AND2X1 U2851 ( .A(ram[1564]), .B(n10814), .Y(n12729) );
  INVX1 U2852 ( .A(n12729), .Y(n1553) );
  AND2X1 U2853 ( .A(ram[1551]), .B(n10814), .Y(n12716) );
  INVX1 U2854 ( .A(n12716), .Y(n1554) );
  AND2X1 U2855 ( .A(ram[1539]), .B(n10814), .Y(n12704) );
  INVX1 U2856 ( .A(n12704), .Y(n1555) );
  AND2X1 U2857 ( .A(ram[1531]), .B(n10812), .Y(n12694) );
  INVX1 U2858 ( .A(n12694), .Y(n1556) );
  AND2X1 U2859 ( .A(ram[1518]), .B(n10812), .Y(n12681) );
  INVX1 U2860 ( .A(n12681), .Y(n1557) );
  AND2X1 U2861 ( .A(ram[1505]), .B(n10812), .Y(n12668) );
  INVX1 U2862 ( .A(n12668), .Y(n1558) );
  AND2X1 U2863 ( .A(ram[1492]), .B(n10812), .Y(n12655) );
  INVX1 U2864 ( .A(n12655), .Y(n1559) );
  AND2X1 U2865 ( .A(ram[1480]), .B(n10812), .Y(n12643) );
  INVX1 U2866 ( .A(n12643), .Y(n1560) );
  AND2X1 U2867 ( .A(ram[1468]), .B(n10810), .Y(n12628) );
  INVX1 U2868 ( .A(n12628), .Y(n1561) );
  AND2X1 U2869 ( .A(ram[1455]), .B(n10810), .Y(n12615) );
  INVX1 U2870 ( .A(n12615), .Y(n1562) );
  AND2X1 U2871 ( .A(ram[1442]), .B(n10810), .Y(n12602) );
  INVX1 U2872 ( .A(n12602), .Y(n1563) );
  AND2X1 U2873 ( .A(ram[1429]), .B(n10810), .Y(n12589) );
  INVX1 U2874 ( .A(n12589), .Y(n1564) );
  AND2X1 U2875 ( .A(ram[1417]), .B(n10810), .Y(n12577) );
  INVX1 U2876 ( .A(n12577), .Y(n1565) );
  AND2X1 U2877 ( .A(ram[1405]), .B(n10808), .Y(n12563) );
  INVX1 U2878 ( .A(n12563), .Y(n1566) );
  AND2X1 U2879 ( .A(ram[1392]), .B(n10808), .Y(n12550) );
  INVX1 U2880 ( .A(n12550), .Y(n1567) );
  AND2X1 U2881 ( .A(ram[1379]), .B(n10808), .Y(n12537) );
  INVX1 U2882 ( .A(n12537), .Y(n1568) );
  AND2X1 U2883 ( .A(ram[1366]), .B(n10808), .Y(n12524) );
  INVX1 U2884 ( .A(n12524), .Y(n1569) );
  AND2X1 U2885 ( .A(ram[1354]), .B(n10808), .Y(n12512) );
  INVX1 U2886 ( .A(n12512), .Y(n1570) );
  AND2X1 U2887 ( .A(ram[1342]), .B(n10806), .Y(n12498) );
  INVX1 U2888 ( .A(n12498), .Y(n1571) );
  AND2X1 U2889 ( .A(ram[1329]), .B(n10806), .Y(n12485) );
  INVX1 U2890 ( .A(n12485), .Y(n1572) );
  AND2X1 U2891 ( .A(ram[1316]), .B(n10806), .Y(n12472) );
  INVX1 U2892 ( .A(n12472), .Y(n1573) );
  AND2X1 U2893 ( .A(ram[1303]), .B(n10806), .Y(n12459) );
  INVX1 U2894 ( .A(n12459), .Y(n1574) );
  AND2X1 U2895 ( .A(ram[1291]), .B(n10806), .Y(n12447) );
  INVX1 U2896 ( .A(n12447), .Y(n1575) );
  AND2X1 U2897 ( .A(ram[1271]), .B(n10804), .Y(n12425) );
  INVX1 U2898 ( .A(n12425), .Y(n1576) );
  AND2X1 U2899 ( .A(ram[1258]), .B(n10804), .Y(n12412) );
  INVX1 U2900 ( .A(n12412), .Y(n1577) );
  AND2X1 U2901 ( .A(ram[1245]), .B(n10804), .Y(n12399) );
  INVX1 U2902 ( .A(n12399), .Y(n1578) );
  AND2X1 U2903 ( .A(ram[1232]), .B(n10804), .Y(n12386) );
  INVX1 U2904 ( .A(n12386), .Y(n1579) );
  AND2X1 U2905 ( .A(ram[1220]), .B(n10804), .Y(n12374) );
  INVX1 U2906 ( .A(n12374), .Y(n1580) );
  AND2X1 U2907 ( .A(ram[1208]), .B(n10802), .Y(n12360) );
  INVX1 U2908 ( .A(n12360), .Y(n1581) );
  AND2X1 U2909 ( .A(ram[1195]), .B(n10802), .Y(n12347) );
  INVX1 U2910 ( .A(n12347), .Y(n1582) );
  AND2X1 U2911 ( .A(ram[1182]), .B(n10802), .Y(n12334) );
  INVX1 U2912 ( .A(n12334), .Y(n1583) );
  AND2X1 U2913 ( .A(ram[1169]), .B(n10802), .Y(n12321) );
  INVX1 U2914 ( .A(n12321), .Y(n1584) );
  AND2X1 U2915 ( .A(ram[1157]), .B(n10802), .Y(n12309) );
  INVX1 U2916 ( .A(n12309), .Y(n1585) );
  AND2X1 U2917 ( .A(ram[1145]), .B(n10800), .Y(n12295) );
  INVX1 U2918 ( .A(n12295), .Y(n1586) );
  AND2X1 U2919 ( .A(ram[1132]), .B(n10800), .Y(n12282) );
  INVX1 U2920 ( .A(n12282), .Y(n1587) );
  AND2X1 U2921 ( .A(ram[1119]), .B(n10800), .Y(n12269) );
  INVX1 U2922 ( .A(n12269), .Y(n1588) );
  AND2X1 U2923 ( .A(ram[1106]), .B(n10800), .Y(n12256) );
  INVX1 U2924 ( .A(n12256), .Y(n1589) );
  AND2X1 U2925 ( .A(ram[1094]), .B(n10800), .Y(n12244) );
  INVX1 U2926 ( .A(n12244), .Y(n1590) );
  AND2X1 U2927 ( .A(ram[1082]), .B(n10798), .Y(n12230) );
  INVX1 U2928 ( .A(n12230), .Y(n1591) );
  AND2X1 U2929 ( .A(ram[1069]), .B(n10798), .Y(n12217) );
  INVX1 U2930 ( .A(n12217), .Y(n1592) );
  AND2X1 U2931 ( .A(ram[1056]), .B(n10798), .Y(n12204) );
  INVX1 U2932 ( .A(n12204), .Y(n1593) );
  AND2X1 U2933 ( .A(ram[1043]), .B(n10798), .Y(n12191) );
  INVX1 U2934 ( .A(n12191), .Y(n1594) );
  AND2X1 U2935 ( .A(ram[1031]), .B(n10798), .Y(n12179) );
  INVX1 U2936 ( .A(n12179), .Y(n1595) );
  AND2X1 U2937 ( .A(ram[1011]), .B(n10796), .Y(n12157) );
  INVX1 U2938 ( .A(n12157), .Y(n1596) );
  AND2X1 U2939 ( .A(ram[998]), .B(n10796), .Y(n12144) );
  INVX1 U2940 ( .A(n12144), .Y(n1597) );
  AND2X1 U2941 ( .A(ram[985]), .B(n10796), .Y(n12131) );
  INVX1 U2942 ( .A(n12131), .Y(n1598) );
  AND2X1 U2943 ( .A(ram[972]), .B(n10796), .Y(n12118) );
  INVX1 U2944 ( .A(n12118), .Y(n1599) );
  AND2X1 U2945 ( .A(ram[960]), .B(n10796), .Y(n12106) );
  INVX1 U2946 ( .A(n12106), .Y(n1600) );
  AND2X1 U2947 ( .A(ram[948]), .B(n10794), .Y(n12091) );
  INVX1 U2948 ( .A(n12091), .Y(n1601) );
  AND2X1 U2949 ( .A(ram[935]), .B(n10794), .Y(n12078) );
  INVX1 U2950 ( .A(n12078), .Y(n1602) );
  AND2X1 U2951 ( .A(ram[922]), .B(n10794), .Y(n12065) );
  INVX1 U2952 ( .A(n12065), .Y(n1603) );
  AND2X1 U2953 ( .A(ram[909]), .B(n10794), .Y(n12052) );
  INVX1 U2954 ( .A(n12052), .Y(n1604) );
  AND2X1 U2955 ( .A(ram[897]), .B(n10794), .Y(n12040) );
  INVX1 U2956 ( .A(n12040), .Y(n1605) );
  AND2X1 U2957 ( .A(ram[885]), .B(n10792), .Y(n12026) );
  INVX1 U2958 ( .A(n12026), .Y(n1606) );
  AND2X1 U2959 ( .A(ram[872]), .B(n10792), .Y(n12013) );
  INVX1 U2960 ( .A(n12013), .Y(n1607) );
  AND2X1 U2961 ( .A(ram[859]), .B(n10792), .Y(n12000) );
  INVX1 U2962 ( .A(n12000), .Y(n1608) );
  AND2X1 U2963 ( .A(ram[846]), .B(n10792), .Y(n11987) );
  INVX1 U2964 ( .A(n11987), .Y(n1609) );
  AND2X1 U2965 ( .A(ram[834]), .B(n10792), .Y(n11975) );
  INVX1 U2966 ( .A(n11975), .Y(n1610) );
  AND2X1 U2967 ( .A(ram[822]), .B(n10790), .Y(n11961) );
  INVX1 U2968 ( .A(n11961), .Y(n1611) );
  AND2X1 U2969 ( .A(ram[809]), .B(n10790), .Y(n11948) );
  INVX1 U2970 ( .A(n11948), .Y(n1612) );
  AND2X1 U2971 ( .A(ram[796]), .B(n10790), .Y(n11935) );
  INVX1 U2972 ( .A(n11935), .Y(n1613) );
  AND2X1 U2973 ( .A(ram[783]), .B(n10790), .Y(n11922) );
  INVX1 U2974 ( .A(n11922), .Y(n1614) );
  AND2X1 U2975 ( .A(ram[771]), .B(n10790), .Y(n11910) );
  INVX1 U2976 ( .A(n11910), .Y(n1615) );
  AND2X1 U2977 ( .A(ram[763]), .B(n10788), .Y(n11900) );
  INVX1 U2978 ( .A(n11900), .Y(n1616) );
  AND2X1 U2979 ( .A(ram[750]), .B(n10788), .Y(n11887) );
  INVX1 U2980 ( .A(n11887), .Y(n1617) );
  AND2X1 U2981 ( .A(ram[737]), .B(n10788), .Y(n11874) );
  INVX1 U2982 ( .A(n11874), .Y(n1618) );
  AND2X1 U2983 ( .A(ram[724]), .B(n10788), .Y(n11861) );
  INVX1 U2984 ( .A(n11861), .Y(n1619) );
  AND2X1 U2985 ( .A(ram[712]), .B(n10788), .Y(n11849) );
  INVX1 U2986 ( .A(n11849), .Y(n1620) );
  AND2X1 U2987 ( .A(ram[700]), .B(n10786), .Y(n11835) );
  INVX1 U2988 ( .A(n11835), .Y(n1621) );
  AND2X1 U2989 ( .A(ram[687]), .B(n10786), .Y(n11822) );
  INVX1 U2990 ( .A(n11822), .Y(n1622) );
  AND2X1 U2991 ( .A(ram[674]), .B(n10786), .Y(n11809) );
  INVX1 U2992 ( .A(n11809), .Y(n1623) );
  AND2X1 U2993 ( .A(ram[661]), .B(n10786), .Y(n11796) );
  INVX1 U2994 ( .A(n11796), .Y(n1624) );
  AND2X1 U2995 ( .A(ram[649]), .B(n10786), .Y(n11784) );
  INVX1 U2996 ( .A(n11784), .Y(n1625) );
  AND2X1 U2997 ( .A(ram[637]), .B(n10784), .Y(n11770) );
  INVX1 U2998 ( .A(n11770), .Y(n1626) );
  AND2X1 U2999 ( .A(ram[624]), .B(n10784), .Y(n11757) );
  INVX1 U3000 ( .A(n11757), .Y(n1627) );
  AND2X1 U3001 ( .A(ram[611]), .B(n10784), .Y(n11744) );
  INVX1 U3002 ( .A(n11744), .Y(n1628) );
  AND2X1 U3003 ( .A(ram[598]), .B(n10784), .Y(n11731) );
  INVX1 U3004 ( .A(n11731), .Y(n1629) );
  AND2X1 U3005 ( .A(ram[586]), .B(n10784), .Y(n11719) );
  INVX1 U3006 ( .A(n11719), .Y(n1630) );
  AND2X1 U3007 ( .A(ram[574]), .B(n10782), .Y(n11705) );
  INVX1 U3008 ( .A(n11705), .Y(n1631) );
  AND2X1 U3009 ( .A(ram[561]), .B(n10782), .Y(n11692) );
  INVX1 U3010 ( .A(n11692), .Y(n1632) );
  AND2X1 U3011 ( .A(ram[548]), .B(n10782), .Y(n11679) );
  INVX1 U3012 ( .A(n11679), .Y(n1633) );
  AND2X1 U3013 ( .A(ram[535]), .B(n10782), .Y(n11666) );
  INVX1 U3014 ( .A(n11666), .Y(n1634) );
  AND2X1 U3015 ( .A(ram[523]), .B(n10782), .Y(n11654) );
  INVX1 U3016 ( .A(n11654), .Y(n1635) );
  AND2X1 U3017 ( .A(ram[503]), .B(n10780), .Y(n11632) );
  INVX1 U3018 ( .A(n11632), .Y(n1636) );
  AND2X1 U3019 ( .A(ram[490]), .B(n10780), .Y(n11619) );
  INVX1 U3020 ( .A(n11619), .Y(n1637) );
  AND2X1 U3021 ( .A(ram[477]), .B(n10780), .Y(n11606) );
  INVX1 U3022 ( .A(n11606), .Y(n1638) );
  AND2X1 U3023 ( .A(ram[464]), .B(n10780), .Y(n11593) );
  INVX1 U3024 ( .A(n11593), .Y(n1639) );
  AND2X1 U3025 ( .A(ram[452]), .B(n10780), .Y(n11581) );
  INVX1 U3026 ( .A(n11581), .Y(n1640) );
  AND2X1 U3027 ( .A(ram[440]), .B(n10778), .Y(n11566) );
  INVX1 U3028 ( .A(n11566), .Y(n1641) );
  AND2X1 U3029 ( .A(ram[427]), .B(n10778), .Y(n11553) );
  INVX1 U3030 ( .A(n11553), .Y(n1642) );
  AND2X1 U3031 ( .A(ram[414]), .B(n10778), .Y(n11540) );
  INVX1 U3032 ( .A(n11540), .Y(n1643) );
  AND2X1 U3033 ( .A(ram[401]), .B(n10778), .Y(n11527) );
  INVX1 U3034 ( .A(n11527), .Y(n1644) );
  AND2X1 U3035 ( .A(ram[389]), .B(n10778), .Y(n11515) );
  INVX1 U3036 ( .A(n11515), .Y(n1645) );
  AND2X1 U3037 ( .A(ram[377]), .B(n10776), .Y(n11501) );
  INVX1 U3038 ( .A(n11501), .Y(n1646) );
  AND2X1 U3039 ( .A(ram[364]), .B(n10776), .Y(n11488) );
  INVX1 U3040 ( .A(n11488), .Y(n1647) );
  AND2X1 U3041 ( .A(ram[351]), .B(n10776), .Y(n11475) );
  INVX1 U3042 ( .A(n11475), .Y(n1648) );
  AND2X1 U3043 ( .A(ram[338]), .B(n10776), .Y(n11462) );
  INVX1 U3044 ( .A(n11462), .Y(n1649) );
  AND2X1 U3045 ( .A(ram[326]), .B(n10776), .Y(n11450) );
  INVX1 U3046 ( .A(n11450), .Y(n1650) );
  AND2X1 U3047 ( .A(ram[314]), .B(n10774), .Y(n11436) );
  INVX1 U3048 ( .A(n11436), .Y(n1651) );
  AND2X1 U3049 ( .A(ram[301]), .B(n10774), .Y(n11423) );
  INVX1 U3050 ( .A(n11423), .Y(n1652) );
  AND2X1 U3051 ( .A(ram[288]), .B(n10774), .Y(n11410) );
  INVX1 U3052 ( .A(n11410), .Y(n1653) );
  AND2X1 U3053 ( .A(ram[275]), .B(n10774), .Y(n11397) );
  INVX1 U3054 ( .A(n11397), .Y(n1654) );
  AND2X1 U3055 ( .A(ram[263]), .B(n10774), .Y(n11385) );
  INVX1 U3056 ( .A(n11385), .Y(n1655) );
  AND2X1 U3057 ( .A(ram[243]), .B(n10772), .Y(n11363) );
  INVX1 U3058 ( .A(n11363), .Y(n1656) );
  AND2X1 U3059 ( .A(ram[230]), .B(n10772), .Y(n11350) );
  INVX1 U3060 ( .A(n11350), .Y(n1657) );
  AND2X1 U3061 ( .A(ram[217]), .B(n10772), .Y(n11337) );
  INVX1 U3062 ( .A(n11337), .Y(n1658) );
  AND2X1 U3063 ( .A(ram[204]), .B(n10772), .Y(n11324) );
  INVX1 U3064 ( .A(n11324), .Y(n1659) );
  AND2X1 U3065 ( .A(ram[192]), .B(n10772), .Y(n11312) );
  INVX1 U3066 ( .A(n11312), .Y(n1660) );
  AND2X1 U3067 ( .A(ram[180]), .B(n10770), .Y(n11298) );
  INVX1 U3068 ( .A(n11298), .Y(n1661) );
  AND2X1 U3069 ( .A(ram[167]), .B(n10770), .Y(n11285) );
  INVX1 U3070 ( .A(n11285), .Y(n1662) );
  AND2X1 U3071 ( .A(ram[154]), .B(n10770), .Y(n11272) );
  INVX1 U3072 ( .A(n11272), .Y(n1663) );
  AND2X1 U3073 ( .A(ram[141]), .B(n10770), .Y(n11259) );
  INVX1 U3074 ( .A(n11259), .Y(n1664) );
  AND2X1 U3075 ( .A(ram[129]), .B(n10770), .Y(n11247) );
  INVX1 U3076 ( .A(n11247), .Y(n1665) );
  AND2X1 U3077 ( .A(ram[117]), .B(n10768), .Y(n11233) );
  INVX1 U3078 ( .A(n11233), .Y(n1666) );
  AND2X1 U3079 ( .A(ram[104]), .B(n10768), .Y(n11220) );
  INVX1 U3080 ( .A(n11220), .Y(n1667) );
  AND2X1 U3081 ( .A(ram[91]), .B(n10768), .Y(n11207) );
  INVX1 U3082 ( .A(n11207), .Y(n1668) );
  AND2X1 U3083 ( .A(ram[78]), .B(n10768), .Y(n11194) );
  INVX1 U3084 ( .A(n11194), .Y(n1669) );
  AND2X1 U3085 ( .A(ram[66]), .B(n10768), .Y(n11182) );
  INVX1 U3086 ( .A(n11182), .Y(n1670) );
  AND2X1 U3087 ( .A(ram[54]), .B(n10766), .Y(n11168) );
  INVX1 U3088 ( .A(n11168), .Y(n1671) );
  AND2X1 U3089 ( .A(ram[41]), .B(n10766), .Y(n11155) );
  INVX1 U3090 ( .A(n11155), .Y(n1672) );
  AND2X1 U3091 ( .A(ram[28]), .B(n10766), .Y(n11142) );
  INVX1 U3092 ( .A(n11142), .Y(n1673) );
  AND2X1 U3093 ( .A(ram[15]), .B(n10766), .Y(n11129) );
  INVX1 U3094 ( .A(n11129), .Y(n1674) );
  AND2X1 U3095 ( .A(ram[3]), .B(n10766), .Y(n11117) );
  INVX1 U3096 ( .A(n11117), .Y(n1675) );
  AND2X1 U3097 ( .A(n1993), .B(n1836), .Y(n11033) );
  INVX1 U3098 ( .A(n11033), .Y(n1676) );
  BUFX2 U3099 ( .A(n10977), .Y(n1677) );
  BUFX2 U3100 ( .A(n2986), .Y(n1678) );
  BUFX2 U3101 ( .A(n13096), .Y(n1679) );
  AND2X1 U3102 ( .A(ram[1975]), .B(n10952), .Y(n13208) );
  INVX1 U3103 ( .A(n13208), .Y(n1680) );
  AND2X1 U3104 ( .A(ram[1962]), .B(n10952), .Y(n13182) );
  INVX1 U3105 ( .A(n13182), .Y(n1681) );
  AND2X1 U3106 ( .A(ram[1949]), .B(n10952), .Y(n13156) );
  INVX1 U3107 ( .A(n13156), .Y(n1682) );
  AND2X1 U3108 ( .A(ram[1936]), .B(n10952), .Y(n13130) );
  INVX1 U3109 ( .A(n13130), .Y(n1683) );
  AND2X1 U3110 ( .A(ram[1924]), .B(n10952), .Y(n13106) );
  INVX1 U3111 ( .A(n13106), .Y(n1684) );
  AND2X1 U3112 ( .A(ram[1914]), .B(n10824), .Y(n13089) );
  INVX1 U3113 ( .A(n13089), .Y(n1685) );
  AND2X1 U3114 ( .A(ram[1901]), .B(n10824), .Y(n13076) );
  INVX1 U3115 ( .A(n13076), .Y(n1686) );
  AND2X1 U3116 ( .A(ram[1888]), .B(n10824), .Y(n13063) );
  INVX1 U3117 ( .A(n13063), .Y(n1687) );
  AND2X1 U3118 ( .A(ram[1875]), .B(n10824), .Y(n13050) );
  INVX1 U3119 ( .A(n13050), .Y(n1688) );
  AND2X1 U3120 ( .A(ram[1863]), .B(n10824), .Y(n13038) );
  INVX1 U3121 ( .A(n13038), .Y(n1689) );
  AND2X1 U3122 ( .A(ram[1849]), .B(n10822), .Y(n13022) );
  INVX1 U3123 ( .A(n13022), .Y(n1690) );
  AND2X1 U3124 ( .A(ram[1836]), .B(n10822), .Y(n13009) );
  INVX1 U3125 ( .A(n13009), .Y(n1691) );
  AND2X1 U3126 ( .A(ram[1823]), .B(n10822), .Y(n12996) );
  INVX1 U3127 ( .A(n12996), .Y(n1692) );
  AND2X1 U3128 ( .A(ram[1810]), .B(n10822), .Y(n12983) );
  INVX1 U3129 ( .A(n12983), .Y(n1693) );
  AND2X1 U3130 ( .A(ram[1798]), .B(n10822), .Y(n12971) );
  INVX1 U3131 ( .A(n12971), .Y(n1694) );
  AND2X1 U3132 ( .A(ram[1780]), .B(n10820), .Y(n12951) );
  INVX1 U3133 ( .A(n12951), .Y(n1695) );
  AND2X1 U3134 ( .A(ram[1767]), .B(n10820), .Y(n12938) );
  INVX1 U3135 ( .A(n12938), .Y(n1696) );
  AND2X1 U3136 ( .A(ram[1754]), .B(n10820), .Y(n12925) );
  INVX1 U3137 ( .A(n12925), .Y(n1697) );
  AND2X1 U3138 ( .A(ram[1741]), .B(n10820), .Y(n12912) );
  INVX1 U3139 ( .A(n12912), .Y(n1698) );
  AND2X1 U3140 ( .A(ram[1729]), .B(n10820), .Y(n12900) );
  INVX1 U3141 ( .A(n12900), .Y(n1699) );
  AND2X1 U3142 ( .A(ram[1715]), .B(n10818), .Y(n12884) );
  INVX1 U3143 ( .A(n12884), .Y(n1700) );
  AND2X1 U3144 ( .A(ram[1702]), .B(n10818), .Y(n12871) );
  INVX1 U3145 ( .A(n12871), .Y(n1701) );
  AND2X1 U3146 ( .A(ram[1689]), .B(n10818), .Y(n12858) );
  INVX1 U3147 ( .A(n12858), .Y(n1702) );
  AND2X1 U3148 ( .A(ram[1676]), .B(n10818), .Y(n12845) );
  INVX1 U3149 ( .A(n12845), .Y(n1703) );
  AND2X1 U3150 ( .A(ram[1664]), .B(n10818), .Y(n12833) );
  INVX1 U3151 ( .A(n12833), .Y(n1704) );
  AND2X1 U3152 ( .A(ram[1654]), .B(n10816), .Y(n12821) );
  INVX1 U3153 ( .A(n12821), .Y(n1705) );
  AND2X1 U3154 ( .A(ram[1641]), .B(n10816), .Y(n12808) );
  INVX1 U3155 ( .A(n12808), .Y(n1706) );
  AND2X1 U3156 ( .A(ram[1628]), .B(n10816), .Y(n12795) );
  INVX1 U3157 ( .A(n12795), .Y(n1707) );
  AND2X1 U3158 ( .A(ram[1615]), .B(n10816), .Y(n12782) );
  INVX1 U3159 ( .A(n12782), .Y(n1708) );
  AND2X1 U3160 ( .A(ram[1603]), .B(n10816), .Y(n12770) );
  INVX1 U3161 ( .A(n12770), .Y(n1709) );
  AND2X1 U3162 ( .A(ram[1589]), .B(n10814), .Y(n12754) );
  INVX1 U3163 ( .A(n12754), .Y(n1710) );
  AND2X1 U3164 ( .A(ram[1576]), .B(n10814), .Y(n12741) );
  INVX1 U3165 ( .A(n12741), .Y(n1711) );
  AND2X1 U3166 ( .A(ram[1563]), .B(n10814), .Y(n12728) );
  INVX1 U3167 ( .A(n12728), .Y(n1712) );
  AND2X1 U3168 ( .A(ram[1550]), .B(n10814), .Y(n12715) );
  INVX1 U3169 ( .A(n12715), .Y(n1713) );
  AND2X1 U3170 ( .A(ram[1538]), .B(n10814), .Y(n12703) );
  INVX1 U3171 ( .A(n12703), .Y(n1714) );
  AND2X1 U3172 ( .A(ram[1532]), .B(n10812), .Y(n12695) );
  INVX1 U3173 ( .A(n12695), .Y(n1715) );
  AND2X1 U3174 ( .A(ram[1519]), .B(n10812), .Y(n12682) );
  INVX1 U3175 ( .A(n12682), .Y(n1716) );
  AND2X1 U3176 ( .A(ram[1506]), .B(n10812), .Y(n12669) );
  INVX1 U3177 ( .A(n12669), .Y(n1717) );
  AND2X1 U3178 ( .A(ram[1493]), .B(n10812), .Y(n12656) );
  INVX1 U3179 ( .A(n12656), .Y(n1718) );
  AND2X1 U3180 ( .A(ram[1481]), .B(n10812), .Y(n12644) );
  INVX1 U3181 ( .A(n12644), .Y(n1719) );
  AND2X1 U3182 ( .A(ram[1467]), .B(n10810), .Y(n12627) );
  INVX1 U3183 ( .A(n12627), .Y(n1720) );
  AND2X1 U3184 ( .A(ram[1454]), .B(n10810), .Y(n12614) );
  INVX1 U3185 ( .A(n12614), .Y(n1721) );
  AND2X1 U3186 ( .A(ram[1441]), .B(n10810), .Y(n12601) );
  INVX1 U3187 ( .A(n12601), .Y(n1722) );
  AND2X1 U3188 ( .A(ram[1428]), .B(n10810), .Y(n12588) );
  INVX1 U3189 ( .A(n12588), .Y(n1723) );
  AND2X1 U3190 ( .A(ram[1416]), .B(n10810), .Y(n12576) );
  INVX1 U3191 ( .A(n12576), .Y(n1724) );
  AND2X1 U3192 ( .A(ram[1406]), .B(n10808), .Y(n12564) );
  INVX1 U3193 ( .A(n12564), .Y(n1725) );
  AND2X1 U3194 ( .A(ram[1393]), .B(n10808), .Y(n12551) );
  INVX1 U3195 ( .A(n12551), .Y(n1726) );
  AND2X1 U3196 ( .A(ram[1380]), .B(n10808), .Y(n12538) );
  INVX1 U3197 ( .A(n12538), .Y(n1727) );
  AND2X1 U3198 ( .A(ram[1367]), .B(n10808), .Y(n12525) );
  INVX1 U3199 ( .A(n12525), .Y(n1728) );
  AND2X1 U3200 ( .A(ram[1355]), .B(n10808), .Y(n12513) );
  INVX1 U3201 ( .A(n12513), .Y(n1729) );
  AND2X1 U3202 ( .A(ram[1341]), .B(n10806), .Y(n12497) );
  INVX1 U3203 ( .A(n12497), .Y(n1730) );
  AND2X1 U3204 ( .A(ram[1328]), .B(n10806), .Y(n12484) );
  INVX1 U3205 ( .A(n12484), .Y(n1731) );
  AND2X1 U3206 ( .A(ram[1315]), .B(n10806), .Y(n12471) );
  INVX1 U3207 ( .A(n12471), .Y(n1732) );
  AND2X1 U3208 ( .A(ram[1302]), .B(n10806), .Y(n12458) );
  INVX1 U3209 ( .A(n12458), .Y(n1733) );
  AND2X1 U3210 ( .A(ram[1290]), .B(n10806), .Y(n12446) );
  INVX1 U3211 ( .A(n12446), .Y(n1734) );
  AND2X1 U3212 ( .A(ram[1272]), .B(n10804), .Y(n12426) );
  INVX1 U3213 ( .A(n12426), .Y(n1735) );
  AND2X1 U3214 ( .A(ram[1259]), .B(n10804), .Y(n12413) );
  INVX1 U3215 ( .A(n12413), .Y(n1736) );
  AND2X1 U3216 ( .A(ram[1246]), .B(n10804), .Y(n12400) );
  INVX1 U3217 ( .A(n12400), .Y(n1737) );
  AND2X1 U3218 ( .A(ram[1233]), .B(n10804), .Y(n12387) );
  INVX1 U3219 ( .A(n12387), .Y(n1738) );
  AND2X1 U3220 ( .A(ram[1221]), .B(n10804), .Y(n12375) );
  INVX1 U3221 ( .A(n12375), .Y(n1739) );
  AND2X1 U3222 ( .A(ram[1207]), .B(n10802), .Y(n12359) );
  INVX1 U3223 ( .A(n12359), .Y(n1740) );
  AND2X1 U3224 ( .A(ram[1194]), .B(n10802), .Y(n12346) );
  INVX1 U3225 ( .A(n12346), .Y(n1741) );
  AND2X1 U3226 ( .A(ram[1181]), .B(n10802), .Y(n12333) );
  INVX1 U3227 ( .A(n12333), .Y(n1742) );
  AND2X1 U3228 ( .A(ram[1168]), .B(n10802), .Y(n12320) );
  INVX1 U3229 ( .A(n12320), .Y(n1743) );
  AND2X1 U3230 ( .A(ram[1156]), .B(n10802), .Y(n12308) );
  INVX1 U3231 ( .A(n12308), .Y(n1744) );
  AND2X1 U3232 ( .A(ram[1146]), .B(n10800), .Y(n12296) );
  INVX1 U3233 ( .A(n12296), .Y(n1745) );
  AND2X1 U3234 ( .A(ram[1133]), .B(n10800), .Y(n12283) );
  INVX1 U3235 ( .A(n12283), .Y(n1746) );
  AND2X1 U3236 ( .A(ram[1120]), .B(n10800), .Y(n12270) );
  INVX1 U3237 ( .A(n12270), .Y(n1747) );
  AND2X1 U3238 ( .A(ram[1107]), .B(n10800), .Y(n12257) );
  INVX1 U3239 ( .A(n12257), .Y(n1748) );
  AND2X1 U3240 ( .A(ram[1095]), .B(n10800), .Y(n12245) );
  INVX1 U3241 ( .A(n12245), .Y(n1749) );
  AND2X1 U3242 ( .A(ram[1081]), .B(n10798), .Y(n12229) );
  INVX1 U3243 ( .A(n12229), .Y(n1750) );
  AND2X1 U3244 ( .A(ram[1068]), .B(n10798), .Y(n12216) );
  INVX1 U3245 ( .A(n12216), .Y(n1751) );
  AND2X1 U3246 ( .A(ram[1055]), .B(n10798), .Y(n12203) );
  INVX1 U3247 ( .A(n12203), .Y(n1752) );
  AND2X1 U3248 ( .A(ram[1042]), .B(n10798), .Y(n12190) );
  INVX1 U3249 ( .A(n12190), .Y(n1753) );
  AND2X1 U3250 ( .A(ram[1030]), .B(n10798), .Y(n12178) );
  INVX1 U3251 ( .A(n12178), .Y(n1754) );
  AND2X1 U3252 ( .A(ram[1012]), .B(n10796), .Y(n12158) );
  INVX1 U3253 ( .A(n12158), .Y(n1755) );
  AND2X1 U3254 ( .A(ram[999]), .B(n10796), .Y(n12145) );
  INVX1 U3255 ( .A(n12145), .Y(n1756) );
  AND2X1 U3256 ( .A(ram[986]), .B(n10796), .Y(n12132) );
  INVX1 U3257 ( .A(n12132), .Y(n1757) );
  AND2X1 U3258 ( .A(ram[973]), .B(n10796), .Y(n12119) );
  INVX1 U3259 ( .A(n12119), .Y(n1758) );
  AND2X1 U3260 ( .A(ram[961]), .B(n10796), .Y(n12107) );
  INVX1 U3261 ( .A(n12107), .Y(n1759) );
  AND2X1 U3262 ( .A(ram[947]), .B(n10794), .Y(n12090) );
  INVX1 U3263 ( .A(n12090), .Y(n1760) );
  AND2X1 U3264 ( .A(ram[934]), .B(n10794), .Y(n12077) );
  INVX1 U3265 ( .A(n12077), .Y(n1761) );
  AND2X1 U3266 ( .A(ram[921]), .B(n10794), .Y(n12064) );
  INVX1 U3267 ( .A(n12064), .Y(n1762) );
  AND2X1 U3268 ( .A(ram[908]), .B(n10794), .Y(n12051) );
  INVX1 U3269 ( .A(n12051), .Y(n1763) );
  AND2X1 U3270 ( .A(ram[896]), .B(n10794), .Y(n12039) );
  INVX1 U3271 ( .A(n12039), .Y(n1764) );
  AND2X1 U3272 ( .A(ram[886]), .B(n10792), .Y(n12027) );
  INVX1 U3273 ( .A(n12027), .Y(n1765) );
  AND2X1 U3274 ( .A(ram[873]), .B(n10792), .Y(n12014) );
  INVX1 U3275 ( .A(n12014), .Y(n1766) );
  AND2X1 U3276 ( .A(ram[860]), .B(n10792), .Y(n12001) );
  INVX1 U3277 ( .A(n12001), .Y(n1767) );
  AND2X1 U3278 ( .A(ram[847]), .B(n10792), .Y(n11988) );
  INVX1 U3279 ( .A(n11988), .Y(n1768) );
  AND2X1 U3280 ( .A(ram[835]), .B(n10792), .Y(n11976) );
  INVX1 U3281 ( .A(n11976), .Y(n1769) );
  AND2X1 U3282 ( .A(ram[821]), .B(n10790), .Y(n11960) );
  INVX1 U3283 ( .A(n11960), .Y(n1770) );
  AND2X1 U3284 ( .A(ram[808]), .B(n10790), .Y(n11947) );
  INVX1 U3285 ( .A(n11947), .Y(n1771) );
  AND2X1 U3286 ( .A(ram[795]), .B(n10790), .Y(n11934) );
  INVX1 U3287 ( .A(n11934), .Y(n1772) );
  AND2X1 U3288 ( .A(ram[782]), .B(n10790), .Y(n11921) );
  INVX1 U3289 ( .A(n11921), .Y(n1773) );
  AND2X1 U3290 ( .A(ram[770]), .B(n10790), .Y(n11909) );
  INVX1 U3291 ( .A(n11909), .Y(n1774) );
  AND2X1 U3292 ( .A(ram[764]), .B(n10788), .Y(n11901) );
  INVX1 U3293 ( .A(n11901), .Y(n1775) );
  AND2X1 U3294 ( .A(ram[751]), .B(n10788), .Y(n11888) );
  INVX1 U3295 ( .A(n11888), .Y(n1776) );
  AND2X1 U3296 ( .A(ram[738]), .B(n10788), .Y(n11875) );
  INVX1 U3297 ( .A(n11875), .Y(n1777) );
  AND2X1 U3298 ( .A(ram[725]), .B(n10788), .Y(n11862) );
  INVX1 U3299 ( .A(n11862), .Y(n1778) );
  AND2X1 U3300 ( .A(ram[713]), .B(n10788), .Y(n11850) );
  INVX1 U3301 ( .A(n11850), .Y(n1779) );
  AND2X1 U3302 ( .A(ram[699]), .B(n10786), .Y(n11834) );
  INVX1 U3303 ( .A(n11834), .Y(n1780) );
  AND2X1 U3304 ( .A(ram[686]), .B(n10786), .Y(n11821) );
  INVX1 U3305 ( .A(n11821), .Y(n1781) );
  AND2X1 U3306 ( .A(ram[673]), .B(n10786), .Y(n11808) );
  INVX1 U3307 ( .A(n11808), .Y(n1782) );
  AND2X1 U3308 ( .A(ram[660]), .B(n10786), .Y(n11795) );
  INVX1 U3309 ( .A(n11795), .Y(n1783) );
  AND2X1 U3310 ( .A(ram[648]), .B(n10786), .Y(n11783) );
  INVX1 U3311 ( .A(n11783), .Y(n1784) );
  AND2X1 U3312 ( .A(ram[638]), .B(n10784), .Y(n11771) );
  INVX1 U3313 ( .A(n11771), .Y(n1785) );
  AND2X1 U3314 ( .A(ram[625]), .B(n10784), .Y(n11758) );
  INVX1 U3315 ( .A(n11758), .Y(n1786) );
  AND2X1 U3316 ( .A(ram[612]), .B(n10784), .Y(n11745) );
  INVX1 U3317 ( .A(n11745), .Y(n1787) );
  AND2X1 U3318 ( .A(ram[599]), .B(n10784), .Y(n11732) );
  INVX1 U3319 ( .A(n11732), .Y(n1788) );
  AND2X1 U3320 ( .A(ram[587]), .B(n10784), .Y(n11720) );
  INVX1 U3321 ( .A(n11720), .Y(n1789) );
  AND2X1 U3322 ( .A(ram[573]), .B(n10782), .Y(n11704) );
  INVX1 U3323 ( .A(n11704), .Y(n1790) );
  AND2X1 U3324 ( .A(ram[560]), .B(n10782), .Y(n11691) );
  INVX1 U3325 ( .A(n11691), .Y(n1791) );
  AND2X1 U3326 ( .A(ram[547]), .B(n10782), .Y(n11678) );
  INVX1 U3327 ( .A(n11678), .Y(n1792) );
  AND2X1 U3328 ( .A(ram[534]), .B(n10782), .Y(n11665) );
  INVX1 U3329 ( .A(n11665), .Y(n1793) );
  AND2X1 U3330 ( .A(ram[522]), .B(n10782), .Y(n11653) );
  INVX1 U3331 ( .A(n11653), .Y(n1794) );
  AND2X1 U3332 ( .A(ram[504]), .B(n10780), .Y(n11633) );
  INVX1 U3333 ( .A(n11633), .Y(n1795) );
  AND2X1 U3334 ( .A(ram[491]), .B(n10780), .Y(n11620) );
  INVX1 U3335 ( .A(n11620), .Y(n1796) );
  AND2X1 U3336 ( .A(ram[478]), .B(n10780), .Y(n11607) );
  INVX1 U3337 ( .A(n11607), .Y(n1797) );
  AND2X1 U3338 ( .A(ram[465]), .B(n10780), .Y(n11594) );
  INVX1 U3339 ( .A(n11594), .Y(n1798) );
  AND2X1 U3340 ( .A(ram[453]), .B(n10780), .Y(n11582) );
  INVX1 U3341 ( .A(n11582), .Y(n1799) );
  AND2X1 U3342 ( .A(ram[439]), .B(n10778), .Y(n11565) );
  INVX1 U3343 ( .A(n11565), .Y(n1800) );
  AND2X1 U3344 ( .A(ram[426]), .B(n10778), .Y(n11552) );
  INVX1 U3345 ( .A(n11552), .Y(n1801) );
  AND2X1 U3346 ( .A(ram[413]), .B(n10778), .Y(n11539) );
  INVX1 U3347 ( .A(n11539), .Y(n1802) );
  AND2X1 U3348 ( .A(ram[400]), .B(n10778), .Y(n11526) );
  INVX1 U3349 ( .A(n11526), .Y(n1803) );
  AND2X1 U3350 ( .A(ram[388]), .B(n10778), .Y(n11514) );
  INVX1 U3351 ( .A(n11514), .Y(n1804) );
  AND2X1 U3352 ( .A(ram[378]), .B(n10776), .Y(n11502) );
  INVX1 U3353 ( .A(n11502), .Y(n1805) );
  AND2X1 U3354 ( .A(ram[365]), .B(n10776), .Y(n11489) );
  INVX1 U3355 ( .A(n11489), .Y(n1806) );
  AND2X1 U3356 ( .A(ram[352]), .B(n10776), .Y(n11476) );
  INVX1 U3357 ( .A(n11476), .Y(n1807) );
  AND2X1 U3358 ( .A(ram[339]), .B(n10776), .Y(n11463) );
  INVX1 U3359 ( .A(n11463), .Y(n1808) );
  AND2X1 U3360 ( .A(ram[327]), .B(n10776), .Y(n11451) );
  INVX1 U3361 ( .A(n11451), .Y(n1809) );
  AND2X1 U3362 ( .A(ram[313]), .B(n10774), .Y(n11435) );
  INVX1 U3363 ( .A(n11435), .Y(n1810) );
  AND2X1 U3364 ( .A(ram[300]), .B(n10774), .Y(n11422) );
  INVX1 U3365 ( .A(n11422), .Y(n1811) );
  AND2X1 U3367 ( .A(ram[287]), .B(n10774), .Y(n11409) );
  INVX1 U3368 ( .A(n11409), .Y(n1812) );
  AND2X1 U3369 ( .A(ram[274]), .B(n10774), .Y(n11396) );
  INVX1 U3370 ( .A(n11396), .Y(n1813) );
  AND2X1 U3371 ( .A(ram[262]), .B(n10774), .Y(n11384) );
  INVX1 U3372 ( .A(n11384), .Y(n1814) );
  AND2X1 U3373 ( .A(ram[244]), .B(n10772), .Y(n11364) );
  INVX1 U3374 ( .A(n11364), .Y(n1815) );
  AND2X1 U3375 ( .A(ram[231]), .B(n10772), .Y(n11351) );
  INVX1 U3376 ( .A(n11351), .Y(n1816) );
  AND2X1 U3377 ( .A(ram[218]), .B(n10772), .Y(n11338) );
  INVX1 U3378 ( .A(n11338), .Y(n1817) );
  AND2X1 U3379 ( .A(ram[205]), .B(n10772), .Y(n11325) );
  INVX1 U3380 ( .A(n11325), .Y(n1818) );
  AND2X1 U3381 ( .A(ram[193]), .B(n10772), .Y(n11313) );
  INVX1 U3382 ( .A(n11313), .Y(n1819) );
  AND2X1 U3383 ( .A(ram[179]), .B(n10770), .Y(n11297) );
  INVX1 U3384 ( .A(n11297), .Y(n1820) );
  AND2X1 U3385 ( .A(ram[166]), .B(n10770), .Y(n11284) );
  INVX1 U3386 ( .A(n11284), .Y(n1821) );
  AND2X1 U3387 ( .A(ram[153]), .B(n10770), .Y(n11271) );
  INVX1 U3388 ( .A(n11271), .Y(n1822) );
  AND2X1 U3389 ( .A(ram[140]), .B(n10770), .Y(n11258) );
  INVX1 U3390 ( .A(n11258), .Y(n1823) );
  AND2X1 U3391 ( .A(ram[128]), .B(n10770), .Y(n11246) );
  INVX1 U3392 ( .A(n11246), .Y(n1824) );
  AND2X1 U3393 ( .A(ram[118]), .B(n10768), .Y(n11234) );
  INVX1 U3394 ( .A(n11234), .Y(n1825) );
  AND2X1 U3395 ( .A(ram[105]), .B(n10768), .Y(n11221) );
  INVX1 U3396 ( .A(n11221), .Y(n1826) );
  AND2X1 U3397 ( .A(ram[92]), .B(n10768), .Y(n11208) );
  INVX1 U3398 ( .A(n11208), .Y(n1827) );
  AND2X1 U3399 ( .A(ram[79]), .B(n10768), .Y(n11195) );
  INVX1 U3400 ( .A(n11195), .Y(n1828) );
  AND2X1 U3401 ( .A(ram[67]), .B(n10768), .Y(n11183) );
  INVX1 U3402 ( .A(n11183), .Y(n1829) );
  AND2X1 U3403 ( .A(ram[53]), .B(n10766), .Y(n11167) );
  INVX1 U3404 ( .A(n11167), .Y(n1830) );
  AND2X1 U3405 ( .A(ram[40]), .B(n10766), .Y(n11154) );
  INVX1 U3406 ( .A(n11154), .Y(n1831) );
  AND2X1 U3407 ( .A(ram[27]), .B(n10766), .Y(n11141) );
  INVX1 U3408 ( .A(n11141), .Y(n1832) );
  AND2X1 U3409 ( .A(ram[14]), .B(n10766), .Y(n11128) );
  INVX1 U3410 ( .A(n11128), .Y(n1833) );
  AND2X1 U3411 ( .A(ram[2]), .B(n10766), .Y(n11116) );
  INVX1 U3412 ( .A(n11116), .Y(n1834) );
  AND2X1 U3413 ( .A(n1993), .B(n2152), .Y(n10994) );
  INVX1 U3414 ( .A(n10994), .Y(n1835) );
  BUFX2 U3415 ( .A(n11014), .Y(n1836) );
  BUFX2 U3416 ( .A(n12633), .Y(n1837) );
  AND2X1 U3417 ( .A(ram[1978]), .B(n10952), .Y(n13214) );
  INVX1 U3418 ( .A(n13214), .Y(n1838) );
  AND2X1 U3419 ( .A(ram[1965]), .B(n10952), .Y(n13188) );
  INVX1 U3420 ( .A(n13188), .Y(n1839) );
  AND2X1 U3421 ( .A(ram[1952]), .B(n10952), .Y(n13162) );
  INVX1 U3422 ( .A(n13162), .Y(n1840) );
  AND2X1 U3423 ( .A(ram[1939]), .B(n10952), .Y(n13136) );
  INVX1 U3424 ( .A(n13136), .Y(n1841) );
  AND2X1 U3425 ( .A(ram[1927]), .B(n10952), .Y(n13112) );
  INVX1 U3426 ( .A(n13112), .Y(n1842) );
  AND2X1 U3427 ( .A(ram[1911]), .B(n10824), .Y(n13086) );
  INVX1 U3428 ( .A(n13086), .Y(n1843) );
  AND2X1 U3429 ( .A(ram[1898]), .B(n10824), .Y(n13073) );
  INVX1 U3430 ( .A(n13073), .Y(n1844) );
  AND2X1 U3431 ( .A(ram[1885]), .B(n10824), .Y(n13060) );
  INVX1 U3432 ( .A(n13060), .Y(n1845) );
  AND2X1 U3433 ( .A(ram[1872]), .B(n10824), .Y(n13047) );
  INVX1 U3434 ( .A(n13047), .Y(n1846) );
  AND2X1 U3435 ( .A(ram[1860]), .B(n10824), .Y(n13035) );
  INVX1 U3436 ( .A(n13035), .Y(n1847) );
  AND2X1 U3437 ( .A(ram[1848]), .B(n10822), .Y(n13021) );
  INVX1 U3438 ( .A(n13021), .Y(n1848) );
  AND2X1 U3439 ( .A(ram[1835]), .B(n10822), .Y(n13008) );
  INVX1 U3440 ( .A(n13008), .Y(n1849) );
  AND2X1 U3441 ( .A(ram[1822]), .B(n10822), .Y(n12995) );
  INVX1 U3442 ( .A(n12995), .Y(n1850) );
  AND2X1 U3443 ( .A(ram[1809]), .B(n10822), .Y(n12982) );
  INVX1 U3444 ( .A(n12982), .Y(n1851) );
  AND2X1 U3445 ( .A(ram[1797]), .B(n10822), .Y(n12970) );
  INVX1 U3446 ( .A(n12970), .Y(n1852) );
  AND2X1 U3447 ( .A(ram[1781]), .B(n10820), .Y(n12952) );
  INVX1 U3448 ( .A(n12952), .Y(n1853) );
  AND2X1 U3449 ( .A(ram[1768]), .B(n10820), .Y(n12939) );
  INVX1 U3450 ( .A(n12939), .Y(n1854) );
  AND2X1 U3451 ( .A(ram[1755]), .B(n10820), .Y(n12926) );
  INVX1 U3452 ( .A(n12926), .Y(n1855) );
  AND2X1 U3453 ( .A(ram[1742]), .B(n10820), .Y(n12913) );
  INVX1 U3454 ( .A(n12913), .Y(n1856) );
  AND2X1 U3455 ( .A(ram[1730]), .B(n10820), .Y(n12901) );
  INVX1 U3456 ( .A(n12901), .Y(n1857) );
  AND2X1 U3457 ( .A(ram[1718]), .B(n10818), .Y(n12887) );
  INVX1 U3458 ( .A(n12887), .Y(n1858) );
  AND2X1 U3459 ( .A(ram[1705]), .B(n10818), .Y(n12874) );
  INVX1 U3460 ( .A(n12874), .Y(n1859) );
  AND2X1 U3461 ( .A(ram[1692]), .B(n10818), .Y(n12861) );
  INVX1 U3462 ( .A(n12861), .Y(n1860) );
  AND2X1 U3463 ( .A(ram[1679]), .B(n10818), .Y(n12848) );
  INVX1 U3464 ( .A(n12848), .Y(n1861) );
  AND2X1 U3465 ( .A(ram[1667]), .B(n10818), .Y(n12836) );
  INVX1 U3466 ( .A(n12836), .Y(n1862) );
  AND2X1 U3467 ( .A(ram[1651]), .B(n10816), .Y(n12818) );
  INVX1 U3468 ( .A(n12818), .Y(n1863) );
  AND2X1 U3469 ( .A(ram[1638]), .B(n10816), .Y(n12805) );
  INVX1 U3470 ( .A(n12805), .Y(n1864) );
  AND2X1 U3471 ( .A(ram[1625]), .B(n10816), .Y(n12792) );
  INVX1 U3472 ( .A(n12792), .Y(n1865) );
  AND2X1 U3473 ( .A(ram[1612]), .B(n10816), .Y(n12779) );
  INVX1 U3474 ( .A(n12779), .Y(n1866) );
  AND2X1 U3475 ( .A(ram[1600]), .B(n10816), .Y(n12767) );
  INVX1 U3476 ( .A(n12767), .Y(n1867) );
  AND2X1 U3477 ( .A(ram[1588]), .B(n10814), .Y(n12753) );
  INVX1 U3478 ( .A(n12753), .Y(n1868) );
  AND2X1 U3479 ( .A(ram[1575]), .B(n10814), .Y(n12740) );
  INVX1 U3480 ( .A(n12740), .Y(n1869) );
  AND2X1 U3481 ( .A(ram[1562]), .B(n10814), .Y(n12727) );
  INVX1 U3482 ( .A(n12727), .Y(n1870) );
  AND2X1 U3483 ( .A(ram[1549]), .B(n10814), .Y(n12714) );
  INVX1 U3484 ( .A(n12714), .Y(n1871) );
  AND2X1 U3485 ( .A(ram[1537]), .B(n10814), .Y(n12702) );
  INVX1 U3486 ( .A(n12702), .Y(n1872) );
  AND2X1 U3487 ( .A(ram[1533]), .B(n10812), .Y(n12696) );
  INVX1 U3488 ( .A(n12696), .Y(n1873) );
  AND2X1 U3489 ( .A(ram[1520]), .B(n10812), .Y(n12683) );
  INVX1 U3490 ( .A(n12683), .Y(n1874) );
  AND2X1 U3491 ( .A(ram[1507]), .B(n10812), .Y(n12670) );
  INVX1 U3492 ( .A(n12670), .Y(n1875) );
  AND2X1 U3493 ( .A(ram[1494]), .B(n10812), .Y(n12657) );
  INVX1 U3494 ( .A(n12657), .Y(n1876) );
  AND2X1 U3495 ( .A(ram[1482]), .B(n10812), .Y(n12645) );
  INVX1 U3496 ( .A(n12645), .Y(n1877) );
  AND2X1 U3498 ( .A(ram[1470]), .B(n10810), .Y(n12630) );
  INVX1 U3499 ( .A(n12630), .Y(n1878) );
  AND2X1 U3500 ( .A(ram[1457]), .B(n10810), .Y(n12617) );
  INVX1 U3501 ( .A(n12617), .Y(n1879) );
  AND2X1 U3502 ( .A(ram[1444]), .B(n10810), .Y(n12604) );
  INVX1 U3503 ( .A(n12604), .Y(n1880) );
  AND2X1 U3504 ( .A(ram[1431]), .B(n10810), .Y(n12591) );
  INVX1 U3505 ( .A(n12591), .Y(n1881) );
  AND2X1 U3506 ( .A(ram[1419]), .B(n10810), .Y(n12579) );
  INVX1 U3507 ( .A(n12579), .Y(n1882) );
  AND2X1 U3508 ( .A(ram[1403]), .B(n10808), .Y(n12561) );
  INVX1 U3509 ( .A(n12561), .Y(n1883) );
  AND2X1 U3510 ( .A(ram[1390]), .B(n10808), .Y(n12548) );
  INVX1 U3511 ( .A(n12548), .Y(n1884) );
  AND2X1 U3512 ( .A(ram[1377]), .B(n10808), .Y(n12535) );
  INVX1 U3513 ( .A(n12535), .Y(n1885) );
  AND2X1 U3514 ( .A(ram[1364]), .B(n10808), .Y(n12522) );
  INVX1 U3515 ( .A(n12522), .Y(n1886) );
  AND2X1 U3516 ( .A(ram[1352]), .B(n10808), .Y(n12510) );
  INVX1 U3517 ( .A(n12510), .Y(n1887) );
  AND2X1 U3518 ( .A(ram[1340]), .B(n10806), .Y(n12496) );
  INVX1 U3519 ( .A(n12496), .Y(n1888) );
  AND2X1 U3520 ( .A(ram[1327]), .B(n10806), .Y(n12483) );
  INVX1 U3521 ( .A(n12483), .Y(n1889) );
  AND2X1 U3522 ( .A(ram[1314]), .B(n10806), .Y(n12470) );
  INVX1 U3523 ( .A(n12470), .Y(n1890) );
  AND2X1 U3524 ( .A(ram[1301]), .B(n10806), .Y(n12457) );
  INVX1 U3525 ( .A(n12457), .Y(n1891) );
  AND2X1 U3526 ( .A(ram[1289]), .B(n10806), .Y(n12445) );
  INVX1 U3527 ( .A(n12445), .Y(n1892) );
  AND2X1 U3528 ( .A(ram[1273]), .B(n10804), .Y(n12427) );
  INVX1 U3529 ( .A(n12427), .Y(n1893) );
  AND2X1 U3530 ( .A(ram[1260]), .B(n10804), .Y(n12414) );
  INVX1 U3531 ( .A(n12414), .Y(n1894) );
  AND2X1 U3532 ( .A(ram[1247]), .B(n10804), .Y(n12401) );
  INVX1 U3533 ( .A(n12401), .Y(n1895) );
  AND2X1 U3534 ( .A(ram[1234]), .B(n10804), .Y(n12388) );
  INVX1 U3535 ( .A(n12388), .Y(n1896) );
  AND2X1 U3536 ( .A(ram[1222]), .B(n10804), .Y(n12376) );
  INVX1 U3537 ( .A(n12376), .Y(n1897) );
  AND2X1 U3538 ( .A(ram[1210]), .B(n10802), .Y(n12362) );
  INVX1 U3539 ( .A(n12362), .Y(n1898) );
  AND2X1 U3540 ( .A(ram[1197]), .B(n10802), .Y(n12349) );
  INVX1 U3541 ( .A(n12349), .Y(n1899) );
  AND2X1 U3542 ( .A(ram[1184]), .B(n10802), .Y(n12336) );
  INVX1 U3543 ( .A(n12336), .Y(n1900) );
  AND2X1 U3544 ( .A(ram[1171]), .B(n10802), .Y(n12323) );
  INVX1 U3545 ( .A(n12323), .Y(n1901) );
  AND2X1 U3546 ( .A(ram[1159]), .B(n10802), .Y(n12311) );
  INVX1 U3547 ( .A(n12311), .Y(n1902) );
  AND2X1 U3548 ( .A(ram[1143]), .B(n10800), .Y(n12293) );
  INVX1 U3549 ( .A(n12293), .Y(n1903) );
  AND2X1 U3550 ( .A(ram[1130]), .B(n10800), .Y(n12280) );
  INVX1 U3551 ( .A(n12280), .Y(n1904) );
  AND2X1 U3552 ( .A(ram[1117]), .B(n10800), .Y(n12267) );
  INVX1 U3553 ( .A(n12267), .Y(n1905) );
  AND2X1 U3554 ( .A(ram[1104]), .B(n10800), .Y(n12254) );
  INVX1 U3555 ( .A(n12254), .Y(n1906) );
  AND2X1 U3556 ( .A(ram[1092]), .B(n10800), .Y(n12242) );
  INVX1 U3557 ( .A(n12242), .Y(n1907) );
  AND2X1 U3558 ( .A(ram[1080]), .B(n10798), .Y(n12228) );
  INVX1 U3559 ( .A(n12228), .Y(n1908) );
  AND2X1 U3560 ( .A(ram[1067]), .B(n10798), .Y(n12215) );
  INVX1 U3561 ( .A(n12215), .Y(n1909) );
  AND2X1 U3562 ( .A(ram[1054]), .B(n10798), .Y(n12202) );
  INVX1 U3563 ( .A(n12202), .Y(n1910) );
  AND2X1 U3564 ( .A(ram[1041]), .B(n10798), .Y(n12189) );
  INVX1 U3565 ( .A(n12189), .Y(n1911) );
  AND2X1 U3566 ( .A(ram[1029]), .B(n10798), .Y(n12177) );
  INVX1 U3567 ( .A(n12177), .Y(n1912) );
  AND2X1 U3568 ( .A(ram[1013]), .B(n10796), .Y(n12159) );
  INVX1 U3569 ( .A(n12159), .Y(n1913) );
  AND2X1 U3570 ( .A(ram[1000]), .B(n10796), .Y(n12146) );
  INVX1 U3571 ( .A(n12146), .Y(n1914) );
  AND2X1 U3572 ( .A(ram[987]), .B(n10796), .Y(n12133) );
  INVX1 U3573 ( .A(n12133), .Y(n1915) );
  AND2X1 U3574 ( .A(ram[974]), .B(n10796), .Y(n12120) );
  INVX1 U3575 ( .A(n12120), .Y(n1916) );
  AND2X1 U3576 ( .A(ram[962]), .B(n10796), .Y(n12108) );
  INVX1 U3577 ( .A(n12108), .Y(n1917) );
  AND2X1 U3578 ( .A(ram[950]), .B(n10794), .Y(n12093) );
  INVX1 U3579 ( .A(n12093), .Y(n1918) );
  AND2X1 U3580 ( .A(ram[937]), .B(n10794), .Y(n12080) );
  INVX1 U3581 ( .A(n12080), .Y(n1919) );
  AND2X1 U3582 ( .A(ram[924]), .B(n10794), .Y(n12067) );
  INVX1 U3583 ( .A(n12067), .Y(n1920) );
  AND2X1 U3584 ( .A(ram[911]), .B(n10794), .Y(n12054) );
  INVX1 U3585 ( .A(n12054), .Y(n1921) );
  AND2X1 U3586 ( .A(ram[899]), .B(n10794), .Y(n12042) );
  INVX1 U3587 ( .A(n12042), .Y(n1922) );
  AND2X1 U3588 ( .A(ram[883]), .B(n10792), .Y(n12024) );
  INVX1 U3589 ( .A(n12024), .Y(n1923) );
  AND2X1 U3590 ( .A(ram[870]), .B(n10792), .Y(n12011) );
  INVX1 U3591 ( .A(n12011), .Y(n1924) );
  AND2X1 U3592 ( .A(ram[857]), .B(n10792), .Y(n11998) );
  INVX1 U3593 ( .A(n11998), .Y(n1925) );
  AND2X1 U3594 ( .A(ram[844]), .B(n10792), .Y(n11985) );
  INVX1 U3595 ( .A(n11985), .Y(n1926) );
  AND2X1 U3596 ( .A(ram[832]), .B(n10792), .Y(n11973) );
  INVX1 U3597 ( .A(n11973), .Y(n1927) );
  AND2X1 U3598 ( .A(ram[820]), .B(n10790), .Y(n11959) );
  INVX1 U3599 ( .A(n11959), .Y(n1928) );
  AND2X1 U3600 ( .A(ram[807]), .B(n10790), .Y(n11946) );
  INVX1 U3601 ( .A(n11946), .Y(n1929) );
  AND2X1 U3602 ( .A(ram[794]), .B(n10790), .Y(n11933) );
  INVX1 U3603 ( .A(n11933), .Y(n1930) );
  AND2X1 U3604 ( .A(ram[781]), .B(n10790), .Y(n11920) );
  INVX1 U3605 ( .A(n11920), .Y(n1931) );
  AND2X1 U3606 ( .A(ram[769]), .B(n10790), .Y(n11908) );
  INVX1 U3607 ( .A(n11908), .Y(n1932) );
  AND2X1 U3608 ( .A(ram[765]), .B(n10788), .Y(n11902) );
  INVX1 U3609 ( .A(n11902), .Y(n1933) );
  AND2X1 U3610 ( .A(ram[752]), .B(n10788), .Y(n11889) );
  INVX1 U3611 ( .A(n11889), .Y(n1934) );
  AND2X1 U3612 ( .A(ram[739]), .B(n10788), .Y(n11876) );
  INVX1 U3613 ( .A(n11876), .Y(n1935) );
  AND2X1 U3614 ( .A(ram[726]), .B(n10788), .Y(n11863) );
  INVX1 U3615 ( .A(n11863), .Y(n1936) );
  AND2X1 U3616 ( .A(ram[714]), .B(n10788), .Y(n11851) );
  INVX1 U3617 ( .A(n11851), .Y(n1937) );
  AND2X1 U3618 ( .A(ram[702]), .B(n10786), .Y(n11837) );
  INVX1 U3619 ( .A(n11837), .Y(n1938) );
  AND2X1 U3620 ( .A(ram[689]), .B(n10786), .Y(n11824) );
  INVX1 U3621 ( .A(n11824), .Y(n1939) );
  AND2X1 U3622 ( .A(ram[676]), .B(n10786), .Y(n11811) );
  INVX1 U3623 ( .A(n11811), .Y(n1940) );
  AND2X1 U3624 ( .A(ram[663]), .B(n10786), .Y(n11798) );
  INVX1 U3625 ( .A(n11798), .Y(n1941) );
  AND2X1 U3626 ( .A(ram[651]), .B(n10786), .Y(n11786) );
  INVX1 U3627 ( .A(n11786), .Y(n1942) );
  AND2X1 U3629 ( .A(ram[635]), .B(n10784), .Y(n11768) );
  INVX1 U3630 ( .A(n11768), .Y(n1943) );
  AND2X1 U3631 ( .A(ram[622]), .B(n10784), .Y(n11755) );
  INVX1 U3632 ( .A(n11755), .Y(n1944) );
  AND2X1 U3633 ( .A(ram[609]), .B(n10784), .Y(n11742) );
  INVX1 U3634 ( .A(n11742), .Y(n1945) );
  AND2X1 U3635 ( .A(ram[596]), .B(n10784), .Y(n11729) );
  INVX1 U3636 ( .A(n11729), .Y(n1946) );
  AND2X1 U3637 ( .A(ram[584]), .B(n10784), .Y(n11717) );
  INVX1 U3638 ( .A(n11717), .Y(n1947) );
  AND2X1 U3639 ( .A(ram[572]), .B(n10782), .Y(n11703) );
  INVX1 U3640 ( .A(n11703), .Y(n1948) );
  AND2X1 U3641 ( .A(ram[559]), .B(n10782), .Y(n11690) );
  INVX1 U3642 ( .A(n11690), .Y(n1949) );
  AND2X1 U3643 ( .A(ram[546]), .B(n10782), .Y(n11677) );
  INVX1 U3644 ( .A(n11677), .Y(n1950) );
  AND2X1 U3645 ( .A(ram[533]), .B(n10782), .Y(n11664) );
  INVX1 U3646 ( .A(n11664), .Y(n1951) );
  AND2X1 U3647 ( .A(ram[521]), .B(n10782), .Y(n11652) );
  INVX1 U3648 ( .A(n11652), .Y(n1952) );
  AND2X1 U3649 ( .A(ram[505]), .B(n10780), .Y(n11634) );
  INVX1 U3650 ( .A(n11634), .Y(n1953) );
  AND2X1 U3651 ( .A(ram[492]), .B(n10780), .Y(n11621) );
  INVX1 U3652 ( .A(n11621), .Y(n1954) );
  AND2X1 U3653 ( .A(ram[479]), .B(n10780), .Y(n11608) );
  INVX1 U3654 ( .A(n11608), .Y(n1955) );
  AND2X1 U3655 ( .A(ram[466]), .B(n10780), .Y(n11595) );
  INVX1 U3656 ( .A(n11595), .Y(n1956) );
  AND2X1 U3657 ( .A(ram[454]), .B(n10780), .Y(n11583) );
  INVX1 U3658 ( .A(n11583), .Y(n1957) );
  AND2X1 U3659 ( .A(ram[442]), .B(n10778), .Y(n11568) );
  INVX1 U3660 ( .A(n11568), .Y(n1958) );
  AND2X1 U3661 ( .A(ram[429]), .B(n10778), .Y(n11555) );
  INVX1 U3662 ( .A(n11555), .Y(n1959) );
  AND2X1 U3663 ( .A(ram[416]), .B(n10778), .Y(n11542) );
  INVX1 U3664 ( .A(n11542), .Y(n1960) );
  AND2X1 U3665 ( .A(ram[403]), .B(n10778), .Y(n11529) );
  INVX1 U3666 ( .A(n11529), .Y(n1961) );
  AND2X1 U3667 ( .A(ram[391]), .B(n10778), .Y(n11517) );
  INVX1 U3668 ( .A(n11517), .Y(n1962) );
  AND2X1 U3669 ( .A(ram[375]), .B(n10776), .Y(n11499) );
  INVX1 U3670 ( .A(n11499), .Y(n1963) );
  AND2X1 U3671 ( .A(ram[362]), .B(n10776), .Y(n11486) );
  INVX1 U3672 ( .A(n11486), .Y(n1964) );
  AND2X1 U3673 ( .A(ram[349]), .B(n10776), .Y(n11473) );
  INVX1 U3674 ( .A(n11473), .Y(n1965) );
  AND2X1 U3675 ( .A(ram[336]), .B(n10776), .Y(n11460) );
  INVX1 U3676 ( .A(n11460), .Y(n1966) );
  AND2X1 U3677 ( .A(ram[324]), .B(n10776), .Y(n11448) );
  INVX1 U3678 ( .A(n11448), .Y(n1967) );
  AND2X1 U3679 ( .A(ram[312]), .B(n10774), .Y(n11434) );
  INVX1 U3680 ( .A(n11434), .Y(n1968) );
  AND2X1 U3681 ( .A(ram[299]), .B(n10774), .Y(n11421) );
  INVX1 U3682 ( .A(n11421), .Y(n1969) );
  AND2X1 U3683 ( .A(ram[286]), .B(n10774), .Y(n11408) );
  INVX1 U3684 ( .A(n11408), .Y(n1970) );
  AND2X1 U3685 ( .A(ram[273]), .B(n10774), .Y(n11395) );
  INVX1 U3686 ( .A(n11395), .Y(n1971) );
  AND2X1 U3687 ( .A(ram[261]), .B(n10774), .Y(n11383) );
  INVX1 U3688 ( .A(n11383), .Y(n1972) );
  AND2X1 U3689 ( .A(ram[245]), .B(n10772), .Y(n11365) );
  INVX1 U3690 ( .A(n11365), .Y(n1973) );
  AND2X1 U3691 ( .A(ram[232]), .B(n10772), .Y(n11352) );
  INVX1 U3692 ( .A(n11352), .Y(n1974) );
  AND2X1 U3693 ( .A(ram[219]), .B(n10772), .Y(n11339) );
  INVX1 U3694 ( .A(n11339), .Y(n1975) );
  AND2X1 U3695 ( .A(ram[206]), .B(n10772), .Y(n11326) );
  INVX1 U3696 ( .A(n11326), .Y(n1976) );
  AND2X1 U3697 ( .A(ram[194]), .B(n10772), .Y(n11314) );
  INVX1 U3698 ( .A(n11314), .Y(n1977) );
  AND2X1 U3699 ( .A(ram[182]), .B(n10770), .Y(n11300) );
  INVX1 U3700 ( .A(n11300), .Y(n1978) );
  AND2X1 U3701 ( .A(ram[169]), .B(n10770), .Y(n11287) );
  INVX1 U3702 ( .A(n11287), .Y(n1979) );
  AND2X1 U3703 ( .A(ram[156]), .B(n10770), .Y(n11274) );
  INVX1 U3704 ( .A(n11274), .Y(n1980) );
  AND2X1 U3705 ( .A(ram[143]), .B(n10770), .Y(n11261) );
  INVX1 U3706 ( .A(n11261), .Y(n1981) );
  AND2X1 U3707 ( .A(ram[131]), .B(n10770), .Y(n11249) );
  INVX1 U3708 ( .A(n11249), .Y(n1982) );
  AND2X1 U3709 ( .A(ram[115]), .B(n10768), .Y(n11231) );
  INVX1 U3710 ( .A(n11231), .Y(n1983) );
  AND2X1 U3711 ( .A(ram[102]), .B(n10768), .Y(n11218) );
  INVX1 U3712 ( .A(n11218), .Y(n1984) );
  AND2X1 U3713 ( .A(ram[89]), .B(n10768), .Y(n11205) );
  INVX1 U3714 ( .A(n11205), .Y(n1985) );
  AND2X1 U3715 ( .A(ram[76]), .B(n10768), .Y(n11192) );
  INVX1 U3716 ( .A(n11192), .Y(n1986) );
  AND2X1 U3717 ( .A(ram[64]), .B(n10768), .Y(n11180) );
  INVX1 U3718 ( .A(n11180), .Y(n1987) );
  AND2X1 U3719 ( .A(ram[52]), .B(n10766), .Y(n11166) );
  INVX1 U3720 ( .A(n11166), .Y(n1988) );
  AND2X1 U3721 ( .A(ram[39]), .B(n10766), .Y(n11153) );
  INVX1 U3722 ( .A(n11153), .Y(n1989) );
  AND2X1 U3723 ( .A(ram[26]), .B(n10766), .Y(n11140) );
  INVX1 U3724 ( .A(n11140), .Y(n1990) );
  AND2X1 U3725 ( .A(ram[13]), .B(n10766), .Y(n11127) );
  INVX1 U3726 ( .A(n11127), .Y(n1991) );
  AND2X1 U3727 ( .A(ram[1]), .B(n10766), .Y(n11115) );
  INVX1 U3728 ( .A(n11115), .Y(n1992) );
  AND2X1 U3729 ( .A(n13228), .B(n13227), .Y(n4668) );
  INVX1 U3730 ( .A(n4668), .Y(n1993) );
  BUFX2 U3731 ( .A(n12104), .Y(n1994) );
  AND2X1 U3732 ( .A(ram[1977]), .B(n10952), .Y(n13212) );
  INVX1 U3733 ( .A(n13212), .Y(n1995) );
  AND2X1 U3734 ( .A(ram[1964]), .B(n10952), .Y(n13186) );
  INVX1 U3735 ( .A(n13186), .Y(n1996) );
  AND2X1 U3736 ( .A(ram[1951]), .B(n10952), .Y(n13160) );
  INVX1 U3737 ( .A(n13160), .Y(n1997) );
  AND2X1 U3738 ( .A(ram[1938]), .B(n10952), .Y(n13134) );
  INVX1 U3739 ( .A(n13134), .Y(n1998) );
  AND2X1 U3740 ( .A(ram[1926]), .B(n10952), .Y(n13110) );
  INVX1 U3741 ( .A(n13110), .Y(n1999) );
  AND2X1 U3742 ( .A(ram[1912]), .B(n10824), .Y(n13087) );
  INVX1 U3743 ( .A(n13087), .Y(n2000) );
  AND2X1 U3744 ( .A(ram[1899]), .B(n10824), .Y(n13074) );
  INVX1 U3745 ( .A(n13074), .Y(n2001) );
  AND2X1 U3746 ( .A(ram[1886]), .B(n10824), .Y(n13061) );
  INVX1 U3747 ( .A(n13061), .Y(n2002) );
  AND2X1 U3748 ( .A(ram[1873]), .B(n10824), .Y(n13048) );
  INVX1 U3749 ( .A(n13048), .Y(n2003) );
  AND2X1 U3750 ( .A(ram[1861]), .B(n10824), .Y(n13036) );
  INVX1 U3751 ( .A(n13036), .Y(n2004) );
  AND2X1 U3752 ( .A(ram[1847]), .B(n10822), .Y(n13020) );
  INVX1 U3753 ( .A(n13020), .Y(n2005) );
  AND2X1 U3754 ( .A(ram[1834]), .B(n10822), .Y(n13007) );
  INVX1 U3755 ( .A(n13007), .Y(n2006) );
  AND2X1 U3756 ( .A(ram[1821]), .B(n10822), .Y(n12994) );
  INVX1 U3757 ( .A(n12994), .Y(n2007) );
  AND2X1 U3758 ( .A(ram[1808]), .B(n10822), .Y(n12981) );
  INVX1 U3760 ( .A(n12981), .Y(n2008) );
  AND2X1 U3761 ( .A(ram[1796]), .B(n10822), .Y(n12969) );
  INVX1 U3762 ( .A(n12969), .Y(n2009) );
  AND2X1 U3763 ( .A(ram[1782]), .B(n10820), .Y(n12953) );
  INVX1 U3764 ( .A(n12953), .Y(n2010) );
  AND2X1 U3765 ( .A(ram[1769]), .B(n10820), .Y(n12940) );
  INVX1 U3766 ( .A(n12940), .Y(n2011) );
  AND2X1 U3767 ( .A(ram[1756]), .B(n10820), .Y(n12927) );
  INVX1 U3768 ( .A(n12927), .Y(n2012) );
  AND2X1 U3769 ( .A(ram[1743]), .B(n10820), .Y(n12914) );
  INVX1 U3770 ( .A(n12914), .Y(n2013) );
  AND2X1 U3771 ( .A(ram[1731]), .B(n10820), .Y(n12902) );
  INVX1 U3772 ( .A(n12902), .Y(n2014) );
  AND2X1 U3773 ( .A(ram[1717]), .B(n10818), .Y(n12886) );
  INVX1 U3774 ( .A(n12886), .Y(n2015) );
  AND2X1 U3775 ( .A(ram[1704]), .B(n10818), .Y(n12873) );
  INVX1 U3776 ( .A(n12873), .Y(n2016) );
  AND2X1 U3777 ( .A(ram[1691]), .B(n10818), .Y(n12860) );
  INVX1 U3778 ( .A(n12860), .Y(n2017) );
  AND2X1 U3779 ( .A(ram[1678]), .B(n10818), .Y(n12847) );
  INVX1 U3780 ( .A(n12847), .Y(n2018) );
  AND2X1 U3781 ( .A(ram[1666]), .B(n10818), .Y(n12835) );
  INVX1 U3782 ( .A(n12835), .Y(n2019) );
  AND2X1 U3783 ( .A(ram[1652]), .B(n10816), .Y(n12819) );
  INVX1 U3784 ( .A(n12819), .Y(n2020) );
  AND2X1 U3785 ( .A(ram[1639]), .B(n10816), .Y(n12806) );
  INVX1 U3786 ( .A(n12806), .Y(n2021) );
  AND2X1 U3787 ( .A(ram[1626]), .B(n10816), .Y(n12793) );
  INVX1 U3788 ( .A(n12793), .Y(n2022) );
  AND2X1 U3789 ( .A(ram[1613]), .B(n10816), .Y(n12780) );
  INVX1 U3790 ( .A(n12780), .Y(n2023) );
  AND2X1 U3791 ( .A(ram[1601]), .B(n10816), .Y(n12768) );
  INVX1 U3792 ( .A(n12768), .Y(n2024) );
  AND2X1 U3793 ( .A(ram[1587]), .B(n10814), .Y(n12752) );
  INVX1 U3794 ( .A(n12752), .Y(n2025) );
  AND2X1 U3795 ( .A(ram[1574]), .B(n10814), .Y(n12739) );
  INVX1 U3796 ( .A(n12739), .Y(n2026) );
  AND2X1 U3797 ( .A(ram[1561]), .B(n10814), .Y(n12726) );
  INVX1 U3798 ( .A(n12726), .Y(n2027) );
  AND2X1 U3799 ( .A(ram[1548]), .B(n10814), .Y(n12713) );
  INVX1 U3800 ( .A(n12713), .Y(n2028) );
  AND2X1 U3801 ( .A(ram[1536]), .B(n10814), .Y(n12701) );
  INVX1 U3802 ( .A(n12701), .Y(n2029) );
  AND2X1 U3803 ( .A(ram[1534]), .B(n10812), .Y(n12697) );
  INVX1 U3804 ( .A(n12697), .Y(n2030) );
  AND2X1 U3805 ( .A(ram[1521]), .B(n10812), .Y(n12684) );
  INVX1 U3806 ( .A(n12684), .Y(n2031) );
  AND2X1 U3807 ( .A(ram[1508]), .B(n10812), .Y(n12671) );
  INVX1 U3808 ( .A(n12671), .Y(n2032) );
  AND2X1 U3809 ( .A(ram[1495]), .B(n10812), .Y(n12658) );
  INVX1 U3810 ( .A(n12658), .Y(n2033) );
  AND2X1 U3811 ( .A(ram[1483]), .B(n10812), .Y(n12646) );
  INVX1 U3812 ( .A(n12646), .Y(n2034) );
  AND2X1 U3813 ( .A(ram[1469]), .B(n10810), .Y(n12629) );
  INVX1 U3814 ( .A(n12629), .Y(n2035) );
  AND2X1 U3815 ( .A(ram[1456]), .B(n10810), .Y(n12616) );
  INVX1 U3816 ( .A(n12616), .Y(n2036) );
  AND2X1 U3817 ( .A(ram[1443]), .B(n10810), .Y(n12603) );
  INVX1 U3818 ( .A(n12603), .Y(n2037) );
  AND2X1 U3819 ( .A(ram[1430]), .B(n10810), .Y(n12590) );
  INVX1 U3820 ( .A(n12590), .Y(n2038) );
  AND2X1 U3821 ( .A(ram[1418]), .B(n10810), .Y(n12578) );
  INVX1 U3822 ( .A(n12578), .Y(n2039) );
  AND2X1 U3823 ( .A(ram[1404]), .B(n10808), .Y(n12562) );
  INVX1 U3824 ( .A(n12562), .Y(n2040) );
  AND2X1 U3825 ( .A(ram[1391]), .B(n10808), .Y(n12549) );
  INVX1 U3826 ( .A(n12549), .Y(n2041) );
  AND2X1 U3827 ( .A(ram[1378]), .B(n10808), .Y(n12536) );
  INVX1 U3828 ( .A(n12536), .Y(n2042) );
  AND2X1 U3829 ( .A(ram[1365]), .B(n10808), .Y(n12523) );
  INVX1 U3830 ( .A(n12523), .Y(n2043) );
  AND2X1 U3831 ( .A(ram[1353]), .B(n10808), .Y(n12511) );
  INVX1 U3832 ( .A(n12511), .Y(n2044) );
  AND2X1 U3833 ( .A(ram[1339]), .B(n10806), .Y(n12495) );
  INVX1 U3834 ( .A(n12495), .Y(n2045) );
  AND2X1 U3835 ( .A(ram[1326]), .B(n10806), .Y(n12482) );
  INVX1 U3836 ( .A(n12482), .Y(n2046) );
  AND2X1 U3837 ( .A(ram[1313]), .B(n10806), .Y(n12469) );
  INVX1 U3838 ( .A(n12469), .Y(n2047) );
  AND2X1 U3839 ( .A(ram[1300]), .B(n10806), .Y(n12456) );
  INVX1 U3840 ( .A(n12456), .Y(n2048) );
  AND2X1 U3841 ( .A(ram[1288]), .B(n10806), .Y(n12444) );
  INVX1 U3842 ( .A(n12444), .Y(n2049) );
  AND2X1 U3843 ( .A(ram[1274]), .B(n10804), .Y(n12428) );
  INVX1 U3844 ( .A(n12428), .Y(n2050) );
  AND2X1 U3845 ( .A(ram[1261]), .B(n10804), .Y(n12415) );
  INVX1 U3846 ( .A(n12415), .Y(n2051) );
  AND2X1 U3847 ( .A(ram[1248]), .B(n10804), .Y(n12402) );
  INVX1 U3848 ( .A(n12402), .Y(n2052) );
  AND2X1 U3849 ( .A(ram[1235]), .B(n10804), .Y(n12389) );
  INVX1 U3850 ( .A(n12389), .Y(n2053) );
  AND2X1 U3851 ( .A(ram[1223]), .B(n10804), .Y(n12377) );
  INVX1 U3852 ( .A(n12377), .Y(n2054) );
  AND2X1 U3853 ( .A(ram[1209]), .B(n10802), .Y(n12361) );
  INVX1 U3854 ( .A(n12361), .Y(n2055) );
  AND2X1 U3855 ( .A(ram[1196]), .B(n10802), .Y(n12348) );
  INVX1 U3856 ( .A(n12348), .Y(n2056) );
  AND2X1 U3857 ( .A(ram[1183]), .B(n10802), .Y(n12335) );
  INVX1 U3858 ( .A(n12335), .Y(n2057) );
  AND2X1 U3859 ( .A(ram[1170]), .B(n10802), .Y(n12322) );
  INVX1 U3860 ( .A(n12322), .Y(n2058) );
  AND2X1 U3861 ( .A(ram[1158]), .B(n10802), .Y(n12310) );
  INVX1 U3862 ( .A(n12310), .Y(n2059) );
  AND2X1 U3863 ( .A(ram[1144]), .B(n10800), .Y(n12294) );
  INVX1 U3864 ( .A(n12294), .Y(n2060) );
  AND2X1 U3865 ( .A(ram[1131]), .B(n10800), .Y(n12281) );
  INVX1 U3866 ( .A(n12281), .Y(n2061) );
  AND2X1 U3867 ( .A(ram[1118]), .B(n10800), .Y(n12268) );
  INVX1 U3868 ( .A(n12268), .Y(n2062) );
  AND2X1 U3869 ( .A(ram[1105]), .B(n10800), .Y(n12255) );
  INVX1 U3870 ( .A(n12255), .Y(n2063) );
  AND2X1 U3871 ( .A(ram[1093]), .B(n10800), .Y(n12243) );
  INVX1 U3872 ( .A(n12243), .Y(n2064) );
  AND2X1 U3873 ( .A(ram[1079]), .B(n10798), .Y(n12227) );
  INVX1 U3874 ( .A(n12227), .Y(n2065) );
  AND2X1 U3875 ( .A(ram[1066]), .B(n10798), .Y(n12214) );
  INVX1 U3876 ( .A(n12214), .Y(n2066) );
  AND2X1 U3877 ( .A(ram[1053]), .B(n10798), .Y(n12201) );
  INVX1 U3878 ( .A(n12201), .Y(n2067) );
  AND2X1 U3879 ( .A(ram[1040]), .B(n10798), .Y(n12188) );
  INVX1 U3880 ( .A(n12188), .Y(n2068) );
  AND2X1 U3881 ( .A(ram[1028]), .B(n10798), .Y(n12176) );
  INVX1 U3882 ( .A(n12176), .Y(n2069) );
  AND2X1 U3883 ( .A(ram[1014]), .B(n10796), .Y(n12160) );
  INVX1 U3884 ( .A(n12160), .Y(n2070) );
  AND2X1 U3885 ( .A(ram[1001]), .B(n10796), .Y(n12147) );
  INVX1 U3886 ( .A(n12147), .Y(n2071) );
  AND2X1 U3887 ( .A(ram[988]), .B(n10796), .Y(n12134) );
  INVX1 U3888 ( .A(n12134), .Y(n2072) );
  AND2X1 U3889 ( .A(ram[975]), .B(n10796), .Y(n12121) );
  INVX1 U3891 ( .A(n12121), .Y(n2073) );
  AND2X1 U3892 ( .A(ram[963]), .B(n10796), .Y(n12109) );
  INVX1 U3893 ( .A(n12109), .Y(n2074) );
  AND2X1 U3894 ( .A(ram[949]), .B(n10794), .Y(n12092) );
  INVX1 U3895 ( .A(n12092), .Y(n2075) );
  AND2X1 U3896 ( .A(ram[936]), .B(n10794), .Y(n12079) );
  INVX1 U3897 ( .A(n12079), .Y(n2076) );
  AND2X1 U3898 ( .A(ram[923]), .B(n10794), .Y(n12066) );
  INVX1 U3899 ( .A(n12066), .Y(n2077) );
  AND2X1 U3900 ( .A(ram[910]), .B(n10794), .Y(n12053) );
  INVX1 U3901 ( .A(n12053), .Y(n2078) );
  AND2X1 U3902 ( .A(ram[898]), .B(n10794), .Y(n12041) );
  INVX1 U3903 ( .A(n12041), .Y(n2079) );
  AND2X1 U3904 ( .A(ram[884]), .B(n10792), .Y(n12025) );
  INVX1 U3905 ( .A(n12025), .Y(n2080) );
  AND2X1 U3906 ( .A(ram[871]), .B(n10792), .Y(n12012) );
  INVX1 U3907 ( .A(n12012), .Y(n2081) );
  AND2X1 U3908 ( .A(ram[858]), .B(n10792), .Y(n11999) );
  INVX1 U3909 ( .A(n11999), .Y(n2082) );
  AND2X1 U3910 ( .A(ram[845]), .B(n10792), .Y(n11986) );
  INVX1 U3911 ( .A(n11986), .Y(n2083) );
  AND2X1 U3912 ( .A(ram[833]), .B(n10792), .Y(n11974) );
  INVX1 U3913 ( .A(n11974), .Y(n2084) );
  AND2X1 U3914 ( .A(ram[819]), .B(n10790), .Y(n11958) );
  INVX1 U3915 ( .A(n11958), .Y(n2085) );
  AND2X1 U3916 ( .A(ram[806]), .B(n10790), .Y(n11945) );
  INVX1 U3917 ( .A(n11945), .Y(n2086) );
  AND2X1 U3918 ( .A(ram[793]), .B(n10790), .Y(n11932) );
  INVX1 U3919 ( .A(n11932), .Y(n2087) );
  AND2X1 U3920 ( .A(ram[780]), .B(n10790), .Y(n11919) );
  INVX1 U3921 ( .A(n11919), .Y(n2088) );
  AND2X1 U3922 ( .A(ram[768]), .B(n10790), .Y(n11907) );
  INVX1 U3923 ( .A(n11907), .Y(n2089) );
  AND2X1 U3924 ( .A(ram[766]), .B(n10788), .Y(n11903) );
  INVX1 U3925 ( .A(n11903), .Y(n2090) );
  AND2X1 U3926 ( .A(ram[753]), .B(n10788), .Y(n11890) );
  INVX1 U3927 ( .A(n11890), .Y(n2091) );
  AND2X1 U3928 ( .A(ram[740]), .B(n10788), .Y(n11877) );
  INVX1 U3929 ( .A(n11877), .Y(n2092) );
  AND2X1 U3930 ( .A(ram[727]), .B(n10788), .Y(n11864) );
  INVX1 U3931 ( .A(n11864), .Y(n2093) );
  AND2X1 U3932 ( .A(ram[715]), .B(n10788), .Y(n11852) );
  INVX1 U3933 ( .A(n11852), .Y(n2094) );
  AND2X1 U3934 ( .A(ram[701]), .B(n10786), .Y(n11836) );
  INVX1 U3935 ( .A(n11836), .Y(n2095) );
  AND2X1 U3936 ( .A(ram[688]), .B(n10786), .Y(n11823) );
  INVX1 U3937 ( .A(n11823), .Y(n2096) );
  AND2X1 U3938 ( .A(ram[675]), .B(n10786), .Y(n11810) );
  INVX1 U3939 ( .A(n11810), .Y(n2097) );
  AND2X1 U3940 ( .A(ram[662]), .B(n10786), .Y(n11797) );
  INVX1 U3941 ( .A(n11797), .Y(n2098) );
  AND2X1 U3942 ( .A(ram[650]), .B(n10786), .Y(n11785) );
  INVX1 U3943 ( .A(n11785), .Y(n2099) );
  AND2X1 U3944 ( .A(ram[636]), .B(n10784), .Y(n11769) );
  INVX1 U3945 ( .A(n11769), .Y(n2100) );
  AND2X1 U3946 ( .A(ram[623]), .B(n10784), .Y(n11756) );
  INVX1 U3947 ( .A(n11756), .Y(n2101) );
  AND2X1 U3948 ( .A(ram[610]), .B(n10784), .Y(n11743) );
  INVX1 U3949 ( .A(n11743), .Y(n2102) );
  AND2X1 U3950 ( .A(ram[597]), .B(n10784), .Y(n11730) );
  INVX1 U3951 ( .A(n11730), .Y(n2103) );
  AND2X1 U3952 ( .A(ram[585]), .B(n10784), .Y(n11718) );
  INVX1 U3953 ( .A(n11718), .Y(n2104) );
  AND2X1 U3954 ( .A(ram[571]), .B(n10782), .Y(n11702) );
  INVX1 U3955 ( .A(n11702), .Y(n2105) );
  AND2X1 U3956 ( .A(ram[558]), .B(n10782), .Y(n11689) );
  INVX1 U3957 ( .A(n11689), .Y(n2106) );
  AND2X1 U3958 ( .A(ram[545]), .B(n10782), .Y(n11676) );
  INVX1 U3959 ( .A(n11676), .Y(n2107) );
  AND2X1 U3960 ( .A(ram[532]), .B(n10782), .Y(n11663) );
  INVX1 U3961 ( .A(n11663), .Y(n2108) );
  AND2X1 U3962 ( .A(ram[520]), .B(n10782), .Y(n11651) );
  INVX1 U3963 ( .A(n11651), .Y(n2109) );
  AND2X1 U3964 ( .A(ram[506]), .B(n10780), .Y(n11635) );
  INVX1 U3965 ( .A(n11635), .Y(n2110) );
  AND2X1 U3966 ( .A(ram[493]), .B(n10780), .Y(n11622) );
  INVX1 U3967 ( .A(n11622), .Y(n2111) );
  AND2X1 U3968 ( .A(ram[480]), .B(n10780), .Y(n11609) );
  INVX1 U3969 ( .A(n11609), .Y(n2112) );
  AND2X1 U3970 ( .A(ram[467]), .B(n10780), .Y(n11596) );
  INVX1 U3971 ( .A(n11596), .Y(n2113) );
  AND2X1 U3972 ( .A(ram[455]), .B(n10780), .Y(n11584) );
  INVX1 U3973 ( .A(n11584), .Y(n2114) );
  AND2X1 U3974 ( .A(ram[441]), .B(n10778), .Y(n11567) );
  INVX1 U3975 ( .A(n11567), .Y(n2115) );
  AND2X1 U3976 ( .A(ram[428]), .B(n10778), .Y(n11554) );
  INVX1 U3977 ( .A(n11554), .Y(n2116) );
  AND2X1 U3978 ( .A(ram[415]), .B(n10778), .Y(n11541) );
  INVX1 U3979 ( .A(n11541), .Y(n2117) );
  AND2X1 U3980 ( .A(ram[402]), .B(n10778), .Y(n11528) );
  INVX1 U3981 ( .A(n11528), .Y(n2118) );
  AND2X1 U3982 ( .A(ram[390]), .B(n10778), .Y(n11516) );
  INVX1 U3983 ( .A(n11516), .Y(n2119) );
  AND2X1 U3984 ( .A(ram[376]), .B(n10776), .Y(n11500) );
  INVX1 U3985 ( .A(n11500), .Y(n2120) );
  AND2X1 U3986 ( .A(ram[363]), .B(n10776), .Y(n11487) );
  INVX1 U3987 ( .A(n11487), .Y(n2121) );
  AND2X1 U3988 ( .A(ram[350]), .B(n10776), .Y(n11474) );
  INVX1 U3989 ( .A(n11474), .Y(n2122) );
  AND2X1 U3990 ( .A(ram[337]), .B(n10776), .Y(n11461) );
  INVX1 U3991 ( .A(n11461), .Y(n2123) );
  AND2X1 U3992 ( .A(ram[325]), .B(n10776), .Y(n11449) );
  INVX1 U3993 ( .A(n11449), .Y(n2124) );
  AND2X1 U3994 ( .A(ram[311]), .B(n10774), .Y(n11433) );
  INVX1 U3995 ( .A(n11433), .Y(n2125) );
  AND2X1 U3996 ( .A(ram[298]), .B(n10774), .Y(n11420) );
  INVX1 U3997 ( .A(n11420), .Y(n2126) );
  AND2X1 U3998 ( .A(ram[285]), .B(n10774), .Y(n11407) );
  INVX1 U3999 ( .A(n11407), .Y(n2127) );
  AND2X1 U4000 ( .A(ram[272]), .B(n10774), .Y(n11394) );
  INVX1 U4001 ( .A(n11394), .Y(n2128) );
  AND2X1 U4002 ( .A(ram[260]), .B(n10774), .Y(n11382) );
  INVX1 U4003 ( .A(n11382), .Y(n2129) );
  AND2X1 U4004 ( .A(ram[246]), .B(n10772), .Y(n11366) );
  INVX1 U4005 ( .A(n11366), .Y(n2130) );
  AND2X1 U4006 ( .A(ram[233]), .B(n10772), .Y(n11353) );
  INVX1 U4007 ( .A(n11353), .Y(n2131) );
  AND2X1 U4008 ( .A(ram[220]), .B(n10772), .Y(n11340) );
  INVX1 U4009 ( .A(n11340), .Y(n2132) );
  AND2X1 U4010 ( .A(ram[207]), .B(n10772), .Y(n11327) );
  INVX1 U4011 ( .A(n11327), .Y(n2133) );
  AND2X1 U4012 ( .A(ram[195]), .B(n10772), .Y(n11315) );
  INVX1 U4013 ( .A(n11315), .Y(n2134) );
  AND2X1 U4014 ( .A(ram[181]), .B(n10770), .Y(n11299) );
  INVX1 U4015 ( .A(n11299), .Y(n2135) );
  AND2X1 U4016 ( .A(ram[168]), .B(n10770), .Y(n11286) );
  INVX1 U4017 ( .A(n11286), .Y(n2136) );
  AND2X1 U4018 ( .A(ram[155]), .B(n10770), .Y(n11273) );
  INVX1 U4019 ( .A(n11273), .Y(n2137) );
  AND2X1 U4020 ( .A(ram[142]), .B(n10770), .Y(n11260) );
  INVX1 U4022 ( .A(n11260), .Y(n2138) );
  AND2X1 U4023 ( .A(ram[130]), .B(n10770), .Y(n11248) );
  INVX1 U4024 ( .A(n11248), .Y(n2139) );
  AND2X1 U4025 ( .A(ram[116]), .B(n10768), .Y(n11232) );
  INVX1 U4026 ( .A(n11232), .Y(n2140) );
  AND2X1 U4027 ( .A(ram[103]), .B(n10768), .Y(n11219) );
  INVX1 U4028 ( .A(n11219), .Y(n2141) );
  AND2X1 U4029 ( .A(ram[90]), .B(n10768), .Y(n11206) );
  INVX1 U4030 ( .A(n11206), .Y(n2142) );
  AND2X1 U4031 ( .A(ram[77]), .B(n10768), .Y(n11193) );
  INVX1 U4032 ( .A(n11193), .Y(n2143) );
  AND2X1 U4033 ( .A(ram[65]), .B(n10768), .Y(n11181) );
  INVX1 U4034 ( .A(n11181), .Y(n2144) );
  AND2X1 U4035 ( .A(ram[51]), .B(n10766), .Y(n11165) );
  INVX1 U4036 ( .A(n11165), .Y(n2145) );
  AND2X1 U4037 ( .A(ram[38]), .B(n10766), .Y(n11152) );
  INVX1 U4038 ( .A(n11152), .Y(n2146) );
  AND2X1 U4039 ( .A(ram[25]), .B(n10766), .Y(n11139) );
  INVX1 U4040 ( .A(n11139), .Y(n2147) );
  AND2X1 U4041 ( .A(ram[12]), .B(n10766), .Y(n11126) );
  INVX1 U4042 ( .A(n11126), .Y(n2148) );
  AND2X1 U4043 ( .A(ram[0]), .B(n10766), .Y(n11114) );
  INVX1 U4044 ( .A(n11114), .Y(n2149) );
  BUFX2 U4045 ( .A(n11045), .Y(n2150) );
  BUFX2 U4046 ( .A(n10967), .Y(n2151) );
  BUFX2 U4047 ( .A(n11017), .Y(n2152) );
  BUFX2 U4048 ( .A(n11575), .Y(n2153) );
  INVX1 U4049 ( .A(n4245), .Y(n4257) );
  INVX1 U4050 ( .A(n4245), .Y(n4258) );
  INVX1 U4051 ( .A(n4245), .Y(n4259) );
  INVX1 U4052 ( .A(n4244), .Y(n4260) );
  INVX1 U4053 ( .A(n4244), .Y(n4261) );
  INVX1 U4054 ( .A(n4244), .Y(n4262) );
  INVX1 U4055 ( .A(n4243), .Y(n4263) );
  INVX1 U4056 ( .A(n4243), .Y(n4264) );
  INVX1 U4057 ( .A(n4243), .Y(n4265) );
  INVX1 U4058 ( .A(n4242), .Y(n4266) );
  INVX1 U4059 ( .A(n4242), .Y(n4267) );
  INVX1 U4060 ( .A(n4242), .Y(n4268) );
  INVX1 U4061 ( .A(n4241), .Y(n4269) );
  INVX1 U4062 ( .A(n4241), .Y(n4270) );
  INVX1 U4063 ( .A(n4241), .Y(n4271) );
  INVX1 U4064 ( .A(n4240), .Y(n4272) );
  INVX1 U4065 ( .A(n4240), .Y(n4273) );
  INVX1 U4066 ( .A(n4240), .Y(n4274) );
  INVX1 U4067 ( .A(n4239), .Y(n4275) );
  INVX1 U4068 ( .A(n4239), .Y(n4276) );
  INVX1 U4069 ( .A(n4239), .Y(n4277) );
  INVX1 U4070 ( .A(n4238), .Y(n4278) );
  INVX1 U4071 ( .A(n4238), .Y(n4279) );
  INVX1 U4072 ( .A(n4238), .Y(n4280) );
  INVX1 U4073 ( .A(n4237), .Y(n4281) );
  INVX1 U4074 ( .A(n4237), .Y(n4282) );
  INVX1 U4075 ( .A(n4237), .Y(n4283) );
  INVX1 U4076 ( .A(n4236), .Y(n4284) );
  INVX1 U4077 ( .A(n4236), .Y(n4285) );
  INVX1 U4078 ( .A(n4236), .Y(n4286) );
  INVX1 U4079 ( .A(n4235), .Y(n4287) );
  INVX1 U4080 ( .A(n4235), .Y(n4288) );
  INVX1 U4081 ( .A(n4235), .Y(n4289) );
  INVX1 U4082 ( .A(n4234), .Y(n4290) );
  INVX1 U4083 ( .A(n4234), .Y(n4291) );
  INVX1 U4084 ( .A(n4234), .Y(n4292) );
  INVX1 U4085 ( .A(n4233), .Y(n4293) );
  INVX1 U4086 ( .A(n4233), .Y(n4294) );
  INVX1 U4087 ( .A(n4233), .Y(n4295) );
  INVX1 U4088 ( .A(n4232), .Y(n4296) );
  INVX1 U4089 ( .A(n4232), .Y(n4297) );
  INVX1 U4090 ( .A(n4232), .Y(n4298) );
  INVX1 U4091 ( .A(n4231), .Y(n4299) );
  INVX1 U4092 ( .A(n4231), .Y(n4300) );
  INVX1 U4093 ( .A(n4231), .Y(n4301) );
  INVX1 U4094 ( .A(n4230), .Y(n4302) );
  INVX1 U4095 ( .A(n4230), .Y(n4303) );
  INVX1 U4096 ( .A(n4230), .Y(n4304) );
  INVX1 U4097 ( .A(n4234), .Y(n4305) );
  INVX1 U4098 ( .A(n4236), .Y(n4306) );
  INVX1 U4099 ( .A(n4229), .Y(n4307) );
  INVX1 U4100 ( .A(n4226), .Y(n4308) );
  INVX1 U4101 ( .A(n10636), .Y(n10719) );
  INVX1 U4102 ( .A(n10636), .Y(n10718) );
  INVX1 U4103 ( .A(n10636), .Y(n10717) );
  INVX1 U4104 ( .A(n10637), .Y(n10716) );
  INVX1 U4105 ( .A(n10637), .Y(n10715) );
  INVX1 U4106 ( .A(n10637), .Y(n10714) );
  INVX1 U4107 ( .A(n10638), .Y(n10713) );
  INVX1 U4108 ( .A(n10638), .Y(n10712) );
  INVX1 U4109 ( .A(n10638), .Y(n10711) );
  INVX1 U4110 ( .A(n10639), .Y(n10710) );
  INVX1 U4111 ( .A(n10639), .Y(n10709) );
  INVX1 U4112 ( .A(n10639), .Y(n10708) );
  INVX1 U4113 ( .A(n10640), .Y(n10707) );
  INVX1 U4114 ( .A(n10640), .Y(n10706) );
  INVX1 U4115 ( .A(n10640), .Y(n10705) );
  INVX1 U4116 ( .A(n10641), .Y(n10704) );
  INVX1 U4117 ( .A(n10641), .Y(n10703) );
  INVX1 U4118 ( .A(n10641), .Y(n10702) );
  INVX1 U4119 ( .A(n10642), .Y(n10701) );
  INVX1 U4120 ( .A(n10642), .Y(n10700) );
  INVX1 U4121 ( .A(n10642), .Y(n10699) );
  INVX1 U4122 ( .A(n10643), .Y(n10698) );
  INVX1 U4123 ( .A(n10643), .Y(n10697) );
  INVX1 U4124 ( .A(n10643), .Y(n10696) );
  INVX1 U4125 ( .A(n10644), .Y(n10695) );
  INVX1 U4126 ( .A(n10644), .Y(n10694) );
  INVX1 U4127 ( .A(n10644), .Y(n10693) );
  INVX1 U4128 ( .A(n10645), .Y(n10692) );
  INVX1 U4129 ( .A(n10645), .Y(n10691) );
  INVX1 U4130 ( .A(n10645), .Y(n10690) );
  INVX1 U4131 ( .A(n10646), .Y(n10689) );
  INVX1 U4132 ( .A(n10646), .Y(n10688) );
  INVX1 U4133 ( .A(n10646), .Y(n10687) );
  INVX1 U4134 ( .A(n10647), .Y(n10686) );
  INVX1 U4135 ( .A(n10647), .Y(n10685) );
  INVX1 U4136 ( .A(n10647), .Y(n10684) );
  INVX1 U4137 ( .A(n10648), .Y(n10683) );
  INVX1 U4138 ( .A(n10648), .Y(n10682) );
  INVX1 U4139 ( .A(n10648), .Y(n10681) );
  INVX1 U4140 ( .A(n10649), .Y(n10680) );
  INVX1 U4141 ( .A(n10649), .Y(n10679) );
  INVX1 U4142 ( .A(n10649), .Y(n10678) );
  INVX1 U4143 ( .A(n10650), .Y(n10677) );
  INVX1 U4144 ( .A(n10650), .Y(n10676) );
  INVX1 U4145 ( .A(n10650), .Y(n10675) );
  INVX1 U4146 ( .A(n10651), .Y(n10674) );
  INVX1 U4147 ( .A(n10651), .Y(n10673) );
  INVX1 U4148 ( .A(n10651), .Y(n10672) );
  INVX1 U4149 ( .A(n10652), .Y(n10671) );
  INVX1 U4150 ( .A(n10652), .Y(n10670) );
  INVX1 U4151 ( .A(n10652), .Y(n10669) );
  INVX1 U4152 ( .A(n10653), .Y(n10668) );
  INVX1 U4154 ( .A(n10653), .Y(n10667) );
  INVX1 U4155 ( .A(n10653), .Y(n10666) );
  INVX1 U4156 ( .A(n8478), .Y(n8491) );
  INVX1 U4157 ( .A(n8478), .Y(n8492) );
  INVX1 U4158 ( .A(n8478), .Y(n8493) );
  INVX1 U4159 ( .A(n8477), .Y(n8494) );
  INVX1 U4160 ( .A(n8477), .Y(n8495) );
  INVX1 U4161 ( .A(n8477), .Y(n8496) );
  INVX1 U4162 ( .A(n8476), .Y(n8497) );
  INVX1 U4163 ( .A(n8476), .Y(n8498) );
  INVX1 U4164 ( .A(n8476), .Y(n8499) );
  INVX1 U4165 ( .A(n8475), .Y(n8500) );
  INVX1 U4166 ( .A(n8475), .Y(n8501) );
  INVX1 U4167 ( .A(n8475), .Y(n8502) );
  INVX1 U4168 ( .A(n8474), .Y(n8503) );
  INVX1 U4169 ( .A(n8474), .Y(n8504) );
  INVX1 U4170 ( .A(n8474), .Y(n8505) );
  INVX1 U4171 ( .A(n8473), .Y(n8506) );
  INVX1 U4172 ( .A(n8473), .Y(n8507) );
  INVX1 U4173 ( .A(n8473), .Y(n8508) );
  INVX1 U4174 ( .A(n8472), .Y(n8509) );
  INVX1 U4175 ( .A(n8472), .Y(n8510) );
  INVX1 U4176 ( .A(n8472), .Y(n8511) );
  INVX1 U4177 ( .A(n8471), .Y(n8512) );
  INVX1 U4178 ( .A(n8471), .Y(n8513) );
  INVX1 U4179 ( .A(n8471), .Y(n8514) );
  INVX1 U4180 ( .A(n8470), .Y(n8515) );
  INVX1 U4181 ( .A(n8470), .Y(n8516) );
  INVX1 U4182 ( .A(n8470), .Y(n8517) );
  INVX1 U4183 ( .A(n8469), .Y(n8518) );
  INVX1 U4184 ( .A(n8469), .Y(n8519) );
  INVX1 U4185 ( .A(n8469), .Y(n8520) );
  INVX1 U4186 ( .A(n8468), .Y(n8521) );
  INVX1 U4187 ( .A(n8468), .Y(n8522) );
  INVX1 U4188 ( .A(n8468), .Y(n8523) );
  INVX1 U4189 ( .A(n8467), .Y(n8524) );
  INVX1 U4190 ( .A(n8467), .Y(n8525) );
  INVX1 U4191 ( .A(n8467), .Y(n8526) );
  INVX1 U4192 ( .A(n8466), .Y(n8527) );
  INVX1 U4193 ( .A(n8466), .Y(n8528) );
  INVX1 U4194 ( .A(n8466), .Y(n8529) );
  INVX1 U4195 ( .A(n8465), .Y(n8530) );
  INVX1 U4196 ( .A(n8465), .Y(n8531) );
  INVX1 U4197 ( .A(n8465), .Y(n8532) );
  INVX1 U4198 ( .A(n8464), .Y(n8533) );
  INVX1 U4199 ( .A(n8464), .Y(n8534) );
  INVX1 U4200 ( .A(n8464), .Y(n8535) );
  INVX1 U4201 ( .A(n8463), .Y(n8536) );
  INVX1 U4202 ( .A(n8463), .Y(n8537) );
  INVX1 U4203 ( .A(n8464), .Y(n8538) );
  INVX1 U4204 ( .A(n8463), .Y(n8539) );
  INVX1 U4205 ( .A(n8463), .Y(n8540) );
  INVX1 U4206 ( .A(n8463), .Y(n8541) );
  INVX1 U4207 ( .A(n8475), .Y(n8542) );
  INVX1 U4208 ( .A(n8465), .Y(n8543) );
  INVX1 U4209 ( .A(n8465), .Y(n8544) );
  INVX1 U4210 ( .A(n4229), .Y(n4309) );
  INVX1 U4211 ( .A(n4229), .Y(n4310) );
  INVX1 U4212 ( .A(n4229), .Y(n4311) );
  INVX1 U4213 ( .A(n4228), .Y(n4312) );
  INVX1 U4214 ( .A(n4228), .Y(n4313) );
  INVX1 U4215 ( .A(n4228), .Y(n4314) );
  INVX1 U4216 ( .A(n4227), .Y(n4315) );
  INVX1 U4217 ( .A(n4227), .Y(n4316) );
  INVX1 U4218 ( .A(n4226), .Y(n4317) );
  INVX1 U4219 ( .A(n4226), .Y(n4318) );
  INVX1 U4220 ( .A(n4226), .Y(n4319) );
  INVX1 U4221 ( .A(n4225), .Y(n4320) );
  INVX1 U4222 ( .A(n4225), .Y(n4321) );
  INVX1 U4223 ( .A(n4225), .Y(n4322) );
  INVX1 U4224 ( .A(n4227), .Y(n4323) );
  INVX1 U4225 ( .A(n4225), .Y(n4324) );
  INVX1 U4226 ( .A(n10639), .Y(n10737) );
  INVX1 U4227 ( .A(n10641), .Y(n10736) );
  INVX1 U4228 ( .A(n10655), .Y(n10735) );
  INVX1 U4229 ( .A(n10640), .Y(n10734) );
  INVX1 U4230 ( .A(n10640), .Y(n10733) );
  INVX1 U4231 ( .A(n10641), .Y(n10732) );
  INVX1 U4232 ( .A(n10634), .Y(n10731) );
  INVX1 U4233 ( .A(n10634), .Y(n10730) );
  INVX1 U4234 ( .A(n10634), .Y(n10729) );
  INVX1 U4235 ( .A(n10643), .Y(n10728) );
  INVX1 U4236 ( .A(n10637), .Y(n10727) );
  INVX1 U4237 ( .A(n10654), .Y(n10726) );
  INVX1 U4238 ( .A(n10653), .Y(n10725) );
  INVX1 U4239 ( .A(n10642), .Y(n10724) );
  INVX1 U4240 ( .A(n10638), .Y(n10723) );
  INVX1 U4241 ( .A(n10635), .Y(n10722) );
  INVX1 U4242 ( .A(n10635), .Y(n10721) );
  INVX1 U4243 ( .A(n10635), .Y(n10720) );
  INVX1 U4244 ( .A(n4247), .Y(n4249) );
  INVX1 U4245 ( .A(n4247), .Y(n4250) );
  INVX1 U4246 ( .A(n4246), .Y(n4251) );
  INVX1 U4247 ( .A(n4246), .Y(n4252) );
  INVX1 U4248 ( .A(n4246), .Y(n4253) );
  INVX1 U4249 ( .A(n4246), .Y(n4254) );
  INVX1 U4250 ( .A(n4330), .Y(n4255) );
  INVX1 U4251 ( .A(n4331), .Y(n4256) );
  INVX1 U4252 ( .A(n10656), .Y(n10659) );
  INVX1 U4253 ( .A(n10656), .Y(n10658) );
  INVX1 U4254 ( .A(n10654), .Y(n10665) );
  INVX1 U4255 ( .A(n10654), .Y(n10664) );
  INVX1 U4256 ( .A(n10654), .Y(n10663) );
  INVX1 U4257 ( .A(n10655), .Y(n10662) );
  INVX1 U4258 ( .A(n10655), .Y(n10661) );
  INVX1 U4259 ( .A(n10655), .Y(n10660) );
  INVX1 U4260 ( .A(n4224), .Y(n4325) );
  INVX1 U4261 ( .A(n4224), .Y(n4326) );
  INVX1 U4262 ( .A(n4224), .Y(n4327) );
  INVX1 U4263 ( .A(n10633), .Y(n10740) );
  INVX1 U4264 ( .A(n10633), .Y(n10739) );
  INVX1 U4265 ( .A(n10633), .Y(n10738) );
  INVX1 U4266 ( .A(n4226), .Y(n4328) );
  INVX1 U4267 ( .A(n4226), .Y(n4329) );
  INVX1 U4268 ( .A(n10633), .Y(n10742) );
  INVX1 U4269 ( .A(n10633), .Y(n10741) );
  INVX1 U4270 ( .A(n11178), .Y(n10767) );
  INVX1 U4271 ( .A(n11113), .Y(n10766) );
  INVX1 U4272 ( .A(n4338), .Y(n4245) );
  INVX1 U4273 ( .A(n4338), .Y(n4244) );
  INVX1 U4274 ( .A(n4338), .Y(n4243) );
  INVX1 U4275 ( .A(n4337), .Y(n4242) );
  INVX1 U4276 ( .A(n4337), .Y(n4241) );
  INVX1 U4277 ( .A(n4337), .Y(n4240) );
  INVX1 U4278 ( .A(n4336), .Y(n4239) );
  INVX1 U4279 ( .A(n4336), .Y(n4238) );
  INVX1 U4280 ( .A(n4336), .Y(n4237) );
  INVX1 U4281 ( .A(n4335), .Y(n4236) );
  INVX1 U4282 ( .A(n4335), .Y(n4235) );
  INVX1 U4286 ( .A(n4335), .Y(n4234) );
  INVX1 U4289 ( .A(n4334), .Y(n4233) );
  INVX1 U4290 ( .A(n4334), .Y(n4232) );
  INVX1 U4291 ( .A(n4334), .Y(n4231) );
  INVX1 U4292 ( .A(n4332), .Y(n4230) );
  INVX1 U4293 ( .A(n10744), .Y(n10636) );
  INVX1 U4294 ( .A(n10744), .Y(n10637) );
  INVX1 U4295 ( .A(n10744), .Y(n10638) );
  INVX1 U4296 ( .A(n10747), .Y(n10639) );
  INVX1 U4297 ( .A(n10744), .Y(n10640) );
  INVX1 U4298 ( .A(n10748), .Y(n10641) );
  INVX1 U4299 ( .A(n10744), .Y(n10642) );
  INVX1 U4300 ( .A(n10746), .Y(n10643) );
  INVX1 U4301 ( .A(n10747), .Y(n10644) );
  INVX1 U4302 ( .A(n10745), .Y(n10645) );
  INVX1 U4303 ( .A(n10745), .Y(n10646) );
  INVX1 U4304 ( .A(n10745), .Y(n10647) );
  INVX1 U4305 ( .A(n10746), .Y(n10648) );
  INVX1 U4306 ( .A(n10746), .Y(n10649) );
  INVX1 U4307 ( .A(n10746), .Y(n10650) );
  INVX1 U4308 ( .A(n10747), .Y(n10651) );
  INVX1 U4309 ( .A(n10747), .Y(n10652) );
  INVX1 U4310 ( .A(n10747), .Y(n10653) );
  INVX1 U4311 ( .A(n4247), .Y(n4248) );
  INVX1 U4312 ( .A(n10656), .Y(n10657) );
  INVX1 U4313 ( .A(n8461), .Y(n8545) );
  INVX1 U4314 ( .A(n8462), .Y(n8546) );
  INVX1 U4315 ( .A(n8463), .Y(n8547) );
  INVX1 U4316 ( .A(n8472), .Y(n8548) );
  INVX1 U4317 ( .A(n8476), .Y(n8549) );
  INVX1 U4318 ( .A(n8464), .Y(n8550) );
  INVX1 U4319 ( .A(n8462), .Y(n8551) );
  INVX1 U4320 ( .A(n8462), .Y(n8552) );
  INVX1 U4321 ( .A(n8462), .Y(n8553) );
  INVX1 U4322 ( .A(n8461), .Y(n8554) );
  INVX1 U4323 ( .A(n8461), .Y(n8555) );
  INVX1 U4324 ( .A(n8461), .Y(n8556) );
  INVX1 U4325 ( .A(n8462), .Y(n8557) );
  INVX1 U4326 ( .A(n8476), .Y(n8558) );
  INVX1 U4327 ( .A(n8461), .Y(n8559) );
  INVX1 U4328 ( .A(n8461), .Y(n8560) );
  INVX1 U4329 ( .A(n8461), .Y(n8561) );
  INVX1 U4330 ( .A(n8462), .Y(n8562) );
  INVX1 U4331 ( .A(n8481), .Y(n8483) );
  INVX1 U4332 ( .A(n8481), .Y(n8484) );
  INVX1 U4333 ( .A(n8480), .Y(n8485) );
  INVX1 U4334 ( .A(n8480), .Y(n8486) );
  INVX1 U4335 ( .A(n8480), .Y(n8487) );
  INVX1 U4336 ( .A(n8479), .Y(n8488) );
  INVX1 U4337 ( .A(n8479), .Y(n8489) );
  INVX1 U4338 ( .A(n8479), .Y(n8490) );
  INVX1 U4339 ( .A(n8464), .Y(n8563) );
  INVX1 U4340 ( .A(n8462), .Y(n8564) );
  INVX1 U4341 ( .A(n8465), .Y(n8565) );
  INVX1 U4342 ( .A(n8461), .Y(n8566) );
  INVX1 U4343 ( .A(n8461), .Y(n8567) );
  INVX1 U4344 ( .A(n8574), .Y(n8478) );
  INVX1 U4345 ( .A(n8574), .Y(n8477) );
  INVX1 U4346 ( .A(n8574), .Y(n8476) );
  INVX1 U4347 ( .A(n8573), .Y(n8475) );
  INVX1 U4348 ( .A(n8573), .Y(n8474) );
  INVX1 U4349 ( .A(n8573), .Y(n8473) );
  INVX1 U4350 ( .A(n8572), .Y(n8472) );
  INVX1 U4351 ( .A(n8572), .Y(n8471) );
  INVX1 U4352 ( .A(n8572), .Y(n8470) );
  INVX1 U4353 ( .A(n8571), .Y(n8469) );
  INVX1 U4354 ( .A(n8571), .Y(n8468) );
  INVX1 U4355 ( .A(n8571), .Y(n8467) );
  INVX1 U4356 ( .A(n8570), .Y(n8466) );
  INVX1 U4357 ( .A(n8570), .Y(n8465) );
  INVX1 U4358 ( .A(n8570), .Y(n8464) );
  INVX1 U4359 ( .A(n8570), .Y(n8463) );
  INVX1 U4360 ( .A(n8481), .Y(n8482) );
  INVX1 U4361 ( .A(n4178), .Y(n4201) );
  INVX1 U4362 ( .A(n4178), .Y(n4202) );
  INVX1 U4363 ( .A(n4178), .Y(n4203) );
  INVX1 U4364 ( .A(n4177), .Y(n4204) );
  INVX1 U4365 ( .A(n4181), .Y(n4205) );
  INVX1 U4366 ( .A(n4178), .Y(n4206) );
  INVX1 U4367 ( .A(n4177), .Y(n4207) );
  INVX1 U4368 ( .A(n4177), .Y(n4208) );
  INVX1 U4369 ( .A(n4177), .Y(n4209) );
  INVX1 U4370 ( .A(n4176), .Y(n4210) );
  INVX1 U4371 ( .A(n4176), .Y(n4211) );
  INVX1 U4372 ( .A(n4176), .Y(n4212) );
  INVX1 U4373 ( .A(n4176), .Y(n4213) );
  INVX1 U4374 ( .A(n4176), .Y(n4214) );
  INVX1 U4375 ( .A(n4178), .Y(n4215) );
  INVX1 U4376 ( .A(n4181), .Y(n4216) );
  INVX1 U4377 ( .A(n4177), .Y(n4217) );
  INVX1 U4378 ( .A(n4178), .Y(n4218) );
  INVX1 U4379 ( .A(n4177), .Y(n4219) );
  INVX1 U4380 ( .A(n4179), .Y(n4220) );
  INVX1 U4381 ( .A(n4181), .Y(n4221) );
  INVX1 U4382 ( .A(n4181), .Y(n4222) );
  INVX1 U4383 ( .A(n10962), .Y(n4158) );
  INVX1 U4384 ( .A(n10962), .Y(n4159) );
  INVX1 U4385 ( .A(n10962), .Y(n4160) );
  INVX1 U4386 ( .A(n10962), .Y(n4161) );
  INVX1 U4387 ( .A(n10962), .Y(n4162) );
  INVX1 U4388 ( .A(n10962), .Y(n4163) );
  INVX1 U4389 ( .A(n10962), .Y(n4164) );
  INVX1 U4390 ( .A(n10962), .Y(n4165) );
  INVX1 U4391 ( .A(n10962), .Y(n4166) );
  INVX1 U4392 ( .A(n10962), .Y(n4167) );
  INVX1 U4393 ( .A(n10962), .Y(n4168) );
  INVX1 U4394 ( .A(n10962), .Y(n4169) );
  INVX1 U4395 ( .A(n10962), .Y(n4170) );
  INVX1 U4396 ( .A(n10962), .Y(n4171) );
  INVX1 U4397 ( .A(n10962), .Y(n4172) );
  INVX1 U4398 ( .A(n10962), .Y(n4173) );
  INVX1 U4399 ( .A(n11043), .Y(n10762) );
  INVX1 U4400 ( .A(n11043), .Y(n10761) );
  INVX1 U4401 ( .A(n4182), .Y(n4184) );
  INVX1 U4402 ( .A(n4182), .Y(n4185) );
  INVX1 U4403 ( .A(n4182), .Y(n4186) );
  INVX1 U4404 ( .A(n4180), .Y(n4187) );
  INVX1 U4405 ( .A(n4179), .Y(n4188) );
  INVX1 U4406 ( .A(n4181), .Y(n4189) );
  INVX1 U4407 ( .A(n4181), .Y(n4190) );
  INVX1 U4408 ( .A(n4181), .Y(n4191) );
  INVX1 U4409 ( .A(n4179), .Y(n4192) );
  INVX1 U4410 ( .A(n4181), .Y(n4193) );
  INVX1 U4411 ( .A(n4181), .Y(n4194) );
  INVX1 U4412 ( .A(n4180), .Y(n4195) );
  INVX1 U4413 ( .A(n4180), .Y(n4196) );
  INVX1 U4414 ( .A(n4180), .Y(n4197) );
  INVX1 U4415 ( .A(n4179), .Y(n4198) );
  INVX1 U4416 ( .A(n4179), .Y(n4199) );
  INVX1 U4417 ( .A(n4179), .Y(n4200) );
  INVX1 U4418 ( .A(n10584), .Y(n10631) );
  INVX1 U4419 ( .A(n10584), .Y(n10630) );
  INVX1 U4420 ( .A(n10584), .Y(n10629) );
  INVX1 U4421 ( .A(n10584), .Y(n10628) );
  INVX1 U4422 ( .A(n10584), .Y(n10627) );
  INVX1 U4423 ( .A(n10584), .Y(n10626) );
  INVX1 U4424 ( .A(n10587), .Y(n10625) );
  INVX1 U4425 ( .A(n10588), .Y(n10624) );
  INVX1 U4426 ( .A(n10589), .Y(n10623) );
  INVX1 U4427 ( .A(n10587), .Y(n10622) );
  INVX1 U4428 ( .A(n10588), .Y(n10621) );
  INVX1 U4429 ( .A(n10585), .Y(n10620) );
  INVX1 U4430 ( .A(n10586), .Y(n10619) );
  INVX1 U4431 ( .A(n10585), .Y(n10618) );
  INVX1 U4432 ( .A(n10588), .Y(n10617) );
  INVX1 U4433 ( .A(n10589), .Y(n10616) );
  INVX1 U4434 ( .A(n10586), .Y(n10615) );
  INVX1 U4435 ( .A(n10586), .Y(n10614) );
  INVX1 U4436 ( .A(n10589), .Y(n10613) );
  INVX1 U4437 ( .A(n10587), .Y(n10612) );
  INVX1 U4438 ( .A(n10588), .Y(n10611) );
  INVX1 U4439 ( .A(n10585), .Y(n10610) );
  INVX1 U4440 ( .A(n10587), .Y(n10609) );
  INVX1 U4441 ( .A(n10586), .Y(n10608) );
  INVX1 U4442 ( .A(n10584), .Y(n10607) );
  INVX1 U4443 ( .A(n10589), .Y(n10606) );
  INVX1 U4444 ( .A(n10585), .Y(n10605) );
  INVX1 U4445 ( .A(n10585), .Y(n10604) );
  INVX1 U4446 ( .A(n10585), .Y(n10603) );
  INVX1 U4447 ( .A(n10585), .Y(n10602) );
  INVX1 U4448 ( .A(n10586), .Y(n10601) );
  INVX1 U4449 ( .A(n10586), .Y(n10600) );
  INVX1 U4450 ( .A(n10586), .Y(n10599) );
  INVX1 U4451 ( .A(n10587), .Y(n10598) );
  INVX1 U4452 ( .A(n10587), .Y(n10597) );
  INVX1 U4453 ( .A(n10587), .Y(n10596) );
  INVX1 U4454 ( .A(n10588), .Y(n10595) );
  INVX1 U4455 ( .A(n10588), .Y(n10594) );
  INVX1 U4456 ( .A(n10588), .Y(n10593) );
  INVX1 U4457 ( .A(n10589), .Y(n10592) );
  INVX1 U4458 ( .A(n10589), .Y(n10591) );
  INVX1 U4459 ( .A(n10964), .Y(n4153) );
  INVX1 U4460 ( .A(n10964), .Y(n4154) );
  INVX1 U4461 ( .A(n10964), .Y(n4155) );
  INVX1 U4462 ( .A(n10567), .Y(n10583) );
  INVX1 U4463 ( .A(n10567), .Y(n10582) );
  INVX1 U4464 ( .A(n10567), .Y(n10581) );
  INVX1 U4465 ( .A(n10567), .Y(n10580) );
  INVX1 U4466 ( .A(n10567), .Y(n10579) );
  INVX1 U4467 ( .A(n10567), .Y(n10578) );
  INVX1 U4468 ( .A(n10567), .Y(n10577) );
  INVX1 U4469 ( .A(n10567), .Y(n10576) );
  INVX1 U4470 ( .A(n10567), .Y(n10575) );
  INVX1 U4471 ( .A(n10567), .Y(n10574) );
  INVX1 U4472 ( .A(n10567), .Y(n10573) );
  INVX1 U4473 ( .A(n10567), .Y(n10572) );
  INVX1 U4474 ( .A(n10567), .Y(n10571) );
  INVX1 U4475 ( .A(n10567), .Y(n10570) );
  INVX1 U4476 ( .A(n10567), .Y(n10569) );
  INVX1 U4477 ( .A(n10567), .Y(n10568) );
  INVX1 U4478 ( .A(n10566), .Y(n10565) );
  INVX1 U4479 ( .A(n10566), .Y(n10564) );
  INVX1 U4480 ( .A(n10566), .Y(n10563) );
  INVX1 U4481 ( .A(n10962), .Y(n4174) );
  INVX1 U4482 ( .A(n10962), .Y(n4175) );
  INVX1 U4483 ( .A(n11244), .Y(n10769) );
  INVX1 U4484 ( .A(n11310), .Y(n10771) );
  INVX1 U4485 ( .A(n11376), .Y(n10773) );
  INVX1 U4486 ( .A(n11442), .Y(n10775) );
  INVX1 U4490 ( .A(n11508), .Y(n10777) );
  INVX1 U4495 ( .A(n11574), .Y(n10779) );
  INVX1 U4496 ( .A(n11641), .Y(n10781) );
  INVX1 U4497 ( .A(n11707), .Y(n10783) );
  INVX1 U4498 ( .A(n11773), .Y(n10785) );
  INVX1 U4499 ( .A(n11839), .Y(n10787) );
  INVX1 U4500 ( .A(n11905), .Y(n10789) );
  INVX1 U4501 ( .A(n11971), .Y(n10791) );
  INVX1 U4502 ( .A(n12037), .Y(n10793) );
  INVX1 U4503 ( .A(n12103), .Y(n10795) );
  INVX1 U4504 ( .A(n12170), .Y(n10797) );
  INVX1 U4505 ( .A(n12236), .Y(n10799) );
  INVX1 U4506 ( .A(n12302), .Y(n10801) );
  INVX1 U4507 ( .A(n12368), .Y(n10803) );
  INVX1 U4508 ( .A(n12434), .Y(n10805) );
  INVX1 U4509 ( .A(n12500), .Y(n10807) );
  INVX1 U4510 ( .A(n12566), .Y(n10809) );
  INVX1 U4511 ( .A(n12632), .Y(n10811) );
  INVX1 U4512 ( .A(n12699), .Y(n10813) );
  INVX1 U4513 ( .A(n12765), .Y(n10815) );
  INVX1 U4514 ( .A(n12831), .Y(n10817) );
  INVX1 U4515 ( .A(n12897), .Y(n10819) );
  INVX1 U4516 ( .A(n12963), .Y(n10821) );
  INVX1 U4517 ( .A(n13029), .Y(n10823) );
  INVX1 U4518 ( .A(n13095), .Y(n10825) );
  INVX1 U4519 ( .A(n13225), .Y(n10953) );
  INVX1 U4520 ( .A(n4182), .Y(n4183) );
  INVX1 U4521 ( .A(n11642), .Y(n10782) );
  INVX1 U4522 ( .A(n12171), .Y(n10798) );
  INVX1 U4523 ( .A(n12700), .Y(n10814) );
  INVX1 U4524 ( .A(n11179), .Y(n10768) );
  INVX1 U4525 ( .A(n11245), .Y(n10770) );
  INVX1 U4526 ( .A(n11311), .Y(n10772) );
  INVX1 U4527 ( .A(n11377), .Y(n10774) );
  INVX1 U4528 ( .A(n11443), .Y(n10776) );
  INVX1 U4529 ( .A(n11509), .Y(n10778) );
  INVX1 U4530 ( .A(n11708), .Y(n10784) );
  INVX1 U4531 ( .A(n11774), .Y(n10786) );
  INVX1 U4532 ( .A(n11840), .Y(n10788) );
  INVX1 U4533 ( .A(n11906), .Y(n10790) );
  INVX1 U4534 ( .A(n11972), .Y(n10792) );
  INVX1 U4535 ( .A(n12038), .Y(n10794) );
  INVX1 U4536 ( .A(n12237), .Y(n10800) );
  INVX1 U4537 ( .A(n12303), .Y(n10802) );
  INVX1 U4538 ( .A(n12369), .Y(n10804) );
  INVX1 U4539 ( .A(n12435), .Y(n10806) );
  INVX1 U4540 ( .A(n12501), .Y(n10808) );
  INVX1 U4541 ( .A(n12567), .Y(n10810) );
  INVX1 U4542 ( .A(n12766), .Y(n10816) );
  INVX1 U4543 ( .A(n12832), .Y(n10818) );
  INVX1 U4544 ( .A(n12898), .Y(n10820) );
  INVX1 U4545 ( .A(n12964), .Y(n10822) );
  INVX1 U4546 ( .A(n13030), .Y(n10824) );
  INVX1 U4547 ( .A(n13097), .Y(n10952) );
  INVX1 U4548 ( .A(n11576), .Y(n10780) );
  INVX1 U4549 ( .A(n12105), .Y(n10796) );
  INVX1 U4550 ( .A(n12634), .Y(n10812) );
  INVX1 U4551 ( .A(n10589), .Y(n10590) );
  INVX1 U4552 ( .A(n4330), .Y(n4338) );
  INVX1 U4553 ( .A(n4330), .Y(n4337) );
  INVX1 U4554 ( .A(n4330), .Y(n4336) );
  INVX1 U4555 ( .A(n4331), .Y(n4335) );
  INVX1 U4556 ( .A(n4331), .Y(n4334) );
  INVX1 U4557 ( .A(n10743), .Y(n10744) );
  INVX1 U4558 ( .A(n10633), .Y(n10745) );
  INVX1 U4559 ( .A(n10743), .Y(n10746) );
  INVX1 U4560 ( .A(n10743), .Y(n10747) );
  INVX1 U4561 ( .A(n4333), .Y(n4229) );
  INVX1 U4562 ( .A(n4333), .Y(n4228) );
  INVX1 U4563 ( .A(n4333), .Y(n4227) );
  INVX1 U4564 ( .A(n4332), .Y(n4226) );
  INVX1 U4565 ( .A(n4332), .Y(n4225) );
  INVX1 U4566 ( .A(n10748), .Y(n10634) );
  INVX1 U4567 ( .A(n10745), .Y(n10635) );
  INVX1 U4568 ( .A(n10957), .Y(n4247) );
  INVX1 U4569 ( .A(n10957), .Y(n4246) );
  INVX1 U4570 ( .A(n10748), .Y(n10656) );
  INVX1 U4571 ( .A(n10748), .Y(n10654) );
  INVX1 U4572 ( .A(n10748), .Y(n10655) );
  INVX1 U4573 ( .A(n4332), .Y(n4224) );
  INVX1 U4574 ( .A(read2_addr[4]), .Y(n10633) );
  INVX1 U4575 ( .A(n8395), .Y(n8396) );
  INVX1 U4576 ( .A(n8395), .Y(n8397) );
  INVX1 U4577 ( .A(n8395), .Y(n8398) );
  INVX1 U4578 ( .A(n8395), .Y(n8399) );
  INVX1 U4579 ( .A(n8395), .Y(n8400) );
  INVX1 U4580 ( .A(n8395), .Y(n8401) );
  INVX1 U4581 ( .A(n8395), .Y(n8402) );
  INVX1 U4582 ( .A(n8395), .Y(n8403) );
  INVX1 U4583 ( .A(n8395), .Y(n8404) );
  INVX1 U4584 ( .A(n8395), .Y(n8405) );
  INVX1 U4585 ( .A(n8395), .Y(n8406) );
  INVX1 U4586 ( .A(n8395), .Y(n8407) );
  INVX1 U4587 ( .A(n8395), .Y(n8409) );
  INVX1 U4588 ( .A(n8395), .Y(n8410) );
  INVX1 U4589 ( .A(n11110), .Y(n10765) );
  INVX1 U4590 ( .A(n8414), .Y(n8434) );
  INVX1 U4591 ( .A(n8414), .Y(n8435) );
  INVX1 U4592 ( .A(n8414), .Y(n8436) );
  INVX1 U4593 ( .A(n8413), .Y(n8437) );
  INVX1 U4594 ( .A(n8414), .Y(n8438) );
  INVX1 U4595 ( .A(n8413), .Y(n8439) );
  INVX1 U4596 ( .A(n8413), .Y(n8440) );
  INVX1 U4597 ( .A(n8413), .Y(n8441) );
  INVX1 U4598 ( .A(n8413), .Y(n8442) );
  INVX1 U4599 ( .A(n8412), .Y(n8443) );
  INVX1 U4600 ( .A(n8412), .Y(n8444) );
  INVX1 U4601 ( .A(n8412), .Y(n8445) );
  INVX1 U4602 ( .A(n8411), .Y(n8446) );
  INVX1 U4603 ( .A(n8411), .Y(n8447) );
  INVX1 U4604 ( .A(n8411), .Y(n8448) );
  INVX1 U4605 ( .A(n8412), .Y(n8449) );
  INVX1 U4606 ( .A(n8411), .Y(n8450) );
  INVX1 U4607 ( .A(n8411), .Y(n8451) );
  INVX1 U4608 ( .A(n8412), .Y(n8452) );
  INVX1 U4609 ( .A(n8411), .Y(n8453) );
  INVX1 U4610 ( .A(n8411), .Y(n8454) );
  INVX1 U4611 ( .A(n8412), .Y(n8455) );
  INVX1 U4612 ( .A(n8413), .Y(n8456) );
  INVX1 U4613 ( .A(n8411), .Y(n8457) );
  INVX1 U4614 ( .A(n8459), .Y(n8417) );
  INVX1 U4615 ( .A(n8412), .Y(n8418) );
  INVX1 U4616 ( .A(n8459), .Y(n8419) );
  INVX1 U4617 ( .A(n8415), .Y(n8420) );
  INVX1 U4618 ( .A(n8412), .Y(n8421) );
  INVX1 U4619 ( .A(n8415), .Y(n8422) );
  INVX1 U4620 ( .A(n8415), .Y(n8423) );
  INVX1 U4621 ( .A(n8415), .Y(n8424) );
  INVX1 U4622 ( .A(n8413), .Y(n8425) );
  INVX1 U4623 ( .A(n8411), .Y(n8426) );
  INVX1 U4624 ( .A(n8414), .Y(n8427) );
  INVX1 U4625 ( .A(n8415), .Y(n8428) );
  INVX1 U4626 ( .A(n8413), .Y(n8429) );
  INVX1 U4627 ( .A(n8412), .Y(n8430) );
  INVX1 U4628 ( .A(n8412), .Y(n8431) );
  INVX1 U4629 ( .A(n8414), .Y(n8432) );
  INVX1 U4630 ( .A(n8415), .Y(n8433) );
  INVX1 U4631 ( .A(n8414), .Y(n8416) );
  INVX1 U4632 ( .A(n8569), .Y(n8574) );
  INVX1 U4633 ( .A(n8569), .Y(n8573) );
  INVX1 U4634 ( .A(n8569), .Y(n8572) );
  INVX1 U4635 ( .A(n8569), .Y(n8571) );
  INVX1 U4636 ( .A(n8569), .Y(n8570) );
  INVX1 U4637 ( .A(n8571), .Y(n8462) );
  INVX1 U4638 ( .A(n8571), .Y(n8461) );
  INVX1 U4639 ( .A(n8575), .Y(n8481) );
  INVX1 U4640 ( .A(n8575), .Y(n8480) );
  INVX1 U4641 ( .A(n8575), .Y(n8479) );
  INVX1 U4642 ( .A(n8388), .Y(n8389) );
  INVX1 U4643 ( .A(n8388), .Y(n8390) );
  INVX1 U4644 ( .A(n8388), .Y(n8391) );
  INVX1 U4645 ( .A(n8388), .Y(n8392) );
  INVX1 U4646 ( .A(n8388), .Y(n8393) );
  INVX1 U4647 ( .A(n8395), .Y(n8408) );
  INVX1 U4648 ( .A(n10584), .Y(n10632) );
  INVX1 U4649 ( .A(n10964), .Y(n4156) );
  INVX1 U4650 ( .A(n10964), .Y(n4157) );
  INVX1 U4651 ( .A(n4223), .Y(n4178) );
  INVX1 U4652 ( .A(n4223), .Y(n4177) );
  INVX1 U4653 ( .A(n4223), .Y(n4176) );
  INVX1 U4654 ( .A(n4223), .Y(n4182) );
  INVX1 U4655 ( .A(n4223), .Y(n4181) );
  INVX1 U4656 ( .A(n4223), .Y(n4180) );
  INVX1 U4657 ( .A(n4223), .Y(n4179) );
  INVX1 U4658 ( .A(read2_addr[3]), .Y(n10584) );
  INVX1 U4659 ( .A(n10957), .Y(n4330) );
  INVX1 U4660 ( .A(n10957), .Y(n4331) );
  INVX1 U4661 ( .A(read2_addr[2]), .Y(n10567) );
  INVX1 U4662 ( .A(n10626), .Y(n10585) );
  INVX1 U4663 ( .A(n10632), .Y(n10586) );
  INVX1 U4664 ( .A(n10630), .Y(n10587) );
  INVX1 U4665 ( .A(n10631), .Y(n10588) );
  INVX1 U4666 ( .A(n10628), .Y(n10589) );
  INVX1 U4667 ( .A(n4331), .Y(n4333) );
  INVX1 U4668 ( .A(n4331), .Y(n4332) );
  INVX1 U4669 ( .A(n10743), .Y(n10748) );
  INVX1 U4670 ( .A(n8413), .Y(n8458) );
  INVX1 U4671 ( .A(read1_addr[2]), .Y(n8395) );
  INVX1 U4672 ( .A(n8460), .Y(n8414) );
  INVX1 U4673 ( .A(n8460), .Y(n8413) );
  INVX1 U4674 ( .A(n8460), .Y(n8412) );
  INVX1 U4675 ( .A(n8460), .Y(n8411) );
  INVX1 U4676 ( .A(n8460), .Y(n8415) );
  INVX1 U4677 ( .A(read1_addr[4]), .Y(n8569) );
  INVX1 U4678 ( .A(n8568), .Y(n8575) );
  INVX1 U4679 ( .A(read1_addr[4]), .Y(n8568) );
  INVX1 U4680 ( .A(n10965), .Y(n4152) );
  INVX1 U4681 ( .A(n10965), .Y(n4151) );
  INVX1 U4682 ( .A(n10965), .Y(n4150) );
  INVX1 U4683 ( .A(n10560), .Y(n10561) );
  INVX1 U4684 ( .A(n10560), .Y(n10562) );
  INVX1 U4685 ( .A(n8388), .Y(n8394) );
  INVX1 U4686 ( .A(read1_addr[1]), .Y(n8388) );
  INVX1 U4687 ( .A(n10960), .Y(n4223) );
  INVX1 U4688 ( .A(n11047), .Y(Dout1[63]) );
  INVX1 U4689 ( .A(n8320), .Y(n119) );
  INVX1 U4690 ( .A(n11048), .Y(Dout1[62]) );
  INVX1 U4691 ( .A(n8321), .Y(n118) );
  INVX1 U4692 ( .A(n11049), .Y(Dout1[61]) );
  INVX1 U4693 ( .A(n8322), .Y(n117) );
  INVX1 U4694 ( .A(n11050), .Y(Dout1[60]) );
  INVX1 U4695 ( .A(n8323), .Y(n116) );
  INVX1 U4696 ( .A(n11051), .Y(Dout1[59]) );
  INVX1 U4697 ( .A(n8324), .Y(n115) );
  INVX1 U4698 ( .A(n11052), .Y(Dout1[58]) );
  INVX1 U4699 ( .A(n8325), .Y(n114) );
  INVX1 U4700 ( .A(n11094), .Y(Dout1[16]) );
  INVX1 U4701 ( .A(n8367), .Y(n72) );
  INVX1 U4702 ( .A(n11095), .Y(Dout1[15]) );
  INVX1 U4703 ( .A(n8368), .Y(n71) );
  INVX1 U4704 ( .A(n11096), .Y(Dout1[14]) );
  INVX1 U4705 ( .A(n8369), .Y(n70) );
  INVX1 U4706 ( .A(n11097), .Y(Dout1[13]) );
  INVX1 U4707 ( .A(n8370), .Y(n69) );
  INVX1 U4708 ( .A(n11098), .Y(Dout1[12]) );
  INVX1 U4709 ( .A(n8371), .Y(n68) );
  INVX1 U4710 ( .A(n11099), .Y(Dout1[11]) );
  INVX1 U4711 ( .A(n8372), .Y(n67) );
  INVX1 U4712 ( .A(n11100), .Y(Dout1[10]) );
  INVX1 U4713 ( .A(n8373), .Y(n66) );
  INVX1 U4714 ( .A(n11101), .Y(Dout1[9]) );
  INVX1 U4715 ( .A(n8374), .Y(n65) );
  INVX1 U4716 ( .A(n11102), .Y(Dout1[8]) );
  INVX1 U4717 ( .A(n8375), .Y(n64) );
  INVX1 U4718 ( .A(n11103), .Y(Dout1[7]) );
  INVX1 U4719 ( .A(n8376), .Y(n63) );
  INVX1 U4720 ( .A(n11104), .Y(Dout1[6]) );
  INVX1 U4721 ( .A(n8377), .Y(n62) );
  INVX1 U4722 ( .A(n11105), .Y(Dout1[5]) );
  INVX1 U4723 ( .A(n8378), .Y(n61) );
  INVX1 U4724 ( .A(n11106), .Y(Dout1[4]) );
  INVX1 U4725 ( .A(n8379), .Y(n60) );
  INVX1 U4726 ( .A(n11107), .Y(Dout1[3]) );
  INVX1 U4727 ( .A(n8380), .Y(n59) );
  INVX1 U4728 ( .A(n11108), .Y(Dout1[2]) );
  INVX1 U4729 ( .A(n8381), .Y(n58) );
  INVX1 U4730 ( .A(n11054), .Y(Dout1[56]) );
  INVX1 U4731 ( .A(n8327), .Y(n112) );
  INVX1 U4732 ( .A(n11090), .Y(Dout1[20]) );
  INVX1 U4733 ( .A(n8363), .Y(n76) );
  INVX1 U4734 ( .A(n11111), .Y(Dout1[0]) );
  INVX1 U4735 ( .A(n8383), .Y(n56) );
  INVX1 U4736 ( .A(n11053), .Y(Dout1[57]) );
  INVX1 U4737 ( .A(n8326), .Y(n113) );
  INVX1 U4738 ( .A(n11089), .Y(Dout1[21]) );
  INVX1 U4739 ( .A(n8362), .Y(n77) );
  INVX1 U4740 ( .A(n11093), .Y(Dout1[17]) );
  INVX1 U4741 ( .A(n8366), .Y(n73) );
  INVX1 U4742 ( .A(n11109), .Y(Dout1[1]) );
  INVX1 U4743 ( .A(n8382), .Y(n57) );
  INVX1 U4744 ( .A(n11056), .Y(Dout1[54]) );
  INVX1 U4745 ( .A(n8329), .Y(n110) );
  INVX1 U4746 ( .A(n11060), .Y(Dout1[50]) );
  INVX1 U4747 ( .A(n8333), .Y(n106) );
  INVX1 U4748 ( .A(n11064), .Y(Dout1[46]) );
  INVX1 U4749 ( .A(n8337), .Y(n102) );
  INVX1 U4750 ( .A(n11072), .Y(Dout1[38]) );
  INVX1 U4751 ( .A(n8345), .Y(n94) );
  INVX1 U4752 ( .A(n11080), .Y(Dout1[30]) );
  INVX1 U4753 ( .A(n8353), .Y(n86) );
  INVX1 U4754 ( .A(n11055), .Y(Dout1[55]) );
  INVX1 U4755 ( .A(n8328), .Y(n111) );
  INVX1 U4756 ( .A(n11059), .Y(Dout1[51]) );
  INVX1 U4757 ( .A(n8332), .Y(n107) );
  INVX1 U4758 ( .A(n11063), .Y(Dout1[47]) );
  INVX1 U4759 ( .A(n8336), .Y(n103) );
  INVX1 U4760 ( .A(n11071), .Y(Dout1[39]) );
  INVX1 U4761 ( .A(n8344), .Y(n95) );
  INVX1 U4762 ( .A(n11079), .Y(Dout1[31]) );
  INVX1 U4763 ( .A(n8352), .Y(n87) );
  INVX1 U4764 ( .A(n11057), .Y(Dout1[53]) );
  INVX1 U4765 ( .A(n8330), .Y(n109) );
  INVX1 U4766 ( .A(n11058), .Y(Dout1[52]) );
  INVX1 U4767 ( .A(n8331), .Y(n108) );
  INVX1 U4768 ( .A(n11061), .Y(Dout1[49]) );
  INVX1 U4769 ( .A(n8334), .Y(n105) );
  INVX1 U4770 ( .A(n11062), .Y(Dout1[48]) );
  INVX1 U4771 ( .A(n8335), .Y(n104) );
  INVX1 U4772 ( .A(n11065), .Y(Dout1[45]) );
  INVX1 U4773 ( .A(n8338), .Y(n101) );
  INVX1 U4774 ( .A(n11066), .Y(Dout1[44]) );
  INVX1 U4775 ( .A(n8339), .Y(n100) );
  INVX1 U4776 ( .A(n11067), .Y(Dout1[43]) );
  INVX1 U4777 ( .A(n8340), .Y(n99) );
  INVX1 U4778 ( .A(n11068), .Y(Dout1[42]) );
  INVX1 U4779 ( .A(n8341), .Y(n98) );
  INVX1 U4780 ( .A(n11069), .Y(Dout1[41]) );
  INVX1 U4781 ( .A(n8342), .Y(n97) );
  INVX1 U4782 ( .A(n11070), .Y(Dout1[40]) );
  INVX1 U4783 ( .A(n8343), .Y(n96) );
  INVX1 U4784 ( .A(n11073), .Y(Dout1[37]) );
  INVX1 U4785 ( .A(n8346), .Y(n93) );
  INVX1 U4786 ( .A(n11074), .Y(Dout1[36]) );
  INVX1 U4787 ( .A(n8347), .Y(n92) );
  INVX1 U4788 ( .A(n11075), .Y(Dout1[35]) );
  INVX1 U4789 ( .A(n8348), .Y(n91) );
  INVX1 U4790 ( .A(n11076), .Y(Dout1[34]) );
  INVX1 U4791 ( .A(n8349), .Y(n90) );
  INVX1 U4792 ( .A(n11077), .Y(Dout1[33]) );
  INVX1 U4793 ( .A(n8350), .Y(n89) );
  INVX1 U4794 ( .A(n11078), .Y(Dout1[32]) );
  INVX1 U4795 ( .A(n8351), .Y(n88) );
  INVX1 U4796 ( .A(n11081), .Y(Dout1[29]) );
  INVX1 U4797 ( .A(n8354), .Y(n85) );
  INVX1 U4798 ( .A(n11082), .Y(Dout1[28]) );
  INVX1 U4799 ( .A(n8355), .Y(n84) );
  INVX1 U4800 ( .A(n11083), .Y(Dout1[27]) );
  INVX1 U4801 ( .A(n8356), .Y(n83) );
  INVX1 U4802 ( .A(n11084), .Y(Dout1[26]) );
  INVX1 U4803 ( .A(n8357), .Y(n82) );
  INVX1 U4804 ( .A(n11085), .Y(Dout1[25]) );
  INVX1 U4805 ( .A(n8358), .Y(n81) );
  INVX1 U4806 ( .A(n11086), .Y(Dout1[24]) );
  INVX1 U4807 ( .A(n8359), .Y(n80) );
  INVX1 U4808 ( .A(n11087), .Y(Dout1[23]) );
  INVX1 U4809 ( .A(n8360), .Y(n79) );
  INVX1 U4810 ( .A(n11088), .Y(Dout1[22]) );
  INVX1 U4811 ( .A(n8361), .Y(n78) );
  INVX1 U4812 ( .A(n11091), .Y(Dout1[19]) );
  INVX1 U4813 ( .A(n8364), .Y(n75) );
  INVX1 U4814 ( .A(n11092), .Y(Dout1[18]) );
  INVX1 U4815 ( .A(n8365), .Y(n74) );
  INVX1 U4816 ( .A(n8459), .Y(n8460) );
  BUFX2 U4817 ( .A(n1835), .Y(n10749) );
  BUFX2 U4818 ( .A(n1519), .Y(n10752) );
  BUFX2 U4819 ( .A(n1835), .Y(n10750) );
  BUFX2 U4820 ( .A(n1519), .Y(n10753) );
  BUFX2 U4821 ( .A(n1676), .Y(n10755) );
  BUFX2 U4822 ( .A(n1393), .Y(n10758) );
  BUFX2 U4823 ( .A(n1676), .Y(n10756) );
  BUFX2 U4824 ( .A(n1393), .Y(n10759) );
  INVX1 U4825 ( .A(n10877), .Y(n10876) );
  INVX1 U4826 ( .A(n13149), .Y(n10877) );
  INVX1 U4827 ( .A(n4111), .Y(current_ram[38]) );
  INVX1 U4828 ( .A(n8384), .Y(n8387) );
  INVX1 U4829 ( .A(n8384), .Y(n8386) );
  INVX1 U4830 ( .A(n8384), .Y(n8385) );
  INVX1 U4831 ( .A(n2155), .Y(n10754) );
  INVX1 U4832 ( .A(n2156), .Y(n10760) );
  INVX1 U4833 ( .A(n2154), .Y(n10751) );
  INVX1 U4834 ( .A(n2157), .Y(n10757) );
  INVX1 U4835 ( .A(read2_addr[0]), .Y(n10560) );
  INVX1 U4836 ( .A(n10875), .Y(n10874) );
  INVX1 U4837 ( .A(n13147), .Y(n10875) );
  INVX1 U4838 ( .A(n4110), .Y(current_ram[39]) );
  INVX1 U4839 ( .A(n10841), .Y(n10840) );
  INVX1 U4840 ( .A(n13113), .Y(n10841) );
  INVX1 U4841 ( .A(n4093), .Y(current_ram[56]) );
  INVX1 U4842 ( .A(n10843), .Y(n10842) );
  INVX1 U4843 ( .A(n13115), .Y(n10843) );
  INVX1 U4844 ( .A(n4094), .Y(current_ram[55]) );
  INVX1 U4845 ( .A(n10847), .Y(n10846) );
  INVX1 U4846 ( .A(n13119), .Y(n10847) );
  INVX1 U4847 ( .A(n4096), .Y(current_ram[53]) );
  INVX1 U4848 ( .A(n10849), .Y(n10848) );
  INVX1 U4849 ( .A(n13121), .Y(n10849) );
  INVX1 U4850 ( .A(n4097), .Y(current_ram[52]) );
  INVX1 U4851 ( .A(n10853), .Y(n10852) );
  INVX1 U4852 ( .A(n13125), .Y(n10853) );
  INVX1 U4853 ( .A(n4099), .Y(current_ram[50]) );
  INVX1 U4854 ( .A(n10855), .Y(n10854) );
  INVX1 U4855 ( .A(n13127), .Y(n10855) );
  INVX1 U4856 ( .A(n4100), .Y(current_ram[49]) );
  INVX1 U4857 ( .A(n10861), .Y(n10860) );
  INVX1 U4858 ( .A(n13133), .Y(n10861) );
  INVX1 U4859 ( .A(n4103), .Y(current_ram[46]) );
  INVX1 U4860 ( .A(n10863), .Y(n10862) );
  INVX1 U4861 ( .A(n13135), .Y(n10863) );
  INVX1 U4862 ( .A(n4104), .Y(current_ram[45]) );
  INVX1 U4863 ( .A(n10867), .Y(n10866) );
  INVX1 U4864 ( .A(n13139), .Y(n10867) );
  INVX1 U4865 ( .A(n4106), .Y(current_ram[43]) );
  INVX1 U4866 ( .A(n10869), .Y(n10868) );
  INVX1 U4867 ( .A(n13141), .Y(n10869) );
  INVX1 U4868 ( .A(n4107), .Y(current_ram[42]) );
  INVX1 U4869 ( .A(n10871), .Y(n10870) );
  INVX1 U4870 ( .A(n13143), .Y(n10871) );
  INVX1 U4871 ( .A(n4108), .Y(current_ram[41]) );
  INVX1 U4872 ( .A(n10873), .Y(n10872) );
  INVX1 U4873 ( .A(n13145), .Y(n10873) );
  INVX1 U4874 ( .A(n4109), .Y(current_ram[40]) );
  INVX1 U4875 ( .A(n10905), .Y(n10904) );
  INVX1 U4876 ( .A(n13177), .Y(n10905) );
  INVX1 U4877 ( .A(n4125), .Y(current_ram[24]) );
  INVX1 U4878 ( .A(n10913), .Y(n10912) );
  INVX1 U4879 ( .A(n13185), .Y(n10913) );
  INVX1 U4880 ( .A(n4129), .Y(current_ram[20]) );
  INVX1 U4881 ( .A(n10917), .Y(n10916) );
  INVX1 U4882 ( .A(n13189), .Y(n10917) );
  INVX1 U4883 ( .A(n4131), .Y(current_ram[18]) );
  INVX1 U4884 ( .A(n10921), .Y(n10920) );
  INVX1 U4885 ( .A(n13193), .Y(n10921) );
  INVX1 U4886 ( .A(n4133), .Y(current_ram[16]) );
  INVX1 U4887 ( .A(n10923), .Y(n10922) );
  INVX1 U4888 ( .A(n13195), .Y(n10923) );
  INVX1 U4889 ( .A(n4134), .Y(current_ram[15]) );
  INVX1 U4890 ( .A(n10925), .Y(n10924) );
  INVX1 U4891 ( .A(n13197), .Y(n10925) );
  INVX1 U4892 ( .A(n4135), .Y(current_ram[14]) );
  INVX1 U4893 ( .A(n10927), .Y(n10926) );
  INVX1 U4894 ( .A(n13199), .Y(n10927) );
  INVX1 U4895 ( .A(n4136), .Y(current_ram[13]) );
  INVX1 U4896 ( .A(n10929), .Y(n10928) );
  INVX1 U4897 ( .A(n13201), .Y(n10929) );
  INVX1 U4898 ( .A(n4137), .Y(current_ram[12]) );
  INVX1 U4899 ( .A(n10931), .Y(n10930) );
  INVX1 U4900 ( .A(n13203), .Y(n10931) );
  INVX1 U4901 ( .A(n4138), .Y(current_ram[11]) );
  INVX1 U4902 ( .A(n10933), .Y(n10932) );
  INVX1 U4903 ( .A(n13205), .Y(n10933) );
  INVX1 U4904 ( .A(n4139), .Y(current_ram[10]) );
  INVX1 U4905 ( .A(n10935), .Y(n10934) );
  INVX1 U4906 ( .A(n13207), .Y(n10935) );
  INVX1 U4907 ( .A(n4140), .Y(current_ram[9]) );
  INVX1 U4908 ( .A(n10937), .Y(n10936) );
  INVX1 U4909 ( .A(n13209), .Y(n10937) );
  INVX1 U4910 ( .A(n4141), .Y(current_ram[8]) );
  INVX1 U4911 ( .A(n10955), .Y(n10954) );
  INVX1 U4912 ( .A(n13226), .Y(n10955) );
  INVX1 U4913 ( .A(n4149), .Y(current_ram[0]) );
  INVX1 U4914 ( .A(n10939), .Y(n10938) );
  INVX1 U4915 ( .A(n13211), .Y(n10939) );
  INVX1 U4916 ( .A(n4142), .Y(current_ram[7]) );
  INVX1 U4917 ( .A(n10851), .Y(n10850) );
  INVX1 U4918 ( .A(n13123), .Y(n10851) );
  INVX1 U4919 ( .A(n4098), .Y(current_ram[51]) );
  INVX1 U4920 ( .A(n10883), .Y(n10882) );
  INVX1 U4921 ( .A(n13155), .Y(n10883) );
  INVX1 U4922 ( .A(n4114), .Y(current_ram[35]) );
  INVX1 U4923 ( .A(n10907), .Y(n10906) );
  INVX1 U4924 ( .A(n13179), .Y(n10907) );
  INVX1 U4925 ( .A(n4126), .Y(current_ram[23]) );
  INVX1 U4926 ( .A(n10911), .Y(n10910) );
  INVX1 U4927 ( .A(n13183), .Y(n10911) );
  INVX1 U4928 ( .A(n4128), .Y(current_ram[21]) );
  INVX1 U4929 ( .A(n10943), .Y(n10942) );
  INVX1 U4930 ( .A(read2_addr[4]), .Y(n10743) );
  INVX1 U4931 ( .A(read2_addr[1]), .Y(n10566) );
  INVX1 U4932 ( .A(reset), .Y(n10956) );
  INVX1 U4933 ( .A(read1_addr[3]), .Y(n8459) );
  INVX1 U4934 ( .A(n10829), .Y(n10828) );
  INVX1 U4935 ( .A(n13101), .Y(n10829) );
  INVX1 U4936 ( .A(n10833), .Y(n10832) );
  INVX1 U4937 ( .A(n13105), .Y(n10833) );
  INVX1 U4938 ( .A(n10837), .Y(n10836) );
  INVX1 U4939 ( .A(n13109), .Y(n10837) );
  INVX1 U4940 ( .A(n10879), .Y(n10878) );
  INVX1 U4941 ( .A(n13151), .Y(n10879) );
  INVX1 U4942 ( .A(n4112), .Y(current_ram[37]) );
  INVX1 U4943 ( .A(n10881), .Y(n10880) );
  INVX1 U4944 ( .A(n13153), .Y(n10881) );
  INVX1 U4945 ( .A(n4113), .Y(current_ram[36]) );
  INVX1 U4946 ( .A(n10885), .Y(n10884) );
  INVX1 U4947 ( .A(n13157), .Y(n10885) );
  INVX1 U4948 ( .A(n4115), .Y(current_ram[34]) );
  INVX1 U4949 ( .A(n10887), .Y(n10886) );
  INVX1 U4950 ( .A(n13159), .Y(n10887) );
  INVX1 U4951 ( .A(n4116), .Y(current_ram[33]) );
  INVX1 U4952 ( .A(n10889), .Y(n10888) );
  INVX1 U4953 ( .A(n13161), .Y(n10889) );
  INVX1 U4954 ( .A(n4117), .Y(current_ram[32]) );
  INVX1 U4955 ( .A(n10919), .Y(n10918) );
  INVX1 U4956 ( .A(n13191), .Y(n10919) );
  INVX1 U4957 ( .A(n4132), .Y(current_ram[17]) );
  INVX1 U4958 ( .A(n10497), .Y(n185) );
  INVX1 U4959 ( .A(n10496), .Y(n186) );
  INVX1 U4960 ( .A(n10534), .Y(n148) );
  INVX1 U4961 ( .A(n10533), .Y(n149) );
  INVX1 U4962 ( .A(n10531), .Y(n151) );
  INVX1 U4963 ( .A(n10530), .Y(n152) );
  INVX1 U4964 ( .A(n10529), .Y(n153) );
  INVX1 U4965 ( .A(n10528), .Y(n154) );
  INVX1 U4966 ( .A(n10501), .Y(n181) );
  INVX1 U4967 ( .A(n10500), .Y(n182) );
  INVX1 U4968 ( .A(n10499), .Y(n183) );
  INVX1 U4969 ( .A(n10498), .Y(n184) );
  INVX1 U4970 ( .A(n11044), .Y(Dout2[0]) );
  INVX1 U4971 ( .A(n11041), .Y(Dout2[1]) );
  INVX1 U4972 ( .A(n11040), .Y(Dout2[2]) );
  INVX1 U4973 ( .A(n11039), .Y(Dout2[3]) );
  INVX1 U4974 ( .A(n11038), .Y(Dout2[4]) );
  INVX1 U4975 ( .A(n11037), .Y(Dout2[5]) );
  INVX1 U4976 ( .A(n11036), .Y(Dout2[6]) );
  INVX1 U4977 ( .A(n11035), .Y(Dout2[7]) );
  INVX1 U4978 ( .A(n11034), .Y(Dout2[8]) );
  INVX1 U4979 ( .A(n11032), .Y(Dout2[9]) );
  INVX1 U4980 ( .A(n11031), .Y(Dout2[10]) );
  INVX1 U4981 ( .A(n11030), .Y(Dout2[11]) );
  INVX1 U4982 ( .A(n11029), .Y(Dout2[12]) );
  INVX1 U4983 ( .A(n11028), .Y(Dout2[13]) );
  INVX1 U4984 ( .A(n11027), .Y(Dout2[14]) );
  INVX1 U4985 ( .A(n11026), .Y(Dout2[15]) );
  INVX1 U4986 ( .A(n11025), .Y(Dout2[16]) );
  INVX1 U4987 ( .A(n11024), .Y(Dout2[17]) );
  INVX1 U4988 ( .A(n11023), .Y(Dout2[18]) );
  INVX1 U4989 ( .A(n11022), .Y(Dout2[19]) );
  INVX1 U4990 ( .A(n11021), .Y(Dout2[20]) );
  INVX1 U4991 ( .A(n11020), .Y(Dout2[21]) );
  INVX1 U4992 ( .A(n11019), .Y(Dout2[22]) );
  INVX1 U4993 ( .A(n11018), .Y(Dout2[23]) );
  INVX1 U4994 ( .A(n11013), .Y(Dout2[24]) );
  INVX1 U4995 ( .A(n11010), .Y(Dout2[27]) );
  INVX1 U4996 ( .A(n11004), .Y(Dout2[32]) );
  INVX1 U4997 ( .A(n11002), .Y(Dout2[33]) );
  INVX1 U4998 ( .A(n11001), .Y(Dout2[34]) );
  INVX1 U4999 ( .A(n11000), .Y(Dout2[35]) );
  INVX1 U5000 ( .A(n10999), .Y(Dout2[36]) );
  INVX1 U5001 ( .A(n10998), .Y(Dout2[37]) );
  INVX1 U5002 ( .A(n10997), .Y(Dout2[38]) );
  INVX1 U5003 ( .A(n10996), .Y(Dout2[39]) );
  INVX1 U5004 ( .A(n10995), .Y(Dout2[40]) );
  INVX1 U5005 ( .A(n10993), .Y(Dout2[41]) );
  INVX1 U5006 ( .A(n10992), .Y(Dout2[42]) );
  INVX1 U5007 ( .A(n10991), .Y(Dout2[43]) );
  INVX1 U5008 ( .A(n10990), .Y(Dout2[44]) );
  INVX1 U5009 ( .A(n10989), .Y(Dout2[45]) );
  INVX1 U5010 ( .A(n10988), .Y(Dout2[46]) );
  INVX1 U5011 ( .A(n10987), .Y(Dout2[47]) );
  INVX1 U5012 ( .A(n10986), .Y(Dout2[48]) );
  INVX1 U5013 ( .A(n10985), .Y(Dout2[49]) );
  INVX1 U5014 ( .A(n10984), .Y(Dout2[50]) );
  INVX1 U5015 ( .A(n10983), .Y(Dout2[51]) );
  INVX1 U5016 ( .A(n10982), .Y(Dout2[52]) );
  INVX1 U5017 ( .A(n10981), .Y(Dout2[53]) );
  INVX1 U5018 ( .A(n10980), .Y(Dout2[54]) );
  INVX1 U5019 ( .A(n10979), .Y(Dout2[55]) );
  INVX1 U5020 ( .A(n10976), .Y(Dout2[56]) );
  INVX1 U5021 ( .A(n10975), .Y(Dout2[57]) );
  INVX1 U5022 ( .A(n10960), .Y(n10959) );
  INVX1 U5023 ( .A(n1678), .Y(n13229) );
  INVX1 U5024 ( .A(n10958), .Y(n10957) );
  INVX1 U5025 ( .A(n10962), .Y(n10961) );
  INVX1 U5026 ( .A(n10966), .Y(n11005) );
  INVX1 U5027 ( .A(n4086), .Y(current_ram[63]) );
  INVX1 U5028 ( .A(n4087), .Y(current_ram[62]) );
  INVX1 U5029 ( .A(n4088), .Y(current_ram[61]) );
  INVX1 U5030 ( .A(n4089), .Y(current_ram[60]) );
  INVX1 U5031 ( .A(n4090), .Y(current_ram[59]) );
  INVX1 U5032 ( .A(n4091), .Y(current_ram[58]) );
  INVX1 U5033 ( .A(n4118), .Y(current_ram[31]) );
  INVX1 U5034 ( .A(n4119), .Y(current_ram[30]) );
  INVX1 U5035 ( .A(n4120), .Y(current_ram[29]) );
  INVX1 U5036 ( .A(n4121), .Y(current_ram[28]) );
  INVX1 U5037 ( .A(n4122), .Y(current_ram[27]) );
  INVX1 U5038 ( .A(n4123), .Y(current_ram[26]) );
  INVX1 U5039 ( .A(n4124), .Y(current_ram[25]) );
  INVX1 U5040 ( .A(n10559), .Y(n123) );
  INVX1 U5041 ( .A(n10558), .Y(n124) );
  INVX1 U5042 ( .A(n10557), .Y(n125) );
  INVX1 U5043 ( .A(n10556), .Y(n126) );
  INVX1 U5044 ( .A(n10555), .Y(n127) );
  INVX1 U5045 ( .A(n10554), .Y(n128) );
  INVX1 U5046 ( .A(n10553), .Y(n129) );
  INVX1 U5047 ( .A(n10552), .Y(n130) );
  INVX1 U5048 ( .A(n10551), .Y(n131) );
  INVX1 U5049 ( .A(n10550), .Y(n132) );
  INVX1 U5050 ( .A(n10549), .Y(n133) );
  INVX1 U5051 ( .A(n10548), .Y(n134) );
  INVX1 U5052 ( .A(n10547), .Y(n135) );
  INVX1 U5053 ( .A(n10546), .Y(n136) );
  INVX1 U5054 ( .A(n10545), .Y(n137) );
  INVX1 U5055 ( .A(n10544), .Y(n138) );
  INVX1 U5056 ( .A(n10543), .Y(n139) );
  INVX1 U5057 ( .A(n10542), .Y(n140) );
  INVX1 U5058 ( .A(n10541), .Y(n141) );
  INVX1 U5059 ( .A(n10540), .Y(n142) );
  INVX1 U5060 ( .A(n10539), .Y(n143) );
  INVX1 U5061 ( .A(n10538), .Y(n144) );
  INVX1 U5062 ( .A(n10537), .Y(n145) );
  INVX1 U5063 ( .A(n10536), .Y(n146) );
  INVX1 U5064 ( .A(n10535), .Y(n147) );
  INVX1 U5065 ( .A(n10532), .Y(n150) );
  INVX1 U5066 ( .A(n10527), .Y(n155) );
  INVX1 U5067 ( .A(n10526), .Y(n156) );
  INVX1 U5068 ( .A(n10525), .Y(n157) );
  INVX1 U5069 ( .A(n10524), .Y(n158) );
  INVX1 U5070 ( .A(n10523), .Y(n159) );
  INVX1 U5071 ( .A(n10522), .Y(n160) );
  INVX1 U5072 ( .A(n10521), .Y(n161) );
  INVX1 U5073 ( .A(n10520), .Y(n162) );
  INVX1 U5074 ( .A(n10519), .Y(n163) );
  INVX1 U5075 ( .A(n10518), .Y(n164) );
  INVX1 U5076 ( .A(n10517), .Y(n165) );
  INVX1 U5077 ( .A(n10516), .Y(n166) );
  INVX1 U5078 ( .A(n10515), .Y(n167) );
  INVX1 U5079 ( .A(n10514), .Y(n168) );
  INVX1 U5080 ( .A(n10513), .Y(n169) );
  INVX1 U5081 ( .A(n10512), .Y(n170) );
  INVX1 U5082 ( .A(n10511), .Y(n171) );
  INVX1 U5083 ( .A(n10510), .Y(n172) );
  INVX1 U5084 ( .A(n10509), .Y(n173) );
  INVX1 U5085 ( .A(n10508), .Y(n174) );
  INVX1 U5086 ( .A(n10507), .Y(n175) );
  INVX1 U5087 ( .A(n10506), .Y(n176) );
  INVX1 U5088 ( .A(n10505), .Y(n177) );
  INVX1 U5089 ( .A(n10504), .Y(n178) );
  INVX1 U5090 ( .A(n10503), .Y(n179) );
  INVX1 U5091 ( .A(n10502), .Y(n180) );
  INVX1 U5092 ( .A(n10964), .Y(n10963) );
  INVX1 U5093 ( .A(read1_addr[0]), .Y(n8384) );
  INVX1 U5094 ( .A(n10827), .Y(n10826) );
  INVX1 U5095 ( .A(n13099), .Y(n10827) );
  INVX1 U5096 ( .A(n10831), .Y(n10830) );
  INVX1 U5097 ( .A(n13103), .Y(n10831) );
  INVX1 U5098 ( .A(n10835), .Y(n10834) );
  INVX1 U5099 ( .A(n13107), .Y(n10835) );
  INVX1 U5100 ( .A(n10891), .Y(n10890) );
  INVX1 U5101 ( .A(n13163), .Y(n10891) );
  INVX1 U5102 ( .A(n10893), .Y(n10892) );
  INVX1 U5103 ( .A(n13165), .Y(n10893) );
  INVX1 U5104 ( .A(n10895), .Y(n10894) );
  INVX1 U5105 ( .A(n13167), .Y(n10895) );
  INVX1 U5106 ( .A(n10897), .Y(n10896) );
  INVX1 U5107 ( .A(n13169), .Y(n10897) );
  INVX1 U5108 ( .A(n10899), .Y(n10898) );
  INVX1 U5109 ( .A(n13171), .Y(n10899) );
  INVX1 U5110 ( .A(n10901), .Y(n10900) );
  INVX1 U5111 ( .A(n13173), .Y(n10901) );
  INVX1 U5112 ( .A(n10903), .Y(n10902) );
  INVX1 U5113 ( .A(n13175), .Y(n10903) );
  INVX1 U5114 ( .A(n10857), .Y(n10856) );
  INVX1 U5115 ( .A(n13129), .Y(n10857) );
  INVX1 U5116 ( .A(n4101), .Y(current_ram[48]) );
  INVX1 U5117 ( .A(n10859), .Y(n10858) );
  INVX1 U5118 ( .A(n13131), .Y(n10859) );
  INVX1 U5119 ( .A(n4102), .Y(current_ram[47]) );
  INVX1 U5120 ( .A(n10865), .Y(n10864) );
  INVX1 U5121 ( .A(n13137), .Y(n10865) );
  INVX1 U5122 ( .A(n4105), .Y(current_ram[44]) );
  INVX1 U5123 ( .A(n10839), .Y(n10838) );
  INVX1 U5124 ( .A(n13111), .Y(n10839) );
  INVX1 U5125 ( .A(n4092), .Y(current_ram[57]) );
  INVX1 U5126 ( .A(n10845), .Y(n10844) );
  INVX1 U5127 ( .A(n13117), .Y(n10845) );
  INVX1 U5128 ( .A(n4095), .Y(current_ram[54]) );
  INVX1 U5129 ( .A(n10909), .Y(n10908) );
  INVX1 U5130 ( .A(n13181), .Y(n10909) );
  INVX1 U5131 ( .A(n4127), .Y(current_ram[22]) );
  INVX1 U5132 ( .A(n10949), .Y(n10948) );
  INVX1 U5133 ( .A(n13221), .Y(n10949) );
  INVX1 U5134 ( .A(n4147), .Y(current_ram[2]) );
  INVX1 U5135 ( .A(n10951), .Y(n10950) );
  INVX1 U5136 ( .A(n13223), .Y(n10951) );
  INVX1 U5137 ( .A(n4148), .Y(current_ram[1]) );
  INVX1 U5138 ( .A(n10915), .Y(n10914) );
  INVX1 U5139 ( .A(n13187), .Y(n10915) );
  INVX1 U5140 ( .A(n4130), .Y(current_ram[19]) );
  INVX1 U5141 ( .A(n10941), .Y(n10940) );
  INVX1 U5142 ( .A(n13213), .Y(n10941) );
  INVX1 U5143 ( .A(n4143), .Y(current_ram[6]) );
  INVX1 U5144 ( .A(n13215), .Y(n10943) );
  INVX1 U5145 ( .A(n4144), .Y(current_ram[5]) );
  INVX1 U5146 ( .A(n10945), .Y(n10944) );
  INVX1 U5147 ( .A(n13217), .Y(n10945) );
  INVX1 U5148 ( .A(n4145), .Y(current_ram[4]) );
  INVX1 U5149 ( .A(n10947), .Y(n10946) );
  INVX1 U5150 ( .A(n13219), .Y(n10947) );
  INVX1 U5151 ( .A(n4146), .Y(current_ram[3]) );
  INVX1 U5152 ( .A(n10970), .Y(Dout2[62]) );
  INVX1 U5153 ( .A(n10969), .Y(Dout2[63]) );
  INVX1 U5154 ( .A(n11012), .Y(Dout2[25]) );
  INVX1 U5155 ( .A(n11011), .Y(Dout2[26]) );
  INVX1 U5156 ( .A(n11009), .Y(Dout2[28]) );
  INVX1 U5157 ( .A(n11008), .Y(Dout2[29]) );
  INVX1 U5158 ( .A(n11007), .Y(Dout2[30]) );
  INVX1 U5159 ( .A(n11006), .Y(Dout2[31]) );
  INVX1 U5160 ( .A(n10974), .Y(Dout2[58]) );
  INVX1 U5161 ( .A(n10973), .Y(Dout2[59]) );
  INVX1 U5162 ( .A(n10972), .Y(Dout2[60]) );
  INVX1 U5163 ( .A(n10971), .Y(Dout2[61]) );
  INVX1 U5164 ( .A(PPP[0]), .Y(n11016) );
  INVX1 U5165 ( .A(write_addr[4]), .Y(n10958) );
  INVX1 U5166 ( .A(write_addr[2]), .Y(n10962) );
  INVX1 U5167 ( .A(write_addr[3]), .Y(n10960) );
  INVX1 U5168 ( .A(write_addr[1]), .Y(n10964) );
  INVX1 U5169 ( .A(write_addr[0]), .Y(n10965) );
  INVX1 U5170 ( .A(PPP[2]), .Y(n13228) );
  INVX1 U5171 ( .A(PPP[1]), .Y(n13227) );
  INVX1 U5172 ( .A(n10978), .Y(n11015) );
  AND2X1 U5173 ( .A(ram[1991]), .B(n10956), .Y(n6660) );
  AND2X1 U5174 ( .A(ram[1992]), .B(n10956), .Y(n6661) );
  AND2X1 U5175 ( .A(ram[1993]), .B(n10956), .Y(n6662) );
  AND2X1 U5176 ( .A(ram[1994]), .B(n10956), .Y(n6663) );
  AND2X1 U5177 ( .A(ram[1995]), .B(n10956), .Y(n6664) );
  AND2X1 U5178 ( .A(ram[1996]), .B(n10956), .Y(n6665) );
  AND2X1 U5179 ( .A(ram[1997]), .B(n10956), .Y(n6666) );
  AND2X1 U5180 ( .A(ram[1998]), .B(n10956), .Y(n6667) );
  AND2X1 U5181 ( .A(ram[1999]), .B(n10956), .Y(n6668) );
  AND2X1 U5182 ( .A(ram[2000]), .B(n10956), .Y(n6669) );
  AND2X1 U5183 ( .A(ram[2001]), .B(n10956), .Y(n6670) );
  AND2X1 U5184 ( .A(ram[2002]), .B(n10956), .Y(n6671) );
  AND2X1 U5185 ( .A(ram[2003]), .B(n10956), .Y(n6672) );
  AND2X1 U5186 ( .A(ram[2004]), .B(n10956), .Y(n6673) );
  AND2X1 U5187 ( .A(ram[2005]), .B(n10956), .Y(n6674) );
  AND2X1 U5188 ( .A(ram[2006]), .B(n10956), .Y(n6675) );
  AND2X1 U5189 ( .A(ram[2007]), .B(n10956), .Y(n6676) );
  AND2X1 U5190 ( .A(ram[2008]), .B(n10956), .Y(n6677) );
  AND2X1 U5191 ( .A(ram[2009]), .B(n10956), .Y(n6678) );
  AND2X1 U5192 ( .A(ram[2010]), .B(n10956), .Y(n6679) );
  AND2X1 U5193 ( .A(ram[2011]), .B(n10956), .Y(n6680) );
  AND2X1 U5194 ( .A(ram[2012]), .B(n10956), .Y(n6681) );
  AND2X1 U5195 ( .A(ram[2013]), .B(n10956), .Y(n6682) );
  AND2X1 U5196 ( .A(ram[2014]), .B(n10956), .Y(n6683) );
  AND2X1 U5197 ( .A(ram[2015]), .B(n10956), .Y(n6684) );
  AND2X1 U5198 ( .A(ram[2016]), .B(n10956), .Y(n6685) );
  AND2X1 U5199 ( .A(ram[2017]), .B(n10956), .Y(n6686) );
  AND2X1 U5200 ( .A(ram[2018]), .B(n10956), .Y(n6687) );
  AND2X1 U5201 ( .A(ram[2019]), .B(n10956), .Y(n6688) );
  AND2X1 U5202 ( .A(ram[2020]), .B(n10956), .Y(n6689) );
  AND2X1 U5203 ( .A(ram[2021]), .B(n10956), .Y(n6690) );
  AND2X1 U5204 ( .A(ram[2022]), .B(n10956), .Y(n6691) );
  AND2X1 U5205 ( .A(ram[2023]), .B(n10956), .Y(n6692) );
  AND2X1 U5206 ( .A(ram[2024]), .B(n10956), .Y(n6693) );
  AND2X1 U5207 ( .A(ram[2025]), .B(n10956), .Y(n6694) );
  AND2X1 U5208 ( .A(ram[2026]), .B(n10956), .Y(n6695) );
  AND2X1 U5209 ( .A(ram[2027]), .B(n10956), .Y(n6696) );
  AND2X1 U5210 ( .A(ram[2028]), .B(n10956), .Y(n6697) );
  AND2X1 U5211 ( .A(ram[2029]), .B(n10956), .Y(n6698) );
  AND2X1 U5212 ( .A(ram[2030]), .B(n10956), .Y(n6699) );
  AND2X1 U5213 ( .A(ram[2031]), .B(n10956), .Y(n6700) );
  AND2X1 U5214 ( .A(ram[2032]), .B(n10956), .Y(n6701) );
  AND2X1 U5215 ( .A(ram[2033]), .B(n10956), .Y(n6702) );
  AND2X1 U5216 ( .A(ram[2034]), .B(n10956), .Y(n6703) );
  AND2X1 U5217 ( .A(ram[2035]), .B(n10956), .Y(n6704) );
  AND2X1 U5218 ( .A(ram[2036]), .B(n10956), .Y(n6705) );
  AND2X1 U5219 ( .A(ram[2037]), .B(n10956), .Y(n6706) );
  AND2X1 U5220 ( .A(ram[2038]), .B(n10956), .Y(n6707) );
  AND2X1 U5221 ( .A(ram[2039]), .B(n10956), .Y(n6708) );
  AND2X1 U5222 ( .A(ram[2040]), .B(n10956), .Y(n6709) );
  AND2X1 U5223 ( .A(ram[2041]), .B(n10956), .Y(n6710) );
  AND2X1 U5224 ( .A(ram[2042]), .B(n10956), .Y(n6711) );
  AND2X1 U5225 ( .A(ram[2043]), .B(n10956), .Y(n6712) );
  AND2X1 U5226 ( .A(ram[2044]), .B(n10956), .Y(n6713) );
  AND2X1 U5227 ( .A(ram[2045]), .B(n10956), .Y(n6714) );
  AND2X1 U5228 ( .A(ram[2046]), .B(n10956), .Y(n6715) );
  AND2X1 U5229 ( .A(ram[1984]), .B(n10956), .Y(n6653) );
  AND2X1 U5230 ( .A(ram[1985]), .B(n10956), .Y(n6654) );
  AND2X1 U5231 ( .A(ram[1986]), .B(n10956), .Y(n6655) );
  AND2X1 U5232 ( .A(ram[1987]), .B(n10956), .Y(n6656) );
  AND2X1 U5233 ( .A(ram[1988]), .B(n10956), .Y(n6657) );
  AND2X1 U5234 ( .A(ram[1989]), .B(n10956), .Y(n6658) );
  AND2X1 U5235 ( .A(ram[1990]), .B(n10956), .Y(n6659) );
  AND2X1 U5236 ( .A(ram[2047]), .B(n10956), .Y(n6716) );
  MUX2X1 U5237 ( .B(n2159), .A(n2160), .S(n4183), .Y(n2158) );
  MUX2X1 U5238 ( .B(n2162), .A(n2163), .S(n4183), .Y(n2161) );
  MUX2X1 U5239 ( .B(n2165), .A(n2166), .S(n4183), .Y(n2164) );
  MUX2X1 U5240 ( .B(n2168), .A(n2169), .S(n4183), .Y(n2167) );
  MUX2X1 U5241 ( .B(n2171), .A(n2172), .S(n4153), .Y(n2170) );
  MUX2X1 U5242 ( .B(n2174), .A(n2175), .S(n4183), .Y(n2173) );
  MUX2X1 U5243 ( .B(n2177), .A(n2178), .S(n4183), .Y(n2176) );
  MUX2X1 U5244 ( .B(n2180), .A(n2181), .S(n4183), .Y(n2179) );
  MUX2X1 U5245 ( .B(n2183), .A(n2184), .S(n4183), .Y(n2182) );
  MUX2X1 U5246 ( .B(n2186), .A(n2187), .S(n4153), .Y(n2185) );
  MUX2X1 U5247 ( .B(n2189), .A(n2190), .S(n4184), .Y(n2188) );
  MUX2X1 U5248 ( .B(n2192), .A(n2193), .S(n4184), .Y(n2191) );
  MUX2X1 U5249 ( .B(n2195), .A(n2196), .S(n4184), .Y(n2194) );
  MUX2X1 U5250 ( .B(n2198), .A(n2199), .S(n4184), .Y(n2197) );
  MUX2X1 U5251 ( .B(n2201), .A(n2202), .S(n4153), .Y(n2200) );
  MUX2X1 U5252 ( .B(n2204), .A(n2205), .S(n4184), .Y(n2203) );
  MUX2X1 U5253 ( .B(n2207), .A(n2208), .S(n4184), .Y(n2206) );
  MUX2X1 U5254 ( .B(n2210), .A(n2211), .S(n4184), .Y(n2209) );
  MUX2X1 U5255 ( .B(n2213), .A(n2214), .S(n4184), .Y(n2212) );
  MUX2X1 U5256 ( .B(n2216), .A(n2217), .S(n4155), .Y(n2215) );
  MUX2X1 U5257 ( .B(n2219), .A(n2220), .S(n4184), .Y(n2218) );
  MUX2X1 U5258 ( .B(n2222), .A(n2223), .S(n4184), .Y(n2221) );
  MUX2X1 U5259 ( .B(n2225), .A(n2226), .S(n4184), .Y(n2224) );
  MUX2X1 U5260 ( .B(n2228), .A(n2229), .S(n4184), .Y(n2227) );
  MUX2X1 U5261 ( .B(n2231), .A(n2232), .S(n4155), .Y(n2230) );
  MUX2X1 U5262 ( .B(n2234), .A(n2235), .S(n4185), .Y(n2233) );
  MUX2X1 U5263 ( .B(n2237), .A(n2238), .S(n4185), .Y(n2236) );
  MUX2X1 U5264 ( .B(n2240), .A(n2241), .S(n4185), .Y(n2239) );
  MUX2X1 U5265 ( .B(n2243), .A(n2244), .S(n4185), .Y(n2242) );
  MUX2X1 U5266 ( .B(n2246), .A(n2247), .S(n4155), .Y(n2245) );
  MUX2X1 U5267 ( .B(n2249), .A(n2250), .S(n4185), .Y(n2248) );
  MUX2X1 U5268 ( .B(n2252), .A(n2253), .S(n4185), .Y(n2251) );
  MUX2X1 U5269 ( .B(n2255), .A(n2256), .S(n4185), .Y(n2254) );
  MUX2X1 U5270 ( .B(n2258), .A(n2259), .S(n4185), .Y(n2257) );
  MUX2X1 U5271 ( .B(n2261), .A(n2262), .S(n4156), .Y(n2260) );
  MUX2X1 U5272 ( .B(n2264), .A(n2265), .S(n4185), .Y(n2263) );
  MUX2X1 U5273 ( .B(n2267), .A(n2268), .S(n4185), .Y(n2266) );
  MUX2X1 U5274 ( .B(n2270), .A(n2271), .S(n4185), .Y(n2269) );
  MUX2X1 U5275 ( .B(n2273), .A(n2274), .S(n4185), .Y(n2272) );
  MUX2X1 U5276 ( .B(n2276), .A(n2277), .S(n4154), .Y(n2275) );
  MUX2X1 U5277 ( .B(n2279), .A(n2280), .S(n4186), .Y(n2278) );
  MUX2X1 U5278 ( .B(n2282), .A(n2283), .S(n4186), .Y(n2281) );
  MUX2X1 U5279 ( .B(n2285), .A(n2286), .S(n4186), .Y(n2284) );
  MUX2X1 U5280 ( .B(n2288), .A(n2289), .S(n4186), .Y(n2287) );
  MUX2X1 U5281 ( .B(n2291), .A(n2292), .S(n4153), .Y(n2290) );
  MUX2X1 U5282 ( .B(n2294), .A(n2295), .S(n4186), .Y(n2293) );
  MUX2X1 U5283 ( .B(n2297), .A(n2298), .S(n4186), .Y(n2296) );
  MUX2X1 U5284 ( .B(n2300), .A(n2301), .S(n4186), .Y(n2299) );
  MUX2X1 U5285 ( .B(n2303), .A(n2304), .S(n4186), .Y(n2302) );
  MUX2X1 U5286 ( .B(n2306), .A(n2307), .S(n4153), .Y(n2305) );
  MUX2X1 U5287 ( .B(n2309), .A(n2310), .S(n4186), .Y(n2308) );
  MUX2X1 U5288 ( .B(n2312), .A(n2313), .S(n4186), .Y(n2311) );
  MUX2X1 U5289 ( .B(n2315), .A(n2316), .S(n4186), .Y(n2314) );
  MUX2X1 U5290 ( .B(n2318), .A(n2319), .S(n4186), .Y(n2317) );
  MUX2X1 U5291 ( .B(n2321), .A(n2322), .S(n4155), .Y(n2320) );
  MUX2X1 U5292 ( .B(n2324), .A(n2325), .S(n4187), .Y(n2323) );
  MUX2X1 U5293 ( .B(n2327), .A(n2328), .S(n4187), .Y(n2326) );
  MUX2X1 U5294 ( .B(n2330), .A(n2331), .S(n4187), .Y(n2329) );
  MUX2X1 U5295 ( .B(n2333), .A(n2334), .S(n4187), .Y(n2332) );
  MUX2X1 U5296 ( .B(n2336), .A(n2337), .S(n4153), .Y(n2335) );
  MUX2X1 U5297 ( .B(n2339), .A(n2340), .S(n4187), .Y(n2338) );
  MUX2X1 U5298 ( .B(n2342), .A(n2343), .S(n4187), .Y(n2341) );
  MUX2X1 U5299 ( .B(n2345), .A(n2346), .S(n4187), .Y(n2344) );
  MUX2X1 U5300 ( .B(n2348), .A(n2349), .S(n4187), .Y(n2347) );
  MUX2X1 U5301 ( .B(n2351), .A(n2352), .S(n4154), .Y(n2350) );
  MUX2X1 U5302 ( .B(n2354), .A(n2355), .S(n4187), .Y(n2353) );
  MUX2X1 U5303 ( .B(n2357), .A(n2358), .S(n4187), .Y(n2356) );
  MUX2X1 U5304 ( .B(n2360), .A(n2361), .S(n4187), .Y(n2359) );
  MUX2X1 U5305 ( .B(n2363), .A(n2364), .S(n4187), .Y(n2362) );
  MUX2X1 U5306 ( .B(n2366), .A(n2367), .S(n4156), .Y(n2365) );
  MUX2X1 U5307 ( .B(n2369), .A(n2370), .S(n4188), .Y(n2368) );
  MUX2X1 U5308 ( .B(n2372), .A(n2373), .S(n4188), .Y(n2371) );
  MUX2X1 U5309 ( .B(n2375), .A(n2376), .S(n4188), .Y(n2374) );
  MUX2X1 U5310 ( .B(n2378), .A(n2379), .S(n4188), .Y(n2377) );
  MUX2X1 U5311 ( .B(n2381), .A(n2382), .S(n4154), .Y(n2380) );
  MUX2X1 U5312 ( .B(n2384), .A(n2385), .S(n4188), .Y(n2383) );
  MUX2X1 U5313 ( .B(n2387), .A(n2388), .S(n4188), .Y(n2386) );
  MUX2X1 U5314 ( .B(n2390), .A(n2391), .S(n4188), .Y(n2389) );
  MUX2X1 U5315 ( .B(n2393), .A(n2394), .S(n4188), .Y(n2392) );
  MUX2X1 U5316 ( .B(n2396), .A(n2397), .S(n4154), .Y(n2395) );
  MUX2X1 U5317 ( .B(n2399), .A(n2400), .S(n4188), .Y(n2398) );
  MUX2X1 U5318 ( .B(n2402), .A(n2403), .S(n4188), .Y(n2401) );
  MUX2X1 U5319 ( .B(n2405), .A(n2406), .S(n4188), .Y(n2404) );
  MUX2X1 U5320 ( .B(n2408), .A(n2409), .S(n4188), .Y(n2407) );
  MUX2X1 U5321 ( .B(n2411), .A(n2412), .S(n4155), .Y(n2410) );
  MUX2X1 U5322 ( .B(n2414), .A(n2415), .S(n4189), .Y(n2413) );
  MUX2X1 U5323 ( .B(n2417), .A(n2418), .S(n4189), .Y(n2416) );
  MUX2X1 U5324 ( .B(n2420), .A(n2421), .S(n4189), .Y(n2419) );
  MUX2X1 U5325 ( .B(n2423), .A(n2424), .S(n4189), .Y(n2422) );
  MUX2X1 U5326 ( .B(n2426), .A(n2427), .S(n4153), .Y(n2425) );
  MUX2X1 U5327 ( .B(n2429), .A(n2430), .S(n4189), .Y(n2428) );
  MUX2X1 U5328 ( .B(n2432), .A(n2433), .S(n4189), .Y(n2431) );
  MUX2X1 U5329 ( .B(n2435), .A(n2436), .S(n4189), .Y(n2434) );
  MUX2X1 U5330 ( .B(n2438), .A(n2439), .S(n4189), .Y(n2437) );
  MUX2X1 U5331 ( .B(n2441), .A(n2442), .S(n4156), .Y(n2440) );
  MUX2X1 U5332 ( .B(n2444), .A(n2445), .S(n4189), .Y(n2443) );
  MUX2X1 U5333 ( .B(n2447), .A(n2448), .S(n4189), .Y(n2446) );
  MUX2X1 U5334 ( .B(n2450), .A(n2451), .S(n4189), .Y(n2449) );
  MUX2X1 U5335 ( .B(n2453), .A(n2454), .S(n4189), .Y(n2452) );
  MUX2X1 U5336 ( .B(n2456), .A(n2457), .S(n4156), .Y(n2455) );
  MUX2X1 U5337 ( .B(n2459), .A(n2460), .S(n4190), .Y(n2458) );
  MUX2X1 U5338 ( .B(n2462), .A(n2463), .S(n4190), .Y(n2461) );
  MUX2X1 U5339 ( .B(n2465), .A(n2466), .S(n4190), .Y(n2464) );
  MUX2X1 U5340 ( .B(n2468), .A(n2469), .S(n4190), .Y(n2467) );
  MUX2X1 U5341 ( .B(n2471), .A(n2472), .S(n4157), .Y(n2470) );
  MUX2X1 U5342 ( .B(n2474), .A(n2475), .S(n4190), .Y(n2473) );
  MUX2X1 U5343 ( .B(n2477), .A(n2478), .S(n4190), .Y(n2476) );
  MUX2X1 U5344 ( .B(n2480), .A(n2481), .S(n4190), .Y(n2479) );
  MUX2X1 U5345 ( .B(n2483), .A(n2484), .S(n4190), .Y(n2482) );
  MUX2X1 U5346 ( .B(n2486), .A(n2487), .S(n4157), .Y(n2485) );
  MUX2X1 U5347 ( .B(n2489), .A(n2490), .S(n4190), .Y(n2488) );
  MUX2X1 U5348 ( .B(n2492), .A(n2493), .S(n4190), .Y(n2491) );
  MUX2X1 U5349 ( .B(n2495), .A(n2496), .S(n4190), .Y(n2494) );
  MUX2X1 U5350 ( .B(n2498), .A(n2499), .S(n4190), .Y(n2497) );
  MUX2X1 U5351 ( .B(n2501), .A(n2502), .S(n4157), .Y(n2500) );
  MUX2X1 U5352 ( .B(n2504), .A(n2505), .S(n4191), .Y(n2503) );
  MUX2X1 U5353 ( .B(n2507), .A(n2508), .S(n4191), .Y(n2506) );
  MUX2X1 U5354 ( .B(n2510), .A(n2511), .S(n4191), .Y(n2509) );
  MUX2X1 U5355 ( .B(n2513), .A(n2514), .S(n4191), .Y(n2512) );
  MUX2X1 U5356 ( .B(n2516), .A(n2518), .S(n4157), .Y(n2515) );
  MUX2X1 U5357 ( .B(n2520), .A(n2521), .S(n4191), .Y(n2519) );
  MUX2X1 U5358 ( .B(n2523), .A(n2524), .S(n4191), .Y(n2522) );
  MUX2X1 U5359 ( .B(n2526), .A(n2527), .S(n4191), .Y(n2525) );
  MUX2X1 U5360 ( .B(n2529), .A(n2530), .S(n4191), .Y(n2528) );
  MUX2X1 U5361 ( .B(n2532), .A(n2533), .S(n4157), .Y(n2531) );
  MUX2X1 U5362 ( .B(n2535), .A(n2536), .S(n4191), .Y(n2534) );
  MUX2X1 U5363 ( .B(n2538), .A(n2539), .S(n4191), .Y(n2537) );
  MUX2X1 U5364 ( .B(n2541), .A(n2542), .S(n4191), .Y(n2540) );
  MUX2X1 U5365 ( .B(n2544), .A(n2545), .S(n4191), .Y(n2543) );
  MUX2X1 U5366 ( .B(n2547), .A(n2548), .S(n4157), .Y(n2546) );
  MUX2X1 U5367 ( .B(n2550), .A(n2551), .S(n4192), .Y(n2549) );
  MUX2X1 U5368 ( .B(n2553), .A(n2554), .S(n4192), .Y(n2552) );
  MUX2X1 U5369 ( .B(n2556), .A(n2557), .S(n4192), .Y(n2555) );
  MUX2X1 U5370 ( .B(n2559), .A(n2560), .S(n4192), .Y(n2558) );
  MUX2X1 U5371 ( .B(n2562), .A(n2563), .S(n4157), .Y(n2561) );
  MUX2X1 U5372 ( .B(n2565), .A(n2566), .S(n4192), .Y(n2564) );
  MUX2X1 U5373 ( .B(n2568), .A(n2569), .S(n4192), .Y(n2567) );
  MUX2X1 U5374 ( .B(n2571), .A(n2572), .S(n4192), .Y(n2570) );
  MUX2X1 U5375 ( .B(n2574), .A(n2575), .S(n4192), .Y(n2573) );
  MUX2X1 U5376 ( .B(n2577), .A(n2578), .S(n4157), .Y(n2576) );
  MUX2X1 U5377 ( .B(n2580), .A(n2581), .S(n4192), .Y(n2579) );
  MUX2X1 U5378 ( .B(n2583), .A(n2585), .S(n4192), .Y(n2582) );
  MUX2X1 U5379 ( .B(n2587), .A(n2588), .S(n4192), .Y(n2586) );
  MUX2X1 U5380 ( .B(n2590), .A(n2591), .S(n4192), .Y(n2589) );
  MUX2X1 U5381 ( .B(n2593), .A(n2594), .S(n4157), .Y(n2592) );
  MUX2X1 U5382 ( .B(n2596), .A(n2597), .S(n4193), .Y(n2595) );
  MUX2X1 U5383 ( .B(n2599), .A(n2600), .S(n4193), .Y(n2598) );
  MUX2X1 U5384 ( .B(n2602), .A(n2603), .S(n4193), .Y(n2601) );
  MUX2X1 U5385 ( .B(n2605), .A(n2606), .S(n4193), .Y(n2604) );
  MUX2X1 U5386 ( .B(n2608), .A(n2609), .S(n4157), .Y(n2607) );
  MUX2X1 U5387 ( .B(n2611), .A(n2612), .S(n4193), .Y(n2610) );
  MUX2X1 U5388 ( .B(n2614), .A(n2615), .S(n4193), .Y(n2613) );
  MUX2X1 U5389 ( .B(n2617), .A(n2618), .S(n4193), .Y(n2616) );
  MUX2X1 U5390 ( .B(n2620), .A(n2621), .S(n4193), .Y(n2619) );
  MUX2X1 U5391 ( .B(n2623), .A(n2624), .S(n10963), .Y(n2622) );
  MUX2X1 U5392 ( .B(n2626), .A(n2627), .S(n4193), .Y(n2625) );
  MUX2X1 U5393 ( .B(n2629), .A(n2630), .S(n4193), .Y(n2628) );
  MUX2X1 U5394 ( .B(n2632), .A(n2633), .S(n4193), .Y(n2631) );
  MUX2X1 U5395 ( .B(n2635), .A(n2636), .S(n4193), .Y(n2634) );
  MUX2X1 U5396 ( .B(n2638), .A(n2639), .S(n4157), .Y(n2637) );
  MUX2X1 U5397 ( .B(n2641), .A(n2642), .S(n4194), .Y(n2640) );
  MUX2X1 U5398 ( .B(n2644), .A(n2645), .S(n4194), .Y(n2643) );
  MUX2X1 U5399 ( .B(n2647), .A(n2648), .S(n4194), .Y(n2646) );
  MUX2X1 U5400 ( .B(n2650), .A(n2652), .S(n4194), .Y(n2649) );
  MUX2X1 U5401 ( .B(n2654), .A(n2655), .S(n4156), .Y(n2653) );
  MUX2X1 U5402 ( .B(n2657), .A(n2658), .S(n4194), .Y(n2656) );
  MUX2X1 U5403 ( .B(n2660), .A(n2661), .S(n4194), .Y(n2659) );
  MUX2X1 U5404 ( .B(n2663), .A(n2664), .S(n4194), .Y(n2662) );
  MUX2X1 U5405 ( .B(n2666), .A(n2667), .S(n4194), .Y(n2665) );
  MUX2X1 U5406 ( .B(n2669), .A(n2670), .S(n4154), .Y(n2668) );
  MUX2X1 U5407 ( .B(n2672), .A(n2673), .S(n4194), .Y(n2671) );
  MUX2X1 U5408 ( .B(n2675), .A(n2676), .S(n4194), .Y(n2674) );
  MUX2X1 U5409 ( .B(n2678), .A(n2679), .S(n4194), .Y(n2677) );
  MUX2X1 U5410 ( .B(n2681), .A(n2682), .S(n4194), .Y(n2680) );
  MUX2X1 U5411 ( .B(n2684), .A(n2685), .S(n4157), .Y(n2683) );
  MUX2X1 U5412 ( .B(n2687), .A(n2688), .S(n4195), .Y(n2686) );
  MUX2X1 U5413 ( .B(n2690), .A(n2691), .S(n4195), .Y(n2689) );
  MUX2X1 U5414 ( .B(n2693), .A(n2694), .S(n4195), .Y(n2692) );
  MUX2X1 U5415 ( .B(n2696), .A(n2697), .S(n4195), .Y(n2695) );
  MUX2X1 U5416 ( .B(n2699), .A(n2700), .S(n4157), .Y(n2698) );
  MUX2X1 U5417 ( .B(n2702), .A(n2703), .S(n4195), .Y(n2701) );
  MUX2X1 U5418 ( .B(n2705), .A(n2706), .S(n4195), .Y(n2704) );
  MUX2X1 U5419 ( .B(n2708), .A(n2709), .S(n4195), .Y(n2707) );
  MUX2X1 U5420 ( .B(n2711), .A(n2712), .S(n4195), .Y(n2710) );
  MUX2X1 U5421 ( .B(n2714), .A(n2715), .S(n4155), .Y(n2713) );
  MUX2X1 U5422 ( .B(n2717), .A(n2719), .S(n4195), .Y(n2716) );
  MUX2X1 U5423 ( .B(n2721), .A(n2722), .S(n4195), .Y(n2720) );
  MUX2X1 U5424 ( .B(n2724), .A(n2725), .S(n4195), .Y(n2723) );
  MUX2X1 U5425 ( .B(n2727), .A(n2728), .S(n4195), .Y(n2726) );
  MUX2X1 U5426 ( .B(n2730), .A(n2731), .S(n4157), .Y(n2729) );
  MUX2X1 U5427 ( .B(n2733), .A(n2734), .S(n4196), .Y(n2732) );
  MUX2X1 U5428 ( .B(n2736), .A(n2737), .S(n4196), .Y(n2735) );
  MUX2X1 U5429 ( .B(n2739), .A(n2740), .S(n4196), .Y(n2738) );
  MUX2X1 U5430 ( .B(n2742), .A(n2743), .S(n4196), .Y(n2741) );
  MUX2X1 U5431 ( .B(n2745), .A(n2746), .S(n4156), .Y(n2744) );
  MUX2X1 U5432 ( .B(n2748), .A(n2749), .S(n4196), .Y(n2747) );
  MUX2X1 U5433 ( .B(n2751), .A(n2752), .S(n4196), .Y(n2750) );
  MUX2X1 U5434 ( .B(n2754), .A(n2755), .S(n4196), .Y(n2753) );
  MUX2X1 U5435 ( .B(n2757), .A(n2758), .S(n4196), .Y(n2756) );
  MUX2X1 U5436 ( .B(n2760), .A(n2761), .S(n4154), .Y(n2759) );
  MUX2X1 U5437 ( .B(n2763), .A(n2764), .S(n4196), .Y(n2762) );
  MUX2X1 U5438 ( .B(n2766), .A(n2767), .S(n4196), .Y(n2765) );
  MUX2X1 U5439 ( .B(n2769), .A(n2770), .S(n4196), .Y(n2768) );
  MUX2X1 U5440 ( .B(n2772), .A(n2773), .S(n4196), .Y(n2771) );
  MUX2X1 U5441 ( .B(n2775), .A(n2776), .S(n4156), .Y(n2774) );
  MUX2X1 U5442 ( .B(n2778), .A(n2779), .S(n4197), .Y(n2777) );
  MUX2X1 U5443 ( .B(n2781), .A(n2782), .S(n4197), .Y(n2780) );
  MUX2X1 U5444 ( .B(n2784), .A(n2786), .S(n4197), .Y(n2783) );
  MUX2X1 U5445 ( .B(n2788), .A(n2789), .S(n4197), .Y(n2787) );
  MUX2X1 U5446 ( .B(n2791), .A(n2792), .S(n4157), .Y(n2790) );
  MUX2X1 U5447 ( .B(n2794), .A(n2795), .S(n4197), .Y(n2793) );
  MUX2X1 U5448 ( .B(n2797), .A(n2798), .S(n4197), .Y(n2796) );
  MUX2X1 U5449 ( .B(n2800), .A(n2801), .S(n4197), .Y(n2799) );
  MUX2X1 U5450 ( .B(n2803), .A(n2804), .S(n4197), .Y(n2802) );
  MUX2X1 U5451 ( .B(n2806), .A(n2807), .S(n4154), .Y(n2805) );
  MUX2X1 U5452 ( .B(n2809), .A(n2810), .S(n4197), .Y(n2808) );
  MUX2X1 U5453 ( .B(n2812), .A(n2813), .S(n4197), .Y(n2811) );
  MUX2X1 U5454 ( .B(n2815), .A(n2816), .S(n4197), .Y(n2814) );
  MUX2X1 U5455 ( .B(n2818), .A(n2819), .S(n4197), .Y(n2817) );
  MUX2X1 U5456 ( .B(n2821), .A(n2822), .S(n4157), .Y(n2820) );
  MUX2X1 U5457 ( .B(n2824), .A(n2825), .S(n4198), .Y(n2823) );
  MUX2X1 U5458 ( .B(n2827), .A(n2828), .S(n4198), .Y(n2826) );
  MUX2X1 U5459 ( .B(n2830), .A(n2831), .S(n4198), .Y(n2829) );
  MUX2X1 U5460 ( .B(n2833), .A(n2834), .S(n4198), .Y(n2832) );
  MUX2X1 U5461 ( .B(n2836), .A(n2837), .S(n4153), .Y(n2835) );
  MUX2X1 U5462 ( .B(n2839), .A(n2840), .S(n4198), .Y(n2838) );
  MUX2X1 U5463 ( .B(n2842), .A(n2843), .S(n4198), .Y(n2841) );
  MUX2X1 U5464 ( .B(n2845), .A(n2846), .S(n4198), .Y(n2844) );
  MUX2X1 U5465 ( .B(n2848), .A(n2849), .S(n4198), .Y(n2847) );
  MUX2X1 U5466 ( .B(n2851), .A(n2853), .S(n4153), .Y(n2850) );
  MUX2X1 U5467 ( .B(n2855), .A(n2856), .S(n4198), .Y(n2854) );
  MUX2X1 U5468 ( .B(n2858), .A(n2859), .S(n4198), .Y(n2857) );
  MUX2X1 U5469 ( .B(n2861), .A(n2862), .S(n4198), .Y(n2860) );
  MUX2X1 U5470 ( .B(n2864), .A(n2865), .S(n4198), .Y(n2863) );
  MUX2X1 U5471 ( .B(n2867), .A(n2868), .S(n4153), .Y(n2866) );
  MUX2X1 U5472 ( .B(n2870), .A(n2871), .S(n4199), .Y(n2869) );
  MUX2X1 U5473 ( .B(n2873), .A(n2874), .S(n4199), .Y(n2872) );
  MUX2X1 U5474 ( .B(n2876), .A(n2877), .S(n4199), .Y(n2875) );
  MUX2X1 U5475 ( .B(n2879), .A(n2880), .S(n4199), .Y(n2878) );
  MUX2X1 U5476 ( .B(n2882), .A(n2883), .S(n4153), .Y(n2881) );
  MUX2X1 U5477 ( .B(n2885), .A(n2886), .S(n4199), .Y(n2884) );
  MUX2X1 U5478 ( .B(n2888), .A(n2889), .S(n4199), .Y(n2887) );
  MUX2X1 U5479 ( .B(n2891), .A(n2892), .S(n4199), .Y(n2890) );
  MUX2X1 U5480 ( .B(n2894), .A(n2895), .S(n4199), .Y(n2893) );
  MUX2X1 U5481 ( .B(n2897), .A(n2898), .S(n4153), .Y(n2896) );
  MUX2X1 U5482 ( .B(n2900), .A(n2901), .S(n4199), .Y(n2899) );
  MUX2X1 U5483 ( .B(n2903), .A(n2904), .S(n4199), .Y(n2902) );
  MUX2X1 U5484 ( .B(n2906), .A(n2907), .S(n4199), .Y(n2905) );
  MUX2X1 U5485 ( .B(n2909), .A(n2910), .S(n4199), .Y(n2908) );
  MUX2X1 U5486 ( .B(n2912), .A(n2913), .S(n4153), .Y(n2911) );
  MUX2X1 U5487 ( .B(n2915), .A(n2916), .S(n4200), .Y(n2914) );
  MUX2X1 U5488 ( .B(n2918), .A(n2920), .S(n4200), .Y(n2917) );
  MUX2X1 U5489 ( .B(n2922), .A(n2923), .S(n4200), .Y(n2921) );
  MUX2X1 U5490 ( .B(n2925), .A(n2926), .S(n4200), .Y(n2924) );
  MUX2X1 U5491 ( .B(n2928), .A(n2929), .S(n4153), .Y(n2927) );
  MUX2X1 U5492 ( .B(n2931), .A(n2932), .S(n4200), .Y(n2930) );
  MUX2X1 U5493 ( .B(n2934), .A(n2935), .S(n4200), .Y(n2933) );
  MUX2X1 U5494 ( .B(n2937), .A(n2938), .S(n4200), .Y(n2936) );
  MUX2X1 U5495 ( .B(n2940), .A(n2941), .S(n4200), .Y(n2939) );
  MUX2X1 U5496 ( .B(n2943), .A(n2944), .S(n4153), .Y(n2942) );
  MUX2X1 U5497 ( .B(n2946), .A(n2947), .S(n4200), .Y(n2945) );
  MUX2X1 U5498 ( .B(n2949), .A(n2950), .S(n4200), .Y(n2948) );
  MUX2X1 U5499 ( .B(n2952), .A(n2953), .S(n4200), .Y(n2951) );
  MUX2X1 U5500 ( .B(n2955), .A(n2956), .S(n4200), .Y(n2954) );
  MUX2X1 U5501 ( .B(n2958), .A(n2959), .S(n4153), .Y(n2957) );
  MUX2X1 U5502 ( .B(n2961), .A(n2962), .S(n4201), .Y(n2960) );
  MUX2X1 U5503 ( .B(n2964), .A(n2965), .S(n4201), .Y(n2963) );
  MUX2X1 U5504 ( .B(n2967), .A(n2968), .S(n4201), .Y(n2966) );
  MUX2X1 U5505 ( .B(n2970), .A(n2971), .S(n4201), .Y(n2969) );
  MUX2X1 U5506 ( .B(n2973), .A(n2974), .S(n4153), .Y(n2972) );
  MUX2X1 U5507 ( .B(n2976), .A(n2977), .S(n4201), .Y(n2975) );
  MUX2X1 U5508 ( .B(n2979), .A(n2980), .S(n4201), .Y(n2978) );
  MUX2X1 U5509 ( .B(n2982), .A(n2983), .S(n4201), .Y(n2981) );
  MUX2X1 U5510 ( .B(n2985), .A(n2987), .S(n4201), .Y(n2984) );
  MUX2X1 U5511 ( .B(n2989), .A(n2990), .S(n4153), .Y(n2988) );
  MUX2X1 U5512 ( .B(n2992), .A(n2993), .S(n4201), .Y(n2991) );
  MUX2X1 U5513 ( .B(n2995), .A(n2996), .S(n4201), .Y(n2994) );
  MUX2X1 U5514 ( .B(n2998), .A(n2999), .S(n4201), .Y(n2997) );
  MUX2X1 U5515 ( .B(n3001), .A(n3002), .S(n4201), .Y(n3000) );
  MUX2X1 U5516 ( .B(n3004), .A(n3005), .S(n4153), .Y(n3003) );
  MUX2X1 U5517 ( .B(n3007), .A(n3008), .S(n4202), .Y(n3006) );
  MUX2X1 U5518 ( .B(n3010), .A(n3011), .S(n4202), .Y(n3009) );
  MUX2X1 U5519 ( .B(n3013), .A(n3014), .S(n4202), .Y(n3012) );
  MUX2X1 U5520 ( .B(n3016), .A(n3017), .S(n4202), .Y(n3015) );
  MUX2X1 U5521 ( .B(n3019), .A(n3020), .S(n4154), .Y(n3018) );
  MUX2X1 U5522 ( .B(n3022), .A(n3023), .S(n4202), .Y(n3021) );
  MUX2X1 U5523 ( .B(n3025), .A(n3026), .S(n4202), .Y(n3024) );
  MUX2X1 U5524 ( .B(n3028), .A(n3029), .S(n4202), .Y(n3027) );
  MUX2X1 U5525 ( .B(n3031), .A(n3032), .S(n4202), .Y(n3030) );
  MUX2X1 U5526 ( .B(n3034), .A(n3035), .S(n4155), .Y(n3033) );
  MUX2X1 U5527 ( .B(n3037), .A(n3038), .S(n4202), .Y(n3036) );
  MUX2X1 U5528 ( .B(n3040), .A(n3041), .S(n4202), .Y(n3039) );
  MUX2X1 U5529 ( .B(n3043), .A(n3044), .S(n4202), .Y(n3042) );
  MUX2X1 U5530 ( .B(n3046), .A(n3047), .S(n4202), .Y(n3045) );
  MUX2X1 U5531 ( .B(n3049), .A(n3050), .S(n4153), .Y(n3048) );
  MUX2X1 U5532 ( .B(n3052), .A(n3053), .S(n4203), .Y(n3051) );
  MUX2X1 U5533 ( .B(n3055), .A(n3056), .S(n4203), .Y(n3054) );
  MUX2X1 U5534 ( .B(n3058), .A(n3059), .S(n4203), .Y(n3057) );
  MUX2X1 U5535 ( .B(n3061), .A(n3062), .S(n4203), .Y(n3060) );
  MUX2X1 U5536 ( .B(n3064), .A(n3065), .S(n4156), .Y(n3063) );
  MUX2X1 U5537 ( .B(n3067), .A(n3068), .S(n4203), .Y(n3066) );
  MUX2X1 U5538 ( .B(n3070), .A(n3071), .S(n4203), .Y(n3069) );
  MUX2X1 U5539 ( .B(n3073), .A(n3074), .S(n4203), .Y(n3072) );
  MUX2X1 U5540 ( .B(n3076), .A(n3077), .S(n4203), .Y(n3075) );
  MUX2X1 U5541 ( .B(n3079), .A(n3080), .S(n4155), .Y(n3078) );
  MUX2X1 U5542 ( .B(n3082), .A(n3083), .S(n4203), .Y(n3081) );
  MUX2X1 U5543 ( .B(n3085), .A(n3086), .S(n4203), .Y(n3084) );
  MUX2X1 U5544 ( .B(n3088), .A(n3089), .S(n4203), .Y(n3087) );
  MUX2X1 U5545 ( .B(n3091), .A(n3092), .S(n4203), .Y(n3090) );
  MUX2X1 U5546 ( .B(n3094), .A(n3095), .S(n4154), .Y(n3093) );
  MUX2X1 U5547 ( .B(n3097), .A(n3098), .S(n4204), .Y(n3096) );
  MUX2X1 U5548 ( .B(n3100), .A(n3101), .S(n4204), .Y(n3099) );
  MUX2X1 U5549 ( .B(n3103), .A(n3104), .S(n4204), .Y(n3102) );
  MUX2X1 U5550 ( .B(n3106), .A(n3107), .S(n4204), .Y(n3105) );
  MUX2X1 U5551 ( .B(n3109), .A(n3110), .S(n4153), .Y(n3108) );
  MUX2X1 U5552 ( .B(n3112), .A(n3113), .S(n4204), .Y(n3111) );
  MUX2X1 U5553 ( .B(n3115), .A(n3116), .S(n4204), .Y(n3114) );
  MUX2X1 U5554 ( .B(n3118), .A(n3119), .S(n4204), .Y(n3117) );
  MUX2X1 U5555 ( .B(n3121), .A(n3122), .S(n4204), .Y(n3120) );
  MUX2X1 U5556 ( .B(n3124), .A(n3125), .S(n4156), .Y(n3123) );
  MUX2X1 U5557 ( .B(n3127), .A(n3128), .S(n4204), .Y(n3126) );
  MUX2X1 U5558 ( .B(n3130), .A(n3131), .S(n4204), .Y(n3129) );
  MUX2X1 U5559 ( .B(n3133), .A(n3134), .S(n4204), .Y(n3132) );
  MUX2X1 U5560 ( .B(n3136), .A(n3137), .S(n4204), .Y(n3135) );
  MUX2X1 U5561 ( .B(n3139), .A(n3140), .S(n4153), .Y(n3138) );
  MUX2X1 U5562 ( .B(n3142), .A(n3143), .S(n4205), .Y(n3141) );
  MUX2X1 U5563 ( .B(n3145), .A(n3146), .S(n4205), .Y(n3144) );
  MUX2X1 U5564 ( .B(n3148), .A(n3149), .S(n4205), .Y(n3147) );
  MUX2X1 U5565 ( .B(n3151), .A(n3152), .S(n4205), .Y(n3150) );
  MUX2X1 U5566 ( .B(n3154), .A(n3155), .S(n4154), .Y(n3153) );
  MUX2X1 U5567 ( .B(n3157), .A(n3158), .S(n4205), .Y(n3156) );
  MUX2X1 U5568 ( .B(n3160), .A(n3161), .S(n4205), .Y(n3159) );
  MUX2X1 U5569 ( .B(n3163), .A(n3164), .S(n4205), .Y(n3162) );
  MUX2X1 U5570 ( .B(n3166), .A(n3167), .S(n4205), .Y(n3165) );
  MUX2X1 U5571 ( .B(n3169), .A(n3170), .S(n4156), .Y(n3168) );
  MUX2X1 U5572 ( .B(n3172), .A(n3173), .S(n4205), .Y(n3171) );
  MUX2X1 U5573 ( .B(n3175), .A(n3176), .S(n4205), .Y(n3174) );
  MUX2X1 U5574 ( .B(n3178), .A(n3179), .S(n4205), .Y(n3177) );
  MUX2X1 U5575 ( .B(n3181), .A(n3182), .S(n4205), .Y(n3180) );
  MUX2X1 U5576 ( .B(n3184), .A(n3185), .S(n4154), .Y(n3183) );
  MUX2X1 U5577 ( .B(n3187), .A(n3188), .S(n4206), .Y(n3186) );
  MUX2X1 U5578 ( .B(n3190), .A(n3191), .S(n4206), .Y(n3189) );
  MUX2X1 U5579 ( .B(n3193), .A(n3194), .S(n4206), .Y(n3192) );
  MUX2X1 U5580 ( .B(n3196), .A(n3197), .S(n4206), .Y(n3195) );
  MUX2X1 U5581 ( .B(n3199), .A(n3200), .S(n4155), .Y(n3198) );
  MUX2X1 U5582 ( .B(n3202), .A(n3203), .S(n4206), .Y(n3201) );
  MUX2X1 U5583 ( .B(n3205), .A(n3206), .S(n4206), .Y(n3204) );
  MUX2X1 U5584 ( .B(n3208), .A(n3209), .S(n4206), .Y(n3207) );
  MUX2X1 U5585 ( .B(n3211), .A(n3212), .S(n4206), .Y(n3210) );
  MUX2X1 U5586 ( .B(n3214), .A(n3215), .S(n4155), .Y(n3213) );
  MUX2X1 U5587 ( .B(n3217), .A(n3218), .S(n4206), .Y(n3216) );
  MUX2X1 U5588 ( .B(n3220), .A(n3221), .S(n4206), .Y(n3219) );
  MUX2X1 U5589 ( .B(n3223), .A(n3224), .S(n4206), .Y(n3222) );
  MUX2X1 U5590 ( .B(n3226), .A(n3227), .S(n4206), .Y(n3225) );
  MUX2X1 U5591 ( .B(n3229), .A(n3230), .S(n4154), .Y(n3228) );
  MUX2X1 U5592 ( .B(n3232), .A(n3233), .S(n4207), .Y(n3231) );
  MUX2X1 U5593 ( .B(n3235), .A(n3236), .S(n4207), .Y(n3234) );
  MUX2X1 U5594 ( .B(n3238), .A(n3239), .S(n4207), .Y(n3237) );
  MUX2X1 U5595 ( .B(n3241), .A(n3242), .S(n4207), .Y(n3240) );
  MUX2X1 U5596 ( .B(n3244), .A(n3245), .S(n4154), .Y(n3243) );
  MUX2X1 U5597 ( .B(n3247), .A(n3248), .S(n4207), .Y(n3246) );
  MUX2X1 U5598 ( .B(n3250), .A(n3251), .S(n4207), .Y(n3249) );
  MUX2X1 U5599 ( .B(n3253), .A(n3254), .S(n4207), .Y(n3252) );
  MUX2X1 U5600 ( .B(n3256), .A(n3257), .S(n4207), .Y(n3255) );
  MUX2X1 U5601 ( .B(n3259), .A(n3260), .S(n4156), .Y(n3258) );
  MUX2X1 U5602 ( .B(n3262), .A(n3263), .S(n4207), .Y(n3261) );
  MUX2X1 U5603 ( .B(n3265), .A(n3266), .S(n4207), .Y(n3264) );
  MUX2X1 U5604 ( .B(n3268), .A(n3269), .S(n4207), .Y(n3267) );
  MUX2X1 U5605 ( .B(n3271), .A(n3272), .S(n4207), .Y(n3270) );
  MUX2X1 U5606 ( .B(n3274), .A(n3275), .S(n4156), .Y(n3273) );
  MUX2X1 U5607 ( .B(n3277), .A(n3278), .S(n4208), .Y(n3276) );
  MUX2X1 U5608 ( .B(n3280), .A(n3281), .S(n4208), .Y(n3279) );
  MUX2X1 U5609 ( .B(n3283), .A(n3284), .S(n4208), .Y(n3282) );
  MUX2X1 U5610 ( .B(n3286), .A(n3287), .S(n4208), .Y(n3285) );
  MUX2X1 U5611 ( .B(n3289), .A(n3290), .S(n4154), .Y(n3288) );
  MUX2X1 U5612 ( .B(n3292), .A(n3293), .S(n4208), .Y(n3291) );
  MUX2X1 U5613 ( .B(n3295), .A(n3296), .S(n4208), .Y(n3294) );
  MUX2X1 U5614 ( .B(n3298), .A(n3299), .S(n4208), .Y(n3297) );
  MUX2X1 U5615 ( .B(n3301), .A(n3302), .S(n4208), .Y(n3300) );
  MUX2X1 U5616 ( .B(n3304), .A(n3305), .S(n4156), .Y(n3303) );
  MUX2X1 U5617 ( .B(n3307), .A(n3308), .S(n4208), .Y(n3306) );
  MUX2X1 U5618 ( .B(n3310), .A(n3311), .S(n4208), .Y(n3309) );
  MUX2X1 U5619 ( .B(n3313), .A(n3314), .S(n4208), .Y(n3312) );
  MUX2X1 U5620 ( .B(n3316), .A(n3317), .S(n4208), .Y(n3315) );
  MUX2X1 U5621 ( .B(n3319), .A(n3320), .S(n4154), .Y(n3318) );
  MUX2X1 U5622 ( .B(n3322), .A(n3323), .S(n4209), .Y(n3321) );
  MUX2X1 U5623 ( .B(n3325), .A(n3326), .S(n4209), .Y(n3324) );
  MUX2X1 U5624 ( .B(n3328), .A(n3329), .S(n4209), .Y(n3327) );
  MUX2X1 U5625 ( .B(n3331), .A(n3332), .S(n4209), .Y(n3330) );
  MUX2X1 U5626 ( .B(n3334), .A(n3335), .S(n4156), .Y(n3333) );
  MUX2X1 U5627 ( .B(n3337), .A(n3338), .S(n4209), .Y(n3336) );
  MUX2X1 U5628 ( .B(n3340), .A(n3341), .S(n4209), .Y(n3339) );
  MUX2X1 U5629 ( .B(n3343), .A(n3344), .S(n4209), .Y(n3342) );
  MUX2X1 U5630 ( .B(n3346), .A(n3347), .S(n4209), .Y(n3345) );
  MUX2X1 U5631 ( .B(n3349), .A(n3350), .S(n4155), .Y(n3348) );
  MUX2X1 U5632 ( .B(n3352), .A(n3353), .S(n4209), .Y(n3351) );
  MUX2X1 U5633 ( .B(n3355), .A(n3356), .S(n4209), .Y(n3354) );
  MUX2X1 U5634 ( .B(n3358), .A(n3359), .S(n4209), .Y(n3357) );
  MUX2X1 U5635 ( .B(n3361), .A(n3362), .S(n4209), .Y(n3360) );
  MUX2X1 U5636 ( .B(n3364), .A(n3365), .S(n4156), .Y(n3363) );
  MUX2X1 U5637 ( .B(n3367), .A(n3368), .S(n4210), .Y(n3366) );
  MUX2X1 U5638 ( .B(n3370), .A(n3371), .S(n4210), .Y(n3369) );
  MUX2X1 U5639 ( .B(n3373), .A(n3374), .S(n4210), .Y(n3372) );
  MUX2X1 U5640 ( .B(n3376), .A(n3377), .S(n4210), .Y(n3375) );
  MUX2X1 U5641 ( .B(n3379), .A(n3380), .S(n4154), .Y(n3378) );
  MUX2X1 U5642 ( .B(n3382), .A(n3383), .S(n4210), .Y(n3381) );
  MUX2X1 U5643 ( .B(n3385), .A(n3386), .S(n4210), .Y(n3384) );
  MUX2X1 U5644 ( .B(n3388), .A(n3389), .S(n4210), .Y(n3387) );
  MUX2X1 U5645 ( .B(n3391), .A(n3392), .S(n4210), .Y(n3390) );
  MUX2X1 U5646 ( .B(n3394), .A(n3395), .S(n4154), .Y(n3393) );
  MUX2X1 U5647 ( .B(n3397), .A(n3398), .S(n4210), .Y(n3396) );
  MUX2X1 U5648 ( .B(n3400), .A(n3401), .S(n4210), .Y(n3399) );
  MUX2X1 U5649 ( .B(n3403), .A(n3404), .S(n4210), .Y(n3402) );
  MUX2X1 U5650 ( .B(n3406), .A(n3407), .S(n4210), .Y(n3405) );
  MUX2X1 U5651 ( .B(n3409), .A(n3410), .S(n4154), .Y(n3408) );
  MUX2X1 U5652 ( .B(n3412), .A(n3413), .S(n4211), .Y(n3411) );
  MUX2X1 U5653 ( .B(n3415), .A(n3416), .S(n4211), .Y(n3414) );
  MUX2X1 U5654 ( .B(n3418), .A(n3419), .S(n4211), .Y(n3417) );
  MUX2X1 U5655 ( .B(n3421), .A(n3422), .S(n4211), .Y(n3420) );
  MUX2X1 U5656 ( .B(n3424), .A(n3425), .S(n4154), .Y(n3423) );
  MUX2X1 U5657 ( .B(n3427), .A(n3428), .S(n4211), .Y(n3426) );
  MUX2X1 U5658 ( .B(n3430), .A(n3431), .S(n4211), .Y(n3429) );
  MUX2X1 U5659 ( .B(n3433), .A(n3434), .S(n4211), .Y(n3432) );
  MUX2X1 U5660 ( .B(n3436), .A(n3437), .S(n4211), .Y(n3435) );
  MUX2X1 U5661 ( .B(n3439), .A(n3440), .S(n4154), .Y(n3438) );
  MUX2X1 U5662 ( .B(n3442), .A(n3443), .S(n4211), .Y(n3441) );
  MUX2X1 U5663 ( .B(n3445), .A(n3446), .S(n4211), .Y(n3444) );
  MUX2X1 U5664 ( .B(n3448), .A(n3449), .S(n4211), .Y(n3447) );
  MUX2X1 U5665 ( .B(n3451), .A(n3452), .S(n4211), .Y(n3450) );
  MUX2X1 U5666 ( .B(n3454), .A(n3455), .S(n4154), .Y(n3453) );
  MUX2X1 U5667 ( .B(n3457), .A(n3458), .S(n4212), .Y(n3456) );
  MUX2X1 U5668 ( .B(n3460), .A(n3461), .S(n4212), .Y(n3459) );
  MUX2X1 U5669 ( .B(n3463), .A(n3464), .S(n4212), .Y(n3462) );
  MUX2X1 U5670 ( .B(n3466), .A(n3467), .S(n4212), .Y(n3465) );
  MUX2X1 U5671 ( .B(n3469), .A(n3470), .S(n4154), .Y(n3468) );
  MUX2X1 U5672 ( .B(n3472), .A(n3473), .S(n4212), .Y(n3471) );
  MUX2X1 U5673 ( .B(n3475), .A(n3476), .S(n4212), .Y(n3474) );
  MUX2X1 U5674 ( .B(n3478), .A(n3479), .S(n4212), .Y(n3477) );
  MUX2X1 U5675 ( .B(n3481), .A(n3482), .S(n4212), .Y(n3480) );
  MUX2X1 U5676 ( .B(n3484), .A(n3485), .S(n4154), .Y(n3483) );
  MUX2X1 U5677 ( .B(n3487), .A(n3488), .S(n4212), .Y(n3486) );
  MUX2X1 U5678 ( .B(n3490), .A(n3491), .S(n4212), .Y(n3489) );
  MUX2X1 U5679 ( .B(n3493), .A(n3494), .S(n4212), .Y(n3492) );
  MUX2X1 U5680 ( .B(n3496), .A(n3497), .S(n4212), .Y(n3495) );
  MUX2X1 U5681 ( .B(n3499), .A(n3500), .S(n4154), .Y(n3498) );
  MUX2X1 U5682 ( .B(n3502), .A(n3503), .S(n4213), .Y(n3501) );
  MUX2X1 U5683 ( .B(n3505), .A(n3506), .S(n4213), .Y(n3504) );
  MUX2X1 U5684 ( .B(n3508), .A(n3509), .S(n4213), .Y(n3507) );
  MUX2X1 U5685 ( .B(n3511), .A(n3512), .S(n4213), .Y(n3510) );
  MUX2X1 U5686 ( .B(n3514), .A(n3515), .S(n4154), .Y(n3513) );
  MUX2X1 U5687 ( .B(n3517), .A(n3518), .S(n4213), .Y(n3516) );
  MUX2X1 U5688 ( .B(n3520), .A(n3521), .S(n4213), .Y(n3519) );
  MUX2X1 U5689 ( .B(n3523), .A(n3524), .S(n4213), .Y(n3522) );
  MUX2X1 U5690 ( .B(n3526), .A(n3527), .S(n4213), .Y(n3525) );
  MUX2X1 U5691 ( .B(n3529), .A(n3530), .S(n4154), .Y(n3528) );
  MUX2X1 U5692 ( .B(n3532), .A(n3533), .S(n4213), .Y(n3531) );
  MUX2X1 U5693 ( .B(n3535), .A(n3536), .S(n4213), .Y(n3534) );
  MUX2X1 U5694 ( .B(n3538), .A(n3539), .S(n4213), .Y(n3537) );
  MUX2X1 U5695 ( .B(n3541), .A(n3542), .S(n4213), .Y(n3540) );
  MUX2X1 U5696 ( .B(n3544), .A(n3545), .S(n4154), .Y(n3543) );
  MUX2X1 U5697 ( .B(n3547), .A(n3548), .S(n4214), .Y(n3546) );
  MUX2X1 U5698 ( .B(n3550), .A(n3551), .S(n4214), .Y(n3549) );
  MUX2X1 U5699 ( .B(n3553), .A(n3554), .S(n4214), .Y(n3552) );
  MUX2X1 U5700 ( .B(n3556), .A(n3557), .S(n4214), .Y(n3555) );
  MUX2X1 U5701 ( .B(n3559), .A(n3560), .S(n4155), .Y(n3558) );
  MUX2X1 U5702 ( .B(n3562), .A(n3563), .S(n4214), .Y(n3561) );
  MUX2X1 U5703 ( .B(n3565), .A(n3566), .S(n4214), .Y(n3564) );
  MUX2X1 U5704 ( .B(n3568), .A(n3569), .S(n4214), .Y(n3567) );
  MUX2X1 U5705 ( .B(n3571), .A(n3572), .S(n4214), .Y(n3570) );
  MUX2X1 U5706 ( .B(n3574), .A(n3575), .S(n4155), .Y(n3573) );
  MUX2X1 U5707 ( .B(n3577), .A(n3578), .S(n4214), .Y(n3576) );
  MUX2X1 U5708 ( .B(n3580), .A(n3581), .S(n4214), .Y(n3579) );
  MUX2X1 U5709 ( .B(n3583), .A(n3584), .S(n4214), .Y(n3582) );
  MUX2X1 U5710 ( .B(n3586), .A(n3587), .S(n4214), .Y(n3585) );
  MUX2X1 U5711 ( .B(n3589), .A(n3590), .S(n4155), .Y(n3588) );
  MUX2X1 U5712 ( .B(n3592), .A(n3593), .S(n4215), .Y(n3591) );
  MUX2X1 U5713 ( .B(n3595), .A(n3596), .S(n4215), .Y(n3594) );
  MUX2X1 U5714 ( .B(n3598), .A(n3599), .S(n4215), .Y(n3597) );
  MUX2X1 U5715 ( .B(n3601), .A(n3602), .S(n4215), .Y(n3600) );
  MUX2X1 U5716 ( .B(n3604), .A(n3605), .S(n4155), .Y(n3603) );
  MUX2X1 U5717 ( .B(n3607), .A(n3608), .S(n4215), .Y(n3606) );
  MUX2X1 U5718 ( .B(n3610), .A(n3611), .S(n4215), .Y(n3609) );
  MUX2X1 U5719 ( .B(n3613), .A(n3614), .S(n4215), .Y(n3612) );
  MUX2X1 U5720 ( .B(n3616), .A(n3617), .S(n4215), .Y(n3615) );
  MUX2X1 U5721 ( .B(n3619), .A(n3620), .S(n4155), .Y(n3618) );
  MUX2X1 U5722 ( .B(n3622), .A(n3623), .S(n4215), .Y(n3621) );
  MUX2X1 U5723 ( .B(n3625), .A(n3626), .S(n4215), .Y(n3624) );
  MUX2X1 U5724 ( .B(n3628), .A(n3629), .S(n4215), .Y(n3627) );
  MUX2X1 U5725 ( .B(n3631), .A(n3632), .S(n4215), .Y(n3630) );
  MUX2X1 U5726 ( .B(n3634), .A(n3635), .S(n4155), .Y(n3633) );
  MUX2X1 U5727 ( .B(n3637), .A(n3638), .S(n4216), .Y(n3636) );
  MUX2X1 U5728 ( .B(n3640), .A(n3641), .S(n4216), .Y(n3639) );
  MUX2X1 U5729 ( .B(n3643), .A(n3644), .S(n4216), .Y(n3642) );
  MUX2X1 U5730 ( .B(n3646), .A(n3647), .S(n4216), .Y(n3645) );
  MUX2X1 U5731 ( .B(n3649), .A(n3650), .S(n4155), .Y(n3648) );
  MUX2X1 U5732 ( .B(n3652), .A(n3653), .S(n4216), .Y(n3651) );
  MUX2X1 U5733 ( .B(n3655), .A(n3656), .S(n4216), .Y(n3654) );
  MUX2X1 U5734 ( .B(n3658), .A(n3659), .S(n4216), .Y(n3657) );
  MUX2X1 U5735 ( .B(n3661), .A(n3662), .S(n4216), .Y(n3660) );
  MUX2X1 U5736 ( .B(n3664), .A(n3665), .S(n4155), .Y(n3663) );
  MUX2X1 U5737 ( .B(n3667), .A(n3668), .S(n4216), .Y(n3666) );
  MUX2X1 U5738 ( .B(n3670), .A(n3671), .S(n4216), .Y(n3669) );
  MUX2X1 U5739 ( .B(n3673), .A(n3674), .S(n4216), .Y(n3672) );
  MUX2X1 U5740 ( .B(n3676), .A(n3677), .S(n4216), .Y(n3675) );
  MUX2X1 U5741 ( .B(n3679), .A(n3680), .S(n4155), .Y(n3678) );
  MUX2X1 U5742 ( .B(n3682), .A(n3683), .S(n4217), .Y(n3681) );
  MUX2X1 U5743 ( .B(n3685), .A(n3686), .S(n4217), .Y(n3684) );
  MUX2X1 U5744 ( .B(n3688), .A(n3689), .S(n4217), .Y(n3687) );
  MUX2X1 U5745 ( .B(n3691), .A(n3692), .S(n4217), .Y(n3690) );
  MUX2X1 U5746 ( .B(n3694), .A(n3695), .S(n4155), .Y(n3693) );
  MUX2X1 U5747 ( .B(n3697), .A(n3698), .S(n4217), .Y(n3696) );
  MUX2X1 U5748 ( .B(n3700), .A(n3701), .S(n4217), .Y(n3699) );
  MUX2X1 U5749 ( .B(n3703), .A(n3704), .S(n4217), .Y(n3702) );
  MUX2X1 U5750 ( .B(n3706), .A(n3707), .S(n4217), .Y(n3705) );
  MUX2X1 U5751 ( .B(n3709), .A(n3710), .S(n4155), .Y(n3708) );
  MUX2X1 U5752 ( .B(n3712), .A(n3713), .S(n4217), .Y(n3711) );
  MUX2X1 U5753 ( .B(n3715), .A(n3716), .S(n4217), .Y(n3714) );
  MUX2X1 U5754 ( .B(n3718), .A(n3719), .S(n4217), .Y(n3717) );
  MUX2X1 U5755 ( .B(n3721), .A(n3722), .S(n4217), .Y(n3720) );
  MUX2X1 U5756 ( .B(n3724), .A(n3725), .S(n4155), .Y(n3723) );
  MUX2X1 U5757 ( .B(n3727), .A(n3728), .S(n4218), .Y(n3726) );
  MUX2X1 U5758 ( .B(n3730), .A(n3731), .S(n4218), .Y(n3729) );
  MUX2X1 U5759 ( .B(n3733), .A(n3734), .S(n4218), .Y(n3732) );
  MUX2X1 U5760 ( .B(n3736), .A(n3737), .S(n4218), .Y(n3735) );
  MUX2X1 U5761 ( .B(n3739), .A(n3740), .S(n4156), .Y(n3738) );
  MUX2X1 U5762 ( .B(n3742), .A(n3743), .S(n4218), .Y(n3741) );
  MUX2X1 U5763 ( .B(n3745), .A(n3746), .S(n4218), .Y(n3744) );
  MUX2X1 U5764 ( .B(n3748), .A(n3749), .S(n4218), .Y(n3747) );
  MUX2X1 U5765 ( .B(n3751), .A(n3752), .S(n4218), .Y(n3750) );
  MUX2X1 U5766 ( .B(n3754), .A(n3755), .S(n4156), .Y(n3753) );
  MUX2X1 U5767 ( .B(n3757), .A(n3758), .S(n4218), .Y(n3756) );
  MUX2X1 U5768 ( .B(n3760), .A(n3761), .S(n4218), .Y(n3759) );
  MUX2X1 U5769 ( .B(n3763), .A(n3764), .S(n4218), .Y(n3762) );
  MUX2X1 U5770 ( .B(n3766), .A(n3767), .S(n4218), .Y(n3765) );
  MUX2X1 U5771 ( .B(n3769), .A(n3770), .S(n4156), .Y(n3768) );
  MUX2X1 U5772 ( .B(n3772), .A(n3773), .S(n4208), .Y(n3771) );
  MUX2X1 U5773 ( .B(n3775), .A(n3776), .S(n4198), .Y(n3774) );
  MUX2X1 U5774 ( .B(n3778), .A(n3779), .S(n4206), .Y(n3777) );
  MUX2X1 U5775 ( .B(n3781), .A(n3782), .S(n4197), .Y(n3780) );
  MUX2X1 U5776 ( .B(n3784), .A(n3785), .S(n4156), .Y(n3783) );
  MUX2X1 U5777 ( .B(n3787), .A(n3788), .S(n4188), .Y(n3786) );
  MUX2X1 U5778 ( .B(n3790), .A(n3791), .S(n4198), .Y(n3789) );
  MUX2X1 U5779 ( .B(n3793), .A(n3794), .S(n4220), .Y(n3792) );
  MUX2X1 U5780 ( .B(n3796), .A(n3797), .S(n4196), .Y(n3795) );
  MUX2X1 U5781 ( .B(n3799), .A(n3800), .S(n4156), .Y(n3798) );
  MUX2X1 U5782 ( .B(n3802), .A(n3803), .S(n4219), .Y(n3801) );
  MUX2X1 U5783 ( .B(n3805), .A(n3806), .S(n4196), .Y(n3804) );
  MUX2X1 U5784 ( .B(n3808), .A(n3809), .S(n4217), .Y(n3807) );
  MUX2X1 U5785 ( .B(n3811), .A(n3812), .S(n4209), .Y(n3810) );
  MUX2X1 U5786 ( .B(n3814), .A(n3815), .S(n4156), .Y(n3813) );
  MUX2X1 U5787 ( .B(n3817), .A(n3818), .S(n4219), .Y(n3816) );
  MUX2X1 U5788 ( .B(n3820), .A(n3821), .S(n4219), .Y(n3819) );
  MUX2X1 U5789 ( .B(n3823), .A(n3824), .S(n4219), .Y(n3822) );
  MUX2X1 U5790 ( .B(n3826), .A(n3827), .S(n4219), .Y(n3825) );
  MUX2X1 U5791 ( .B(n3829), .A(n3830), .S(n4156), .Y(n3828) );
  MUX2X1 U5792 ( .B(n3832), .A(n3833), .S(n4219), .Y(n3831) );
  MUX2X1 U5793 ( .B(n3835), .A(n3836), .S(n4219), .Y(n3834) );
  MUX2X1 U5794 ( .B(n3838), .A(n3839), .S(n4219), .Y(n3837) );
  MUX2X1 U5795 ( .B(n3841), .A(n3842), .S(n4219), .Y(n3840) );
  MUX2X1 U5796 ( .B(n3844), .A(n3845), .S(n4156), .Y(n3843) );
  MUX2X1 U5797 ( .B(n3847), .A(n3848), .S(n4219), .Y(n3846) );
  MUX2X1 U5798 ( .B(n3850), .A(n3851), .S(n4219), .Y(n3849) );
  MUX2X1 U5799 ( .B(n3853), .A(n3854), .S(n4219), .Y(n3852) );
  MUX2X1 U5800 ( .B(n3856), .A(n3857), .S(n4219), .Y(n3855) );
  MUX2X1 U5801 ( .B(n3859), .A(n3860), .S(n4156), .Y(n3858) );
  MUX2X1 U5802 ( .B(n3862), .A(n3863), .S(n4220), .Y(n3861) );
  MUX2X1 U5803 ( .B(n3865), .A(n3866), .S(n4220), .Y(n3864) );
  MUX2X1 U5804 ( .B(n3868), .A(n3869), .S(n4220), .Y(n3867) );
  MUX2X1 U5805 ( .B(n3871), .A(n3872), .S(n4220), .Y(n3870) );
  MUX2X1 U5806 ( .B(n3874), .A(n3875), .S(n4156), .Y(n3873) );
  MUX2X1 U5807 ( .B(n3877), .A(n3878), .S(n4220), .Y(n3876) );
  MUX2X1 U5808 ( .B(n3880), .A(n3881), .S(n4220), .Y(n3879) );
  MUX2X1 U5809 ( .B(n3883), .A(n3884), .S(n4220), .Y(n3882) );
  MUX2X1 U5810 ( .B(n3886), .A(n3887), .S(n4220), .Y(n3885) );
  MUX2X1 U5811 ( .B(n3889), .A(n3890), .S(n4156), .Y(n3888) );
  MUX2X1 U5812 ( .B(n3892), .A(n3893), .S(n4220), .Y(n3891) );
  MUX2X1 U5813 ( .B(n3895), .A(n3896), .S(n4220), .Y(n3894) );
  MUX2X1 U5814 ( .B(n3898), .A(n3899), .S(n4220), .Y(n3897) );
  MUX2X1 U5815 ( .B(n3901), .A(n3902), .S(n4220), .Y(n3900) );
  MUX2X1 U5816 ( .B(n3904), .A(n3905), .S(n4156), .Y(n3903) );
  MUX2X1 U5817 ( .B(n3907), .A(n3908), .S(n4221), .Y(n3906) );
  MUX2X1 U5818 ( .B(n3910), .A(n3911), .S(n4221), .Y(n3909) );
  MUX2X1 U5819 ( .B(n3913), .A(n3914), .S(n4221), .Y(n3912) );
  MUX2X1 U5820 ( .B(n3916), .A(n3917), .S(n4221), .Y(n3915) );
  MUX2X1 U5821 ( .B(n3919), .A(n3920), .S(n4157), .Y(n3918) );
  MUX2X1 U5822 ( .B(n3922), .A(n3923), .S(n4221), .Y(n3921) );
  MUX2X1 U5823 ( .B(n3925), .A(n3926), .S(n4221), .Y(n3924) );
  MUX2X1 U5824 ( .B(n3928), .A(n3929), .S(n4221), .Y(n3927) );
  MUX2X1 U5825 ( .B(n3931), .A(n3932), .S(n4221), .Y(n3930) );
  MUX2X1 U5826 ( .B(n3934), .A(n3935), .S(n4157), .Y(n3933) );
  MUX2X1 U5827 ( .B(n3937), .A(n3938), .S(n4221), .Y(n3936) );
  MUX2X1 U5828 ( .B(n3940), .A(n3941), .S(n4221), .Y(n3939) );
  MUX2X1 U5829 ( .B(n3943), .A(n3944), .S(n4221), .Y(n3942) );
  MUX2X1 U5830 ( .B(n3946), .A(n3947), .S(n4221), .Y(n3945) );
  MUX2X1 U5831 ( .B(n3949), .A(n3950), .S(n4157), .Y(n3948) );
  MUX2X1 U5832 ( .B(n3952), .A(n3953), .S(n4222), .Y(n3951) );
  MUX2X1 U5833 ( .B(n3955), .A(n3956), .S(n4222), .Y(n3954) );
  MUX2X1 U5834 ( .B(n3958), .A(n3959), .S(n4222), .Y(n3957) );
  MUX2X1 U5835 ( .B(n3961), .A(n3962), .S(n4222), .Y(n3960) );
  MUX2X1 U5836 ( .B(n3964), .A(n3965), .S(n4157), .Y(n3963) );
  MUX2X1 U5837 ( .B(n3967), .A(n3968), .S(n4222), .Y(n3966) );
  MUX2X1 U5838 ( .B(n3970), .A(n3971), .S(n4222), .Y(n3969) );
  MUX2X1 U5839 ( .B(n3973), .A(n3974), .S(n4222), .Y(n3972) );
  MUX2X1 U5840 ( .B(n3976), .A(n3977), .S(n4222), .Y(n3975) );
  MUX2X1 U5841 ( .B(n3979), .A(n3980), .S(n4157), .Y(n3978) );
  MUX2X1 U5842 ( .B(n3982), .A(n3983), .S(n4222), .Y(n3981) );
  MUX2X1 U5843 ( .B(n3985), .A(n3986), .S(n4222), .Y(n3984) );
  MUX2X1 U5844 ( .B(n3988), .A(n3989), .S(n4222), .Y(n3987) );
  MUX2X1 U5845 ( .B(n3991), .A(n3992), .S(n4222), .Y(n3990) );
  MUX2X1 U5846 ( .B(n3994), .A(n3995), .S(n4157), .Y(n3993) );
  MUX2X1 U5847 ( .B(n3997), .A(n3998), .S(n4220), .Y(n3996) );
  MUX2X1 U5848 ( .B(n4000), .A(n4001), .S(n4192), .Y(n3999) );
  MUX2X1 U5849 ( .B(n4003), .A(n4004), .S(n4193), .Y(n4002) );
  MUX2X1 U5850 ( .B(n4006), .A(n4007), .S(n4197), .Y(n4005) );
  MUX2X1 U5851 ( .B(n4009), .A(n4010), .S(n4157), .Y(n4008) );
  MUX2X1 U5852 ( .B(n4012), .A(n4013), .S(n4191), .Y(n4011) );
  MUX2X1 U5853 ( .B(n4015), .A(n4016), .S(n4222), .Y(n4014) );
  MUX2X1 U5854 ( .B(n4018), .A(n4019), .S(n4222), .Y(n4017) );
  MUX2X1 U5855 ( .B(n4021), .A(n4022), .S(n4220), .Y(n4020) );
  MUX2X1 U5856 ( .B(n4024), .A(n4025), .S(n4157), .Y(n4023) );
  MUX2X1 U5857 ( .B(n4027), .A(n4028), .S(n4214), .Y(n4026) );
  MUX2X1 U5858 ( .B(n4030), .A(n4031), .S(n4221), .Y(n4029) );
  MUX2X1 U5859 ( .B(n4033), .A(n4034), .S(n4198), .Y(n4032) );
  MUX2X1 U5860 ( .B(n4036), .A(n4037), .S(n4218), .Y(n4035) );
  MUX2X1 U5861 ( .B(n4039), .A(n4040), .S(n4157), .Y(n4038) );
  MUX2X1 U5862 ( .B(n4042), .A(n4043), .S(n4214), .Y(n4041) );
  MUX2X1 U5863 ( .B(n4045), .A(n4046), .S(n4221), .Y(n4044) );
  MUX2X1 U5864 ( .B(n4048), .A(n4049), .S(n4221), .Y(n4047) );
  MUX2X1 U5865 ( .B(n4051), .A(n4052), .S(n4221), .Y(n4050) );
  MUX2X1 U5866 ( .B(n4054), .A(n4055), .S(n4157), .Y(n4053) );
  MUX2X1 U5867 ( .B(n4057), .A(n4058), .S(n4221), .Y(n4056) );
  MUX2X1 U5868 ( .B(n4060), .A(n4061), .S(n4190), .Y(n4059) );
  MUX2X1 U5869 ( .B(n4063), .A(n4064), .S(n4190), .Y(n4062) );
  MUX2X1 U5870 ( .B(n4066), .A(n4067), .S(n4193), .Y(n4065) );
  MUX2X1 U5871 ( .B(n4069), .A(n4070), .S(n4157), .Y(n4068) );
  MUX2X1 U5872 ( .B(n4072), .A(n4073), .S(n4221), .Y(n4071) );
  MUX2X1 U5873 ( .B(n4075), .A(n4076), .S(n4214), .Y(n4074) );
  MUX2X1 U5874 ( .B(n4078), .A(n4079), .S(n4214), .Y(n4077) );
  MUX2X1 U5875 ( .B(n4081), .A(n4082), .S(n4193), .Y(n4080) );
  MUX2X1 U5876 ( .B(n4084), .A(n4085), .S(n4157), .Y(n4083) );
  MUX2X1 U5877 ( .B(ram[64]), .A(ram[0]), .S(n4248), .Y(n2160) );
  MUX2X1 U5878 ( .B(ram[192]), .A(ram[128]), .S(n4248), .Y(n2159) );
  MUX2X1 U5879 ( .B(ram[320]), .A(ram[256]), .S(n4248), .Y(n2163) );
  MUX2X1 U5880 ( .B(ram[448]), .A(ram[384]), .S(n4248), .Y(n2162) );
  MUX2X1 U5881 ( .B(n2161), .A(n2158), .S(n4162), .Y(n2172) );
  MUX2X1 U5882 ( .B(ram[576]), .A(ram[512]), .S(n4249), .Y(n2166) );
  MUX2X1 U5883 ( .B(ram[704]), .A(ram[640]), .S(n4249), .Y(n2165) );
  MUX2X1 U5884 ( .B(ram[832]), .A(ram[768]), .S(n4249), .Y(n2169) );
  MUX2X1 U5885 ( .B(ram[960]), .A(ram[896]), .S(n4249), .Y(n2168) );
  MUX2X1 U5886 ( .B(n2167), .A(n2164), .S(n4163), .Y(n2171) );
  MUX2X1 U5887 ( .B(ram[1088]), .A(ram[1024]), .S(n4249), .Y(n2175) );
  MUX2X1 U5888 ( .B(ram[1216]), .A(ram[1152]), .S(n4249), .Y(n2174) );
  MUX2X1 U5889 ( .B(ram[1344]), .A(ram[1280]), .S(n4249), .Y(n2178) );
  MUX2X1 U5890 ( .B(ram[1472]), .A(ram[1408]), .S(n4249), .Y(n2177) );
  MUX2X1 U5891 ( .B(n2176), .A(n2173), .S(n4165), .Y(n2187) );
  MUX2X1 U5892 ( .B(ram[1600]), .A(ram[1536]), .S(n4249), .Y(n2181) );
  MUX2X1 U5893 ( .B(ram[1728]), .A(ram[1664]), .S(n4249), .Y(n2180) );
  MUX2X1 U5894 ( .B(ram[1856]), .A(ram[1792]), .S(n4249), .Y(n2184) );
  MUX2X1 U5895 ( .B(ram[1984]), .A(ram[1920]), .S(n4249), .Y(n2183) );
  MUX2X1 U5896 ( .B(n2182), .A(n2179), .S(n4160), .Y(n2186) );
  MUX2X1 U5897 ( .B(n2185), .A(n2170), .S(n4151), .Y(n4086) );
  MUX2X1 U5898 ( .B(ram[65]), .A(ram[1]), .S(n4250), .Y(n2190) );
  MUX2X1 U5899 ( .B(ram[193]), .A(ram[129]), .S(n4250), .Y(n2189) );
  MUX2X1 U5900 ( .B(ram[321]), .A(ram[257]), .S(n4250), .Y(n2193) );
  MUX2X1 U5901 ( .B(ram[449]), .A(ram[385]), .S(n4250), .Y(n2192) );
  MUX2X1 U5902 ( .B(n2191), .A(n2188), .S(n4158), .Y(n2202) );
  MUX2X1 U5903 ( .B(ram[577]), .A(ram[513]), .S(n4250), .Y(n2196) );
  MUX2X1 U5904 ( .B(ram[705]), .A(ram[641]), .S(n4250), .Y(n2195) );
  MUX2X1 U5905 ( .B(ram[833]), .A(ram[769]), .S(n4250), .Y(n2199) );
  MUX2X1 U5906 ( .B(ram[961]), .A(ram[897]), .S(n4250), .Y(n2198) );
  MUX2X1 U5907 ( .B(n2197), .A(n2194), .S(n4158), .Y(n2201) );
  MUX2X1 U5908 ( .B(ram[1089]), .A(ram[1025]), .S(n4250), .Y(n2205) );
  MUX2X1 U5909 ( .B(ram[1217]), .A(ram[1153]), .S(n4250), .Y(n2204) );
  MUX2X1 U5910 ( .B(ram[1345]), .A(ram[1281]), .S(n4250), .Y(n2208) );
  MUX2X1 U5911 ( .B(ram[1473]), .A(ram[1409]), .S(n4250), .Y(n2207) );
  MUX2X1 U5912 ( .B(n2206), .A(n2203), .S(n4158), .Y(n2217) );
  MUX2X1 U5913 ( .B(ram[1601]), .A(ram[1537]), .S(n4251), .Y(n2211) );
  MUX2X1 U5914 ( .B(ram[1729]), .A(ram[1665]), .S(n4251), .Y(n2210) );
  MUX2X1 U5915 ( .B(ram[1857]), .A(ram[1793]), .S(n4251), .Y(n2214) );
  MUX2X1 U5916 ( .B(ram[1985]), .A(ram[1921]), .S(n4251), .Y(n2213) );
  MUX2X1 U5917 ( .B(n2212), .A(n2209), .S(n4158), .Y(n2216) );
  MUX2X1 U5918 ( .B(n2215), .A(n2200), .S(n4152), .Y(n4087) );
  MUX2X1 U5919 ( .B(ram[66]), .A(ram[2]), .S(n4251), .Y(n2220) );
  MUX2X1 U5920 ( .B(ram[194]), .A(ram[130]), .S(n4251), .Y(n2219) );
  MUX2X1 U5921 ( .B(ram[322]), .A(ram[258]), .S(n4251), .Y(n2223) );
  MUX2X1 U5922 ( .B(ram[450]), .A(ram[386]), .S(n4251), .Y(n2222) );
  MUX2X1 U5923 ( .B(n2221), .A(n2218), .S(n4158), .Y(n2232) );
  MUX2X1 U5924 ( .B(ram[578]), .A(ram[514]), .S(n4251), .Y(n2226) );
  MUX2X1 U5925 ( .B(ram[706]), .A(ram[642]), .S(n4251), .Y(n2225) );
  MUX2X1 U5926 ( .B(ram[834]), .A(ram[770]), .S(n4251), .Y(n2229) );
  MUX2X1 U5927 ( .B(ram[962]), .A(ram[898]), .S(n4251), .Y(n2228) );
  MUX2X1 U5928 ( .B(n2227), .A(n2224), .S(n4158), .Y(n2231) );
  MUX2X1 U5929 ( .B(ram[1090]), .A(ram[1026]), .S(n4252), .Y(n2235) );
  MUX2X1 U5930 ( .B(ram[1218]), .A(ram[1154]), .S(n4252), .Y(n2234) );
  MUX2X1 U5931 ( .B(ram[1346]), .A(ram[1282]), .S(n4252), .Y(n2238) );
  MUX2X1 U5932 ( .B(ram[1474]), .A(ram[1410]), .S(n4252), .Y(n2237) );
  MUX2X1 U5933 ( .B(n2236), .A(n2233), .S(n4158), .Y(n2247) );
  MUX2X1 U5934 ( .B(ram[1602]), .A(ram[1538]), .S(n4252), .Y(n2241) );
  MUX2X1 U5935 ( .B(ram[1730]), .A(ram[1666]), .S(n4252), .Y(n2240) );
  MUX2X1 U5936 ( .B(ram[1858]), .A(ram[1794]), .S(n4252), .Y(n2244) );
  MUX2X1 U5937 ( .B(ram[1986]), .A(ram[1922]), .S(n4252), .Y(n2243) );
  MUX2X1 U5938 ( .B(n2242), .A(n2239), .S(n4158), .Y(n2246) );
  MUX2X1 U5939 ( .B(n2245), .A(n2230), .S(n4152), .Y(n4088) );
  MUX2X1 U5940 ( .B(ram[67]), .A(ram[3]), .S(n4252), .Y(n2250) );
  MUX2X1 U5941 ( .B(ram[195]), .A(ram[131]), .S(n4252), .Y(n2249) );
  MUX2X1 U5942 ( .B(ram[323]), .A(ram[259]), .S(n4252), .Y(n2253) );
  MUX2X1 U5943 ( .B(ram[451]), .A(ram[387]), .S(n4252), .Y(n2252) );
  MUX2X1 U5944 ( .B(n2251), .A(n2248), .S(n4158), .Y(n2262) );
  MUX2X1 U5945 ( .B(ram[579]), .A(ram[515]), .S(n4253), .Y(n2256) );
  MUX2X1 U5946 ( .B(ram[707]), .A(ram[643]), .S(n4253), .Y(n2255) );
  MUX2X1 U5947 ( .B(ram[835]), .A(ram[771]), .S(n4253), .Y(n2259) );
  MUX2X1 U5948 ( .B(ram[963]), .A(ram[899]), .S(n4253), .Y(n2258) );
  MUX2X1 U5949 ( .B(n2257), .A(n2254), .S(n4158), .Y(n2261) );
  MUX2X1 U5950 ( .B(ram[1091]), .A(ram[1027]), .S(n4253), .Y(n2265) );
  MUX2X1 U5951 ( .B(ram[1219]), .A(ram[1155]), .S(n4253), .Y(n2264) );
  MUX2X1 U5952 ( .B(ram[1347]), .A(ram[1283]), .S(n4253), .Y(n2268) );
  MUX2X1 U5953 ( .B(ram[1475]), .A(ram[1411]), .S(n4253), .Y(n2267) );
  MUX2X1 U5954 ( .B(n2266), .A(n2263), .S(n4158), .Y(n2277) );
  MUX2X1 U5955 ( .B(ram[1603]), .A(ram[1539]), .S(n4253), .Y(n2271) );
  MUX2X1 U5956 ( .B(ram[1731]), .A(ram[1667]), .S(n4253), .Y(n2270) );
  MUX2X1 U5957 ( .B(ram[1859]), .A(ram[1795]), .S(n4253), .Y(n2274) );
  MUX2X1 U5958 ( .B(ram[1987]), .A(ram[1923]), .S(n4253), .Y(n2273) );
  MUX2X1 U5959 ( .B(n2272), .A(n2269), .S(n4158), .Y(n2276) );
  MUX2X1 U5960 ( .B(n2275), .A(n2260), .S(n4152), .Y(n4089) );
  MUX2X1 U5961 ( .B(ram[68]), .A(ram[4]), .S(n4254), .Y(n2280) );
  MUX2X1 U5962 ( .B(ram[196]), .A(ram[132]), .S(n4254), .Y(n2279) );
  MUX2X1 U5963 ( .B(ram[324]), .A(ram[260]), .S(n4254), .Y(n2283) );
  MUX2X1 U5964 ( .B(ram[452]), .A(ram[388]), .S(n4254), .Y(n2282) );
  MUX2X1 U5965 ( .B(n2281), .A(n2278), .S(n4159), .Y(n2292) );
  MUX2X1 U5966 ( .B(ram[580]), .A(ram[516]), .S(n4254), .Y(n2286) );
  MUX2X1 U5967 ( .B(ram[708]), .A(ram[644]), .S(n4254), .Y(n2285) );
  MUX2X1 U5968 ( .B(ram[836]), .A(ram[772]), .S(n4254), .Y(n2289) );
  MUX2X1 U5969 ( .B(ram[964]), .A(ram[900]), .S(n4254), .Y(n2288) );
  MUX2X1 U5970 ( .B(n2287), .A(n2284), .S(n4159), .Y(n2291) );
  MUX2X1 U5971 ( .B(ram[1092]), .A(ram[1028]), .S(n4254), .Y(n2295) );
  MUX2X1 U5972 ( .B(ram[1220]), .A(ram[1156]), .S(n4254), .Y(n2294) );
  MUX2X1 U5973 ( .B(ram[1348]), .A(ram[1284]), .S(n4254), .Y(n2298) );
  MUX2X1 U5974 ( .B(ram[1476]), .A(ram[1412]), .S(n4254), .Y(n2297) );
  MUX2X1 U5975 ( .B(n2296), .A(n2293), .S(n4159), .Y(n2307) );
  MUX2X1 U5976 ( .B(ram[1604]), .A(ram[1540]), .S(n4255), .Y(n2301) );
  MUX2X1 U5977 ( .B(ram[1732]), .A(ram[1668]), .S(n4255), .Y(n2300) );
  MUX2X1 U5978 ( .B(ram[1860]), .A(ram[1796]), .S(n4255), .Y(n2304) );
  MUX2X1 U5979 ( .B(ram[1988]), .A(ram[1924]), .S(n4255), .Y(n2303) );
  MUX2X1 U5980 ( .B(n2302), .A(n2299), .S(n4159), .Y(n2306) );
  MUX2X1 U5981 ( .B(n2305), .A(n2290), .S(n4152), .Y(n4090) );
  MUX2X1 U5982 ( .B(ram[69]), .A(ram[5]), .S(n4255), .Y(n2310) );
  MUX2X1 U5983 ( .B(ram[197]), .A(ram[133]), .S(n4255), .Y(n2309) );
  MUX2X1 U5984 ( .B(ram[325]), .A(ram[261]), .S(n4255), .Y(n2313) );
  MUX2X1 U5985 ( .B(ram[453]), .A(ram[389]), .S(n4255), .Y(n2312) );
  MUX2X1 U5986 ( .B(n2311), .A(n2308), .S(n4159), .Y(n2322) );
  MUX2X1 U5987 ( .B(ram[581]), .A(ram[517]), .S(n4255), .Y(n2316) );
  MUX2X1 U5988 ( .B(ram[709]), .A(ram[645]), .S(n4255), .Y(n2315) );
  MUX2X1 U5989 ( .B(ram[837]), .A(ram[773]), .S(n4255), .Y(n2319) );
  MUX2X1 U5990 ( .B(ram[965]), .A(ram[901]), .S(n4255), .Y(n2318) );
  MUX2X1 U5991 ( .B(n2317), .A(n2314), .S(n4159), .Y(n2321) );
  MUX2X1 U5992 ( .B(ram[1093]), .A(ram[1029]), .S(n4256), .Y(n2325) );
  MUX2X1 U5993 ( .B(ram[1221]), .A(ram[1157]), .S(n4256), .Y(n2324) );
  MUX2X1 U5994 ( .B(ram[1349]), .A(ram[1285]), .S(n4256), .Y(n2328) );
  MUX2X1 U5995 ( .B(ram[1477]), .A(ram[1413]), .S(n4256), .Y(n2327) );
  MUX2X1 U5996 ( .B(n2326), .A(n2323), .S(n4159), .Y(n2337) );
  MUX2X1 U5997 ( .B(ram[1605]), .A(ram[1541]), .S(n4256), .Y(n2331) );
  MUX2X1 U5998 ( .B(ram[1733]), .A(ram[1669]), .S(n4256), .Y(n2330) );
  MUX2X1 U5999 ( .B(ram[1861]), .A(ram[1797]), .S(n4256), .Y(n2334) );
  MUX2X1 U6000 ( .B(ram[1989]), .A(ram[1925]), .S(n4256), .Y(n2333) );
  MUX2X1 U6001 ( .B(n2332), .A(n2329), .S(n4159), .Y(n2336) );
  MUX2X1 U6002 ( .B(n2335), .A(n2320), .S(n4151), .Y(n4091) );
  MUX2X1 U6003 ( .B(ram[70]), .A(ram[6]), .S(n4256), .Y(n2340) );
  MUX2X1 U6004 ( .B(ram[198]), .A(ram[134]), .S(n4256), .Y(n2339) );
  MUX2X1 U6005 ( .B(ram[326]), .A(ram[262]), .S(n4256), .Y(n2343) );
  MUX2X1 U6006 ( .B(ram[454]), .A(ram[390]), .S(n4256), .Y(n2342) );
  MUX2X1 U6007 ( .B(n2341), .A(n2338), .S(n4159), .Y(n2352) );
  MUX2X1 U6008 ( .B(ram[582]), .A(ram[518]), .S(n4257), .Y(n2346) );
  MUX2X1 U6009 ( .B(ram[710]), .A(ram[646]), .S(n4257), .Y(n2345) );
  MUX2X1 U6010 ( .B(ram[838]), .A(ram[774]), .S(n4257), .Y(n2349) );
  MUX2X1 U6011 ( .B(ram[966]), .A(ram[902]), .S(n4257), .Y(n2348) );
  MUX2X1 U6012 ( .B(n2347), .A(n2344), .S(n4159), .Y(n2351) );
  MUX2X1 U6013 ( .B(ram[1094]), .A(ram[1030]), .S(n4257), .Y(n2355) );
  MUX2X1 U6014 ( .B(ram[1222]), .A(ram[1158]), .S(n4257), .Y(n2354) );
  MUX2X1 U6015 ( .B(ram[1350]), .A(ram[1286]), .S(n4257), .Y(n2358) );
  MUX2X1 U6016 ( .B(ram[1478]), .A(ram[1414]), .S(n4257), .Y(n2357) );
  MUX2X1 U6017 ( .B(n2356), .A(n2353), .S(n4159), .Y(n2367) );
  MUX2X1 U6018 ( .B(ram[1606]), .A(ram[1542]), .S(n4257), .Y(n2361) );
  MUX2X1 U6019 ( .B(ram[1734]), .A(ram[1670]), .S(n4257), .Y(n2360) );
  MUX2X1 U6020 ( .B(ram[1862]), .A(ram[1798]), .S(n4257), .Y(n2364) );
  MUX2X1 U6021 ( .B(ram[1990]), .A(ram[1926]), .S(n4257), .Y(n2363) );
  MUX2X1 U6022 ( .B(n2362), .A(n2359), .S(n4159), .Y(n2366) );
  MUX2X1 U6023 ( .B(n2365), .A(n2350), .S(n4151), .Y(n4092) );
  MUX2X1 U6024 ( .B(ram[71]), .A(ram[7]), .S(n4258), .Y(n2370) );
  MUX2X1 U6025 ( .B(ram[199]), .A(ram[135]), .S(n4258), .Y(n2369) );
  MUX2X1 U6026 ( .B(ram[327]), .A(ram[263]), .S(n4258), .Y(n2373) );
  MUX2X1 U6027 ( .B(ram[455]), .A(ram[391]), .S(n4258), .Y(n2372) );
  MUX2X1 U6028 ( .B(n2371), .A(n2368), .S(n4160), .Y(n2382) );
  MUX2X1 U6029 ( .B(ram[583]), .A(ram[519]), .S(n4258), .Y(n2376) );
  MUX2X1 U6030 ( .B(ram[711]), .A(ram[647]), .S(n4258), .Y(n2375) );
  MUX2X1 U6031 ( .B(ram[839]), .A(ram[775]), .S(n4258), .Y(n2379) );
  MUX2X1 U6032 ( .B(ram[967]), .A(ram[903]), .S(n4258), .Y(n2378) );
  MUX2X1 U6033 ( .B(n2377), .A(n2374), .S(n4160), .Y(n2381) );
  MUX2X1 U6034 ( .B(ram[1095]), .A(ram[1031]), .S(n4258), .Y(n2385) );
  MUX2X1 U6035 ( .B(ram[1223]), .A(ram[1159]), .S(n4258), .Y(n2384) );
  MUX2X1 U6036 ( .B(ram[1351]), .A(ram[1287]), .S(n4258), .Y(n2388) );
  MUX2X1 U6037 ( .B(ram[1479]), .A(ram[1415]), .S(n4258), .Y(n2387) );
  MUX2X1 U6038 ( .B(n2386), .A(n2383), .S(n4160), .Y(n2397) );
  MUX2X1 U6039 ( .B(ram[1607]), .A(ram[1543]), .S(n4259), .Y(n2391) );
  MUX2X1 U6040 ( .B(ram[1735]), .A(ram[1671]), .S(n4259), .Y(n2390) );
  MUX2X1 U6041 ( .B(ram[1863]), .A(ram[1799]), .S(n4259), .Y(n2394) );
  MUX2X1 U6042 ( .B(ram[1991]), .A(ram[1927]), .S(n4259), .Y(n2393) );
  MUX2X1 U6043 ( .B(n2392), .A(n2389), .S(n4160), .Y(n2396) );
  MUX2X1 U6044 ( .B(n2395), .A(n2380), .S(n4152), .Y(n4093) );
  MUX2X1 U6045 ( .B(ram[72]), .A(ram[8]), .S(n4259), .Y(n2400) );
  MUX2X1 U6046 ( .B(ram[200]), .A(ram[136]), .S(n4259), .Y(n2399) );
  MUX2X1 U6047 ( .B(ram[328]), .A(ram[264]), .S(n4259), .Y(n2403) );
  MUX2X1 U6048 ( .B(ram[456]), .A(ram[392]), .S(n4259), .Y(n2402) );
  MUX2X1 U6049 ( .B(n2401), .A(n2398), .S(n4160), .Y(n2412) );
  MUX2X1 U6050 ( .B(ram[584]), .A(ram[520]), .S(n4259), .Y(n2406) );
  MUX2X1 U6051 ( .B(ram[712]), .A(ram[648]), .S(n4259), .Y(n2405) );
  MUX2X1 U6052 ( .B(ram[840]), .A(ram[776]), .S(n4259), .Y(n2409) );
  MUX2X1 U6053 ( .B(ram[968]), .A(ram[904]), .S(n4259), .Y(n2408) );
  MUX2X1 U6054 ( .B(n2407), .A(n2404), .S(n4160), .Y(n2411) );
  MUX2X1 U6055 ( .B(ram[1096]), .A(ram[1032]), .S(n4260), .Y(n2415) );
  MUX2X1 U6056 ( .B(ram[1224]), .A(ram[1160]), .S(n4260), .Y(n2414) );
  MUX2X1 U6057 ( .B(ram[1352]), .A(ram[1288]), .S(n4260), .Y(n2418) );
  MUX2X1 U6058 ( .B(ram[1480]), .A(ram[1416]), .S(n4260), .Y(n2417) );
  MUX2X1 U6059 ( .B(n2416), .A(n2413), .S(n4160), .Y(n2427) );
  MUX2X1 U6060 ( .B(ram[1608]), .A(ram[1544]), .S(n4260), .Y(n2421) );
  MUX2X1 U6061 ( .B(ram[1736]), .A(ram[1672]), .S(n4260), .Y(n2420) );
  MUX2X1 U6062 ( .B(ram[1864]), .A(ram[1800]), .S(n4260), .Y(n2424) );
  MUX2X1 U6063 ( .B(ram[1992]), .A(ram[1928]), .S(n4260), .Y(n2423) );
  MUX2X1 U6064 ( .B(n2422), .A(n2419), .S(n4160), .Y(n2426) );
  MUX2X1 U6065 ( .B(n2425), .A(n2410), .S(n4151), .Y(n4094) );
  MUX2X1 U6066 ( .B(ram[73]), .A(ram[9]), .S(n4260), .Y(n2430) );
  MUX2X1 U6067 ( .B(ram[201]), .A(ram[137]), .S(n4260), .Y(n2429) );
  MUX2X1 U6068 ( .B(ram[329]), .A(ram[265]), .S(n4260), .Y(n2433) );
  MUX2X1 U6069 ( .B(ram[457]), .A(ram[393]), .S(n4260), .Y(n2432) );
  MUX2X1 U6070 ( .B(n2431), .A(n2428), .S(n4160), .Y(n2442) );
  MUX2X1 U6071 ( .B(ram[585]), .A(ram[521]), .S(n4261), .Y(n2436) );
  MUX2X1 U6072 ( .B(ram[713]), .A(ram[649]), .S(n4261), .Y(n2435) );
  MUX2X1 U6073 ( .B(ram[841]), .A(ram[777]), .S(n4261), .Y(n2439) );
  MUX2X1 U6074 ( .B(ram[969]), .A(ram[905]), .S(n4261), .Y(n2438) );
  MUX2X1 U6075 ( .B(n2437), .A(n2434), .S(n4160), .Y(n2441) );
  MUX2X1 U6076 ( .B(ram[1097]), .A(ram[1033]), .S(n4261), .Y(n2445) );
  MUX2X1 U6077 ( .B(ram[1225]), .A(ram[1161]), .S(n4261), .Y(n2444) );
  MUX2X1 U6078 ( .B(ram[1353]), .A(ram[1289]), .S(n4261), .Y(n2448) );
  MUX2X1 U6079 ( .B(ram[1481]), .A(ram[1417]), .S(n4261), .Y(n2447) );
  MUX2X1 U6080 ( .B(n2446), .A(n2443), .S(n4160), .Y(n2457) );
  MUX2X1 U6081 ( .B(ram[1609]), .A(ram[1545]), .S(n4261), .Y(n2451) );
  MUX2X1 U6082 ( .B(ram[1737]), .A(ram[1673]), .S(n4261), .Y(n2450) );
  MUX2X1 U6083 ( .B(ram[1865]), .A(ram[1801]), .S(n4261), .Y(n2454) );
  MUX2X1 U6084 ( .B(ram[1993]), .A(ram[1929]), .S(n4261), .Y(n2453) );
  MUX2X1 U6085 ( .B(n2452), .A(n2449), .S(n4160), .Y(n2456) );
  MUX2X1 U6086 ( .B(n2455), .A(n2440), .S(n4151), .Y(n4095) );
  MUX2X1 U6087 ( .B(ram[74]), .A(ram[10]), .S(n4262), .Y(n2460) );
  MUX2X1 U6088 ( .B(ram[202]), .A(ram[138]), .S(n4262), .Y(n2459) );
  MUX2X1 U6089 ( .B(ram[330]), .A(ram[266]), .S(n4262), .Y(n2463) );
  MUX2X1 U6090 ( .B(ram[458]), .A(ram[394]), .S(n4262), .Y(n2462) );
  MUX2X1 U6091 ( .B(n2461), .A(n2458), .S(n4161), .Y(n2472) );
  MUX2X1 U6092 ( .B(ram[586]), .A(ram[522]), .S(n4262), .Y(n2466) );
  MUX2X1 U6093 ( .B(ram[714]), .A(ram[650]), .S(n4262), .Y(n2465) );
  MUX2X1 U6094 ( .B(ram[842]), .A(ram[778]), .S(n4262), .Y(n2469) );
  MUX2X1 U6095 ( .B(ram[970]), .A(ram[906]), .S(n4262), .Y(n2468) );
  MUX2X1 U6096 ( .B(n2467), .A(n2464), .S(n4161), .Y(n2471) );
  MUX2X1 U6097 ( .B(ram[1098]), .A(ram[1034]), .S(n4262), .Y(n2475) );
  MUX2X1 U6098 ( .B(ram[1226]), .A(ram[1162]), .S(n4262), .Y(n2474) );
  MUX2X1 U6099 ( .B(ram[1354]), .A(ram[1290]), .S(n4262), .Y(n2478) );
  MUX2X1 U6100 ( .B(ram[1482]), .A(ram[1418]), .S(n4262), .Y(n2477) );
  MUX2X1 U6101 ( .B(n2476), .A(n2473), .S(n4161), .Y(n2487) );
  MUX2X1 U6102 ( .B(ram[1610]), .A(ram[1546]), .S(n4263), .Y(n2481) );
  MUX2X1 U6103 ( .B(ram[1738]), .A(ram[1674]), .S(n4263), .Y(n2480) );
  MUX2X1 U6104 ( .B(ram[1866]), .A(ram[1802]), .S(n4263), .Y(n2484) );
  MUX2X1 U6105 ( .B(ram[1994]), .A(ram[1930]), .S(n4263), .Y(n2483) );
  MUX2X1 U6106 ( .B(n2482), .A(n2479), .S(n4161), .Y(n2486) );
  MUX2X1 U6107 ( .B(n2485), .A(n2470), .S(n4151), .Y(n4096) );
  MUX2X1 U6108 ( .B(ram[75]), .A(ram[11]), .S(n4263), .Y(n2490) );
  MUX2X1 U6109 ( .B(ram[203]), .A(ram[139]), .S(n4263), .Y(n2489) );
  MUX2X1 U6110 ( .B(ram[331]), .A(ram[267]), .S(n4263), .Y(n2493) );
  MUX2X1 U6111 ( .B(ram[459]), .A(ram[395]), .S(n4263), .Y(n2492) );
  MUX2X1 U6112 ( .B(n2491), .A(n2488), .S(n4161), .Y(n2502) );
  MUX2X1 U6113 ( .B(ram[587]), .A(ram[523]), .S(n4263), .Y(n2496) );
  MUX2X1 U6114 ( .B(ram[715]), .A(ram[651]), .S(n4263), .Y(n2495) );
  MUX2X1 U6115 ( .B(ram[843]), .A(ram[779]), .S(n4263), .Y(n2499) );
  MUX2X1 U6116 ( .B(ram[971]), .A(ram[907]), .S(n4263), .Y(n2498) );
  MUX2X1 U6117 ( .B(n2497), .A(n2494), .S(n4161), .Y(n2501) );
  MUX2X1 U6118 ( .B(ram[1099]), .A(ram[1035]), .S(n4264), .Y(n2505) );
  MUX2X1 U6119 ( .B(ram[1227]), .A(ram[1163]), .S(n4264), .Y(n2504) );
  MUX2X1 U6120 ( .B(ram[1355]), .A(ram[1291]), .S(n4264), .Y(n2508) );
  MUX2X1 U6121 ( .B(ram[1483]), .A(ram[1419]), .S(n4264), .Y(n2507) );
  MUX2X1 U6122 ( .B(n2506), .A(n2503), .S(n4161), .Y(n2518) );
  MUX2X1 U6123 ( .B(ram[1611]), .A(ram[1547]), .S(n4264), .Y(n2511) );
  MUX2X1 U6124 ( .B(ram[1739]), .A(ram[1675]), .S(n4264), .Y(n2510) );
  MUX2X1 U6125 ( .B(ram[1867]), .A(ram[1803]), .S(n4264), .Y(n2514) );
  MUX2X1 U6126 ( .B(ram[1995]), .A(ram[1931]), .S(n4264), .Y(n2513) );
  MUX2X1 U6127 ( .B(n2512), .A(n2509), .S(n4161), .Y(n2516) );
  MUX2X1 U6128 ( .B(n2515), .A(n2500), .S(n4152), .Y(n4097) );
  MUX2X1 U6129 ( .B(ram[76]), .A(ram[12]), .S(n4264), .Y(n2521) );
  MUX2X1 U6130 ( .B(ram[204]), .A(ram[140]), .S(n4264), .Y(n2520) );
  MUX2X1 U6131 ( .B(ram[332]), .A(ram[268]), .S(n4264), .Y(n2524) );
  MUX2X1 U6132 ( .B(ram[460]), .A(ram[396]), .S(n4264), .Y(n2523) );
  MUX2X1 U6133 ( .B(n2522), .A(n2519), .S(n4161), .Y(n2533) );
  MUX2X1 U6134 ( .B(ram[588]), .A(ram[524]), .S(n4265), .Y(n2527) );
  MUX2X1 U6135 ( .B(ram[716]), .A(ram[652]), .S(n4265), .Y(n2526) );
  MUX2X1 U6136 ( .B(ram[844]), .A(ram[780]), .S(n4265), .Y(n2530) );
  MUX2X1 U6137 ( .B(ram[972]), .A(ram[908]), .S(n4265), .Y(n2529) );
  MUX2X1 U6138 ( .B(n2528), .A(n2525), .S(n4161), .Y(n2532) );
  MUX2X1 U6139 ( .B(ram[1100]), .A(ram[1036]), .S(n4265), .Y(n2536) );
  MUX2X1 U6140 ( .B(ram[1228]), .A(ram[1164]), .S(n4265), .Y(n2535) );
  MUX2X1 U6141 ( .B(ram[1356]), .A(ram[1292]), .S(n4265), .Y(n2539) );
  MUX2X1 U6142 ( .B(ram[1484]), .A(ram[1420]), .S(n4265), .Y(n2538) );
  MUX2X1 U6143 ( .B(n2537), .A(n2534), .S(n4161), .Y(n2548) );
  MUX2X1 U6144 ( .B(ram[1612]), .A(ram[1548]), .S(n4265), .Y(n2542) );
  MUX2X1 U6145 ( .B(ram[1740]), .A(ram[1676]), .S(n4265), .Y(n2541) );
  MUX2X1 U6146 ( .B(ram[1868]), .A(ram[1804]), .S(n4265), .Y(n2545) );
  MUX2X1 U6147 ( .B(ram[1996]), .A(ram[1932]), .S(n4265), .Y(n2544) );
  MUX2X1 U6148 ( .B(n2543), .A(n2540), .S(n4161), .Y(n2547) );
  MUX2X1 U6149 ( .B(n2546), .A(n2531), .S(n4152), .Y(n4098) );
  MUX2X1 U6150 ( .B(ram[77]), .A(ram[13]), .S(n4266), .Y(n2551) );
  MUX2X1 U6151 ( .B(ram[205]), .A(ram[141]), .S(n4266), .Y(n2550) );
  MUX2X1 U6152 ( .B(ram[333]), .A(ram[269]), .S(n4266), .Y(n2554) );
  MUX2X1 U6153 ( .B(ram[461]), .A(ram[397]), .S(n4266), .Y(n2553) );
  MUX2X1 U6154 ( .B(n2552), .A(n2549), .S(n4162), .Y(n2563) );
  MUX2X1 U6155 ( .B(ram[589]), .A(ram[525]), .S(n4266), .Y(n2557) );
  MUX2X1 U6156 ( .B(ram[717]), .A(ram[653]), .S(n4266), .Y(n2556) );
  MUX2X1 U6157 ( .B(ram[845]), .A(ram[781]), .S(n4266), .Y(n2560) );
  MUX2X1 U6158 ( .B(ram[973]), .A(ram[909]), .S(n4266), .Y(n2559) );
  MUX2X1 U6159 ( .B(n2558), .A(n2555), .S(n4162), .Y(n2562) );
  MUX2X1 U6160 ( .B(ram[1101]), .A(ram[1037]), .S(n4266), .Y(n2566) );
  MUX2X1 U6161 ( .B(ram[1229]), .A(ram[1165]), .S(n4266), .Y(n2565) );
  MUX2X1 U6162 ( .B(ram[1357]), .A(ram[1293]), .S(n4266), .Y(n2569) );
  MUX2X1 U6163 ( .B(ram[1485]), .A(ram[1421]), .S(n4266), .Y(n2568) );
  MUX2X1 U6164 ( .B(n2567), .A(n2564), .S(n4162), .Y(n2578) );
  MUX2X1 U6165 ( .B(ram[1613]), .A(ram[1549]), .S(n4267), .Y(n2572) );
  MUX2X1 U6166 ( .B(ram[1741]), .A(ram[1677]), .S(n4267), .Y(n2571) );
  MUX2X1 U6167 ( .B(ram[1869]), .A(ram[1805]), .S(n4267), .Y(n2575) );
  MUX2X1 U6168 ( .B(ram[1997]), .A(ram[1933]), .S(n4267), .Y(n2574) );
  MUX2X1 U6169 ( .B(n2573), .A(n2570), .S(n4162), .Y(n2577) );
  MUX2X1 U6170 ( .B(n2576), .A(n2561), .S(n4152), .Y(n4099) );
  MUX2X1 U6171 ( .B(ram[78]), .A(ram[14]), .S(n4267), .Y(n2581) );
  MUX2X1 U6172 ( .B(ram[206]), .A(ram[142]), .S(n4267), .Y(n2580) );
  MUX2X1 U6173 ( .B(ram[334]), .A(ram[270]), .S(n4267), .Y(n2585) );
  MUX2X1 U6174 ( .B(ram[462]), .A(ram[398]), .S(n4267), .Y(n2583) );
  MUX2X1 U6175 ( .B(n2582), .A(n2579), .S(n4162), .Y(n2594) );
  MUX2X1 U6176 ( .B(ram[590]), .A(ram[526]), .S(n4267), .Y(n2588) );
  MUX2X1 U6177 ( .B(ram[718]), .A(ram[654]), .S(n4267), .Y(n2587) );
  MUX2X1 U6178 ( .B(ram[846]), .A(ram[782]), .S(n4267), .Y(n2591) );
  MUX2X1 U6179 ( .B(ram[974]), .A(ram[910]), .S(n4267), .Y(n2590) );
  MUX2X1 U6180 ( .B(n2589), .A(n2586), .S(n4162), .Y(n2593) );
  MUX2X1 U6181 ( .B(ram[1102]), .A(ram[1038]), .S(n4268), .Y(n2597) );
  MUX2X1 U6182 ( .B(ram[1230]), .A(ram[1166]), .S(n4268), .Y(n2596) );
  MUX2X1 U6183 ( .B(ram[1358]), .A(ram[1294]), .S(n4268), .Y(n2600) );
  MUX2X1 U6184 ( .B(ram[1486]), .A(ram[1422]), .S(n4268), .Y(n2599) );
  MUX2X1 U6185 ( .B(n2598), .A(n2595), .S(n4162), .Y(n2609) );
  MUX2X1 U6186 ( .B(ram[1614]), .A(ram[1550]), .S(n4268), .Y(n2603) );
  MUX2X1 U6187 ( .B(ram[1742]), .A(ram[1678]), .S(n4268), .Y(n2602) );
  MUX2X1 U6188 ( .B(ram[1870]), .A(ram[1806]), .S(n4268), .Y(n2606) );
  MUX2X1 U6189 ( .B(ram[1998]), .A(ram[1934]), .S(n4268), .Y(n2605) );
  MUX2X1 U6190 ( .B(n2604), .A(n2601), .S(n4162), .Y(n2608) );
  MUX2X1 U6191 ( .B(n2607), .A(n2592), .S(n4152), .Y(n4100) );
  MUX2X1 U6192 ( .B(ram[79]), .A(ram[15]), .S(n4268), .Y(n2612) );
  MUX2X1 U6193 ( .B(ram[207]), .A(ram[143]), .S(n4268), .Y(n2611) );
  MUX2X1 U6194 ( .B(ram[335]), .A(ram[271]), .S(n4268), .Y(n2615) );
  MUX2X1 U6195 ( .B(ram[463]), .A(ram[399]), .S(n4268), .Y(n2614) );
  MUX2X1 U6196 ( .B(n2613), .A(n2610), .S(n4162), .Y(n2624) );
  MUX2X1 U6197 ( .B(ram[591]), .A(ram[527]), .S(n4269), .Y(n2618) );
  MUX2X1 U6198 ( .B(ram[719]), .A(ram[655]), .S(n4269), .Y(n2617) );
  MUX2X1 U6199 ( .B(ram[847]), .A(ram[783]), .S(n4269), .Y(n2621) );
  MUX2X1 U6200 ( .B(ram[975]), .A(ram[911]), .S(n4269), .Y(n2620) );
  MUX2X1 U6201 ( .B(n2619), .A(n2616), .S(n4162), .Y(n2623) );
  MUX2X1 U6202 ( .B(ram[1103]), .A(ram[1039]), .S(n4269), .Y(n2627) );
  MUX2X1 U6203 ( .B(ram[1231]), .A(ram[1167]), .S(n4269), .Y(n2626) );
  MUX2X1 U6204 ( .B(ram[1359]), .A(ram[1295]), .S(n4269), .Y(n2630) );
  MUX2X1 U6205 ( .B(ram[1487]), .A(ram[1423]), .S(n4269), .Y(n2629) );
  MUX2X1 U6206 ( .B(n2628), .A(n2625), .S(n4162), .Y(n2639) );
  MUX2X1 U6207 ( .B(ram[1615]), .A(ram[1551]), .S(n4269), .Y(n2633) );
  MUX2X1 U6208 ( .B(ram[1743]), .A(ram[1679]), .S(n4269), .Y(n2632) );
  MUX2X1 U6209 ( .B(ram[1871]), .A(ram[1807]), .S(n4269), .Y(n2636) );
  MUX2X1 U6210 ( .B(ram[1999]), .A(ram[1935]), .S(n4269), .Y(n2635) );
  MUX2X1 U6211 ( .B(n2634), .A(n2631), .S(n4162), .Y(n2638) );
  MUX2X1 U6212 ( .B(n2637), .A(n2622), .S(n4152), .Y(n4101) );
  MUX2X1 U6213 ( .B(ram[80]), .A(ram[16]), .S(n4270), .Y(n2642) );
  MUX2X1 U6214 ( .B(ram[208]), .A(ram[144]), .S(n4270), .Y(n2641) );
  MUX2X1 U6215 ( .B(ram[336]), .A(ram[272]), .S(n4270), .Y(n2645) );
  MUX2X1 U6216 ( .B(ram[464]), .A(ram[400]), .S(n4270), .Y(n2644) );
  MUX2X1 U6217 ( .B(n2643), .A(n2640), .S(n4164), .Y(n2655) );
  MUX2X1 U6218 ( .B(ram[592]), .A(ram[528]), .S(n4270), .Y(n2648) );
  MUX2X1 U6219 ( .B(ram[720]), .A(ram[656]), .S(n4270), .Y(n2647) );
  MUX2X1 U6220 ( .B(ram[848]), .A(ram[784]), .S(n4270), .Y(n2652) );
  MUX2X1 U6221 ( .B(ram[976]), .A(ram[912]), .S(n4270), .Y(n2650) );
  MUX2X1 U6222 ( .B(n2649), .A(n2646), .S(n4161), .Y(n2654) );
  MUX2X1 U6223 ( .B(ram[1104]), .A(ram[1040]), .S(n4270), .Y(n2658) );
  MUX2X1 U6224 ( .B(ram[1232]), .A(ram[1168]), .S(n4270), .Y(n2657) );
  MUX2X1 U6225 ( .B(ram[1360]), .A(ram[1296]), .S(n4270), .Y(n2661) );
  MUX2X1 U6226 ( .B(ram[1488]), .A(ram[1424]), .S(n4270), .Y(n2660) );
  MUX2X1 U6227 ( .B(n2659), .A(n2656), .S(n4159), .Y(n2670) );
  MUX2X1 U6228 ( .B(ram[1616]), .A(ram[1552]), .S(n4271), .Y(n2664) );
  MUX2X1 U6229 ( .B(ram[1744]), .A(ram[1680]), .S(n4271), .Y(n2663) );
  MUX2X1 U6230 ( .B(ram[1872]), .A(ram[1808]), .S(n4271), .Y(n2667) );
  MUX2X1 U6231 ( .B(ram[2000]), .A(ram[1936]), .S(n4271), .Y(n2666) );
  MUX2X1 U6232 ( .B(n2665), .A(n2662), .S(n4166), .Y(n2669) );
  MUX2X1 U6233 ( .B(n2668), .A(n2653), .S(n4152), .Y(n4102) );
  MUX2X1 U6234 ( .B(ram[81]), .A(ram[17]), .S(n4271), .Y(n2673) );
  MUX2X1 U6235 ( .B(ram[209]), .A(ram[145]), .S(n4271), .Y(n2672) );
  MUX2X1 U6236 ( .B(ram[337]), .A(ram[273]), .S(n4271), .Y(n2676) );
  MUX2X1 U6237 ( .B(ram[465]), .A(ram[401]), .S(n4271), .Y(n2675) );
  MUX2X1 U6238 ( .B(n2674), .A(n2671), .S(n4158), .Y(n2685) );
  MUX2X1 U6239 ( .B(ram[593]), .A(ram[529]), .S(n4271), .Y(n2679) );
  MUX2X1 U6240 ( .B(ram[721]), .A(ram[657]), .S(n4271), .Y(n2678) );
  MUX2X1 U6241 ( .B(ram[849]), .A(ram[785]), .S(n4271), .Y(n2682) );
  MUX2X1 U6242 ( .B(ram[977]), .A(ram[913]), .S(n4271), .Y(n2681) );
  MUX2X1 U6243 ( .B(n2680), .A(n2677), .S(n4167), .Y(n2684) );
  MUX2X1 U6244 ( .B(ram[1105]), .A(ram[1041]), .S(n4272), .Y(n2688) );
  MUX2X1 U6245 ( .B(ram[1233]), .A(ram[1169]), .S(n4272), .Y(n2687) );
  MUX2X1 U6246 ( .B(ram[1361]), .A(ram[1297]), .S(n4272), .Y(n2691) );
  MUX2X1 U6247 ( .B(ram[1489]), .A(ram[1425]), .S(n4272), .Y(n2690) );
  MUX2X1 U6248 ( .B(n2689), .A(n2686), .S(n4158), .Y(n2700) );
  MUX2X1 U6249 ( .B(ram[1617]), .A(ram[1553]), .S(n4272), .Y(n2694) );
  MUX2X1 U6250 ( .B(ram[1745]), .A(ram[1681]), .S(n4272), .Y(n2693) );
  MUX2X1 U6251 ( .B(ram[1873]), .A(ram[1809]), .S(n4272), .Y(n2697) );
  MUX2X1 U6252 ( .B(ram[2001]), .A(ram[1937]), .S(n4272), .Y(n2696) );
  MUX2X1 U6253 ( .B(n2695), .A(n2692), .S(n4159), .Y(n2699) );
  MUX2X1 U6254 ( .B(n2698), .A(n2683), .S(n4152), .Y(n4103) );
  MUX2X1 U6255 ( .B(ram[82]), .A(ram[18]), .S(n4272), .Y(n2703) );
  MUX2X1 U6256 ( .B(ram[210]), .A(ram[146]), .S(n4272), .Y(n2702) );
  MUX2X1 U6257 ( .B(ram[338]), .A(ram[274]), .S(n4272), .Y(n2706) );
  MUX2X1 U6258 ( .B(ram[466]), .A(ram[402]), .S(n4272), .Y(n2705) );
  MUX2X1 U6259 ( .B(n2704), .A(n2701), .S(n4169), .Y(n2715) );
  MUX2X1 U6260 ( .B(ram[594]), .A(ram[530]), .S(n4273), .Y(n2709) );
  MUX2X1 U6261 ( .B(ram[722]), .A(ram[658]), .S(n4273), .Y(n2708) );
  MUX2X1 U6262 ( .B(ram[850]), .A(ram[786]), .S(n4273), .Y(n2712) );
  MUX2X1 U6263 ( .B(ram[978]), .A(ram[914]), .S(n4273), .Y(n2711) );
  MUX2X1 U6264 ( .B(n2710), .A(n2707), .S(n4174), .Y(n2714) );
  MUX2X1 U6265 ( .B(ram[1106]), .A(ram[1042]), .S(n4273), .Y(n2719) );
  MUX2X1 U6266 ( .B(ram[1234]), .A(ram[1170]), .S(n4273), .Y(n2717) );
  MUX2X1 U6267 ( .B(ram[1362]), .A(ram[1298]), .S(n4273), .Y(n2722) );
  MUX2X1 U6268 ( .B(ram[1490]), .A(ram[1426]), .S(n4273), .Y(n2721) );
  MUX2X1 U6269 ( .B(n2720), .A(n2716), .S(n4171), .Y(n2731) );
  MUX2X1 U6270 ( .B(ram[1618]), .A(ram[1554]), .S(n4273), .Y(n2725) );
  MUX2X1 U6271 ( .B(ram[1746]), .A(ram[1682]), .S(n4273), .Y(n2724) );
  MUX2X1 U6272 ( .B(ram[1874]), .A(ram[1810]), .S(n4273), .Y(n2728) );
  MUX2X1 U6273 ( .B(ram[2002]), .A(ram[1938]), .S(n4273), .Y(n2727) );
  MUX2X1 U6274 ( .B(n2726), .A(n2723), .S(n4172), .Y(n2730) );
  MUX2X1 U6275 ( .B(n2729), .A(n2713), .S(n4152), .Y(n4104) );
  MUX2X1 U6276 ( .B(ram[83]), .A(ram[19]), .S(n4274), .Y(n2734) );
  MUX2X1 U6277 ( .B(ram[211]), .A(ram[147]), .S(n4274), .Y(n2733) );
  MUX2X1 U6278 ( .B(ram[339]), .A(ram[275]), .S(n4274), .Y(n2737) );
  MUX2X1 U6279 ( .B(ram[467]), .A(ram[403]), .S(n4274), .Y(n2736) );
  MUX2X1 U6280 ( .B(n2735), .A(n2732), .S(n4163), .Y(n2746) );
  MUX2X1 U6281 ( .B(ram[595]), .A(ram[531]), .S(n4274), .Y(n2740) );
  MUX2X1 U6282 ( .B(ram[723]), .A(ram[659]), .S(n4274), .Y(n2739) );
  MUX2X1 U6283 ( .B(ram[851]), .A(ram[787]), .S(n4274), .Y(n2743) );
  MUX2X1 U6284 ( .B(ram[979]), .A(ram[915]), .S(n4274), .Y(n2742) );
  MUX2X1 U6285 ( .B(n2741), .A(n2738), .S(n4163), .Y(n2745) );
  MUX2X1 U6286 ( .B(ram[1107]), .A(ram[1043]), .S(n4274), .Y(n2749) );
  MUX2X1 U6287 ( .B(ram[1235]), .A(ram[1171]), .S(n4274), .Y(n2748) );
  MUX2X1 U6288 ( .B(ram[1363]), .A(ram[1299]), .S(n4274), .Y(n2752) );
  MUX2X1 U6289 ( .B(ram[1491]), .A(ram[1427]), .S(n4274), .Y(n2751) );
  MUX2X1 U6290 ( .B(n2750), .A(n2747), .S(n4163), .Y(n2761) );
  MUX2X1 U6291 ( .B(ram[1619]), .A(ram[1555]), .S(n4275), .Y(n2755) );
  MUX2X1 U6292 ( .B(ram[1747]), .A(ram[1683]), .S(n4275), .Y(n2754) );
  MUX2X1 U6293 ( .B(ram[1875]), .A(ram[1811]), .S(n4275), .Y(n2758) );
  MUX2X1 U6294 ( .B(ram[2003]), .A(ram[1939]), .S(n4275), .Y(n2757) );
  MUX2X1 U6295 ( .B(n2756), .A(n2753), .S(n4163), .Y(n2760) );
  MUX2X1 U6296 ( .B(n2759), .A(n2744), .S(n4152), .Y(n4105) );
  MUX2X1 U6297 ( .B(ram[84]), .A(ram[20]), .S(n4275), .Y(n2764) );
  MUX2X1 U6298 ( .B(ram[212]), .A(ram[148]), .S(n4275), .Y(n2763) );
  MUX2X1 U6299 ( .B(ram[340]), .A(ram[276]), .S(n4275), .Y(n2767) );
  MUX2X1 U6300 ( .B(ram[468]), .A(ram[404]), .S(n4275), .Y(n2766) );
  MUX2X1 U6301 ( .B(n2765), .A(n2762), .S(n4163), .Y(n2776) );
  MUX2X1 U6302 ( .B(ram[596]), .A(ram[532]), .S(n4275), .Y(n2770) );
  MUX2X1 U6303 ( .B(ram[724]), .A(ram[660]), .S(n4275), .Y(n2769) );
  MUX2X1 U6304 ( .B(ram[852]), .A(ram[788]), .S(n4275), .Y(n2773) );
  MUX2X1 U6305 ( .B(ram[980]), .A(ram[916]), .S(n4275), .Y(n2772) );
  MUX2X1 U6306 ( .B(n2771), .A(n2768), .S(n4163), .Y(n2775) );
  MUX2X1 U6307 ( .B(ram[1108]), .A(ram[1044]), .S(n4276), .Y(n2779) );
  MUX2X1 U6308 ( .B(ram[1236]), .A(ram[1172]), .S(n4276), .Y(n2778) );
  MUX2X1 U6309 ( .B(ram[1364]), .A(ram[1300]), .S(n4276), .Y(n2782) );
  MUX2X1 U6310 ( .B(ram[1492]), .A(ram[1428]), .S(n4276), .Y(n2781) );
  MUX2X1 U6311 ( .B(n2780), .A(n2777), .S(n4163), .Y(n2792) );
  MUX2X1 U6312 ( .B(ram[1620]), .A(ram[1556]), .S(n4276), .Y(n2786) );
  MUX2X1 U6313 ( .B(ram[1748]), .A(ram[1684]), .S(n4276), .Y(n2784) );
  MUX2X1 U6314 ( .B(ram[1876]), .A(ram[1812]), .S(n4276), .Y(n2789) );
  MUX2X1 U6315 ( .B(ram[2004]), .A(ram[1940]), .S(n4276), .Y(n2788) );
  MUX2X1 U6316 ( .B(n2787), .A(n2783), .S(n4163), .Y(n2791) );
  MUX2X1 U6317 ( .B(n2790), .A(n2774), .S(n4152), .Y(n4106) );
  MUX2X1 U6318 ( .B(ram[85]), .A(ram[21]), .S(n4276), .Y(n2795) );
  MUX2X1 U6319 ( .B(ram[213]), .A(ram[149]), .S(n4276), .Y(n2794) );
  MUX2X1 U6320 ( .B(ram[341]), .A(ram[277]), .S(n4276), .Y(n2798) );
  MUX2X1 U6321 ( .B(ram[469]), .A(ram[405]), .S(n4276), .Y(n2797) );
  MUX2X1 U6322 ( .B(n2796), .A(n2793), .S(n4163), .Y(n2807) );
  MUX2X1 U6323 ( .B(ram[597]), .A(ram[533]), .S(n4277), .Y(n2801) );
  MUX2X1 U6324 ( .B(ram[725]), .A(ram[661]), .S(n4277), .Y(n2800) );
  MUX2X1 U6325 ( .B(ram[853]), .A(ram[789]), .S(n4277), .Y(n2804) );
  MUX2X1 U6326 ( .B(ram[981]), .A(ram[917]), .S(n4277), .Y(n2803) );
  MUX2X1 U6327 ( .B(n2802), .A(n2799), .S(n4163), .Y(n2806) );
  MUX2X1 U6328 ( .B(ram[1109]), .A(ram[1045]), .S(n4277), .Y(n2810) );
  MUX2X1 U6329 ( .B(ram[1237]), .A(ram[1173]), .S(n4277), .Y(n2809) );
  MUX2X1 U6330 ( .B(ram[1365]), .A(ram[1301]), .S(n4277), .Y(n2813) );
  MUX2X1 U6331 ( .B(ram[1493]), .A(ram[1429]), .S(n4277), .Y(n2812) );
  MUX2X1 U6332 ( .B(n2811), .A(n2808), .S(n4163), .Y(n2822) );
  MUX2X1 U6333 ( .B(ram[1621]), .A(ram[1557]), .S(n4277), .Y(n2816) );
  MUX2X1 U6334 ( .B(ram[1749]), .A(ram[1685]), .S(n4277), .Y(n2815) );
  MUX2X1 U6335 ( .B(ram[1877]), .A(ram[1813]), .S(n4277), .Y(n2819) );
  MUX2X1 U6336 ( .B(ram[2005]), .A(ram[1941]), .S(n4277), .Y(n2818) );
  MUX2X1 U6337 ( .B(n2817), .A(n2814), .S(n4163), .Y(n2821) );
  MUX2X1 U6338 ( .B(n2820), .A(n2805), .S(n4152), .Y(n4107) );
  MUX2X1 U6339 ( .B(ram[86]), .A(ram[22]), .S(n4278), .Y(n2825) );
  MUX2X1 U6340 ( .B(ram[214]), .A(ram[150]), .S(n4278), .Y(n2824) );
  MUX2X1 U6341 ( .B(ram[342]), .A(ram[278]), .S(n4278), .Y(n2828) );
  MUX2X1 U6342 ( .B(ram[470]), .A(ram[406]), .S(n4278), .Y(n2827) );
  MUX2X1 U6343 ( .B(n2826), .A(n2823), .S(n4164), .Y(n2837) );
  MUX2X1 U6344 ( .B(ram[598]), .A(ram[534]), .S(n4278), .Y(n2831) );
  MUX2X1 U6345 ( .B(ram[726]), .A(ram[662]), .S(n4278), .Y(n2830) );
  MUX2X1 U6346 ( .B(ram[854]), .A(ram[790]), .S(n4278), .Y(n2834) );
  MUX2X1 U6347 ( .B(ram[982]), .A(ram[918]), .S(n4278), .Y(n2833) );
  MUX2X1 U6348 ( .B(n2832), .A(n2829), .S(n4164), .Y(n2836) );
  MUX2X1 U6349 ( .B(ram[1110]), .A(ram[1046]), .S(n4278), .Y(n2840) );
  MUX2X1 U6350 ( .B(ram[1238]), .A(ram[1174]), .S(n4278), .Y(n2839) );
  MUX2X1 U6351 ( .B(ram[1366]), .A(ram[1302]), .S(n4278), .Y(n2843) );
  MUX2X1 U6352 ( .B(ram[1494]), .A(ram[1430]), .S(n4278), .Y(n2842) );
  MUX2X1 U6353 ( .B(n2841), .A(n2838), .S(n4164), .Y(n2853) );
  MUX2X1 U6354 ( .B(ram[1622]), .A(ram[1558]), .S(n4279), .Y(n2846) );
  MUX2X1 U6355 ( .B(ram[1750]), .A(ram[1686]), .S(n4279), .Y(n2845) );
  MUX2X1 U6356 ( .B(ram[1878]), .A(ram[1814]), .S(n4279), .Y(n2849) );
  MUX2X1 U6357 ( .B(ram[2006]), .A(ram[1942]), .S(n4279), .Y(n2848) );
  MUX2X1 U6358 ( .B(n2847), .A(n2844), .S(n4164), .Y(n2851) );
  MUX2X1 U6359 ( .B(n2850), .A(n2835), .S(n4152), .Y(n4108) );
  MUX2X1 U6360 ( .B(ram[87]), .A(ram[23]), .S(n4279), .Y(n2856) );
  MUX2X1 U6361 ( .B(ram[215]), .A(ram[151]), .S(n4279), .Y(n2855) );
  MUX2X1 U6362 ( .B(ram[343]), .A(ram[279]), .S(n4279), .Y(n2859) );
  MUX2X1 U6363 ( .B(ram[471]), .A(ram[407]), .S(n4279), .Y(n2858) );
  MUX2X1 U6364 ( .B(n2857), .A(n2854), .S(n4164), .Y(n2868) );
  MUX2X1 U6365 ( .B(ram[599]), .A(ram[535]), .S(n4279), .Y(n2862) );
  MUX2X1 U6366 ( .B(ram[727]), .A(ram[663]), .S(n4279), .Y(n2861) );
  MUX2X1 U6367 ( .B(ram[855]), .A(ram[791]), .S(n4279), .Y(n2865) );
  MUX2X1 U6368 ( .B(ram[983]), .A(ram[919]), .S(n4279), .Y(n2864) );
  MUX2X1 U6369 ( .B(n2863), .A(n2860), .S(n4164), .Y(n2867) );
  MUX2X1 U6370 ( .B(ram[1111]), .A(ram[1047]), .S(n4280), .Y(n2871) );
  MUX2X1 U6371 ( .B(ram[1239]), .A(ram[1175]), .S(n4280), .Y(n2870) );
  MUX2X1 U6372 ( .B(ram[1367]), .A(ram[1303]), .S(n4280), .Y(n2874) );
  MUX2X1 U6373 ( .B(ram[1495]), .A(ram[1431]), .S(n4280), .Y(n2873) );
  MUX2X1 U6374 ( .B(n2872), .A(n2869), .S(n4164), .Y(n2883) );
  MUX2X1 U6375 ( .B(ram[1623]), .A(ram[1559]), .S(n4280), .Y(n2877) );
  MUX2X1 U6376 ( .B(ram[1751]), .A(ram[1687]), .S(n4280), .Y(n2876) );
  MUX2X1 U6377 ( .B(ram[1879]), .A(ram[1815]), .S(n4280), .Y(n2880) );
  MUX2X1 U6378 ( .B(ram[2007]), .A(ram[1943]), .S(n4280), .Y(n2879) );
  MUX2X1 U6379 ( .B(n2878), .A(n2875), .S(n4164), .Y(n2882) );
  MUX2X1 U6380 ( .B(n2881), .A(n2866), .S(n4152), .Y(n4109) );
  MUX2X1 U6381 ( .B(ram[88]), .A(ram[24]), .S(n4280), .Y(n2886) );
  MUX2X1 U6382 ( .B(ram[216]), .A(ram[152]), .S(n4280), .Y(n2885) );
  MUX2X1 U6383 ( .B(ram[344]), .A(ram[280]), .S(n4280), .Y(n2889) );
  MUX2X1 U6384 ( .B(ram[472]), .A(ram[408]), .S(n4280), .Y(n2888) );
  MUX2X1 U6385 ( .B(n2887), .A(n2884), .S(n4164), .Y(n2898) );
  MUX2X1 U6386 ( .B(ram[600]), .A(ram[536]), .S(n4281), .Y(n2892) );
  MUX2X1 U6387 ( .B(ram[728]), .A(ram[664]), .S(n4281), .Y(n2891) );
  MUX2X1 U6388 ( .B(ram[856]), .A(ram[792]), .S(n4281), .Y(n2895) );
  MUX2X1 U6389 ( .B(ram[984]), .A(ram[920]), .S(n4281), .Y(n2894) );
  MUX2X1 U6390 ( .B(n2893), .A(n2890), .S(n4164), .Y(n2897) );
  MUX2X1 U6391 ( .B(ram[1112]), .A(ram[1048]), .S(n4281), .Y(n2901) );
  MUX2X1 U6392 ( .B(ram[1240]), .A(ram[1176]), .S(n4281), .Y(n2900) );
  MUX2X1 U6393 ( .B(ram[1368]), .A(ram[1304]), .S(n4281), .Y(n2904) );
  MUX2X1 U6394 ( .B(ram[1496]), .A(ram[1432]), .S(n4281), .Y(n2903) );
  MUX2X1 U6395 ( .B(n2902), .A(n2899), .S(n4164), .Y(n2913) );
  MUX2X1 U6396 ( .B(ram[1624]), .A(ram[1560]), .S(n4281), .Y(n2907) );
  MUX2X1 U6397 ( .B(ram[1752]), .A(ram[1688]), .S(n4281), .Y(n2906) );
  MUX2X1 U6398 ( .B(ram[1880]), .A(ram[1816]), .S(n4281), .Y(n2910) );
  MUX2X1 U6399 ( .B(ram[2008]), .A(ram[1944]), .S(n4281), .Y(n2909) );
  MUX2X1 U6400 ( .B(n2908), .A(n2905), .S(n4164), .Y(n2912) );
  MUX2X1 U6401 ( .B(n2911), .A(n2896), .S(n4152), .Y(n4110) );
  MUX2X1 U6402 ( .B(ram[89]), .A(ram[25]), .S(n4282), .Y(n2916) );
  MUX2X1 U6403 ( .B(ram[217]), .A(ram[153]), .S(n4282), .Y(n2915) );
  MUX2X1 U6404 ( .B(ram[345]), .A(ram[281]), .S(n4282), .Y(n2920) );
  MUX2X1 U6405 ( .B(ram[473]), .A(ram[409]), .S(n4282), .Y(n2918) );
  MUX2X1 U6406 ( .B(n2917), .A(n2914), .S(n4165), .Y(n2929) );
  MUX2X1 U6407 ( .B(ram[601]), .A(ram[537]), .S(n4282), .Y(n2923) );
  MUX2X1 U6408 ( .B(ram[729]), .A(ram[665]), .S(n4282), .Y(n2922) );
  MUX2X1 U6409 ( .B(ram[857]), .A(ram[793]), .S(n4282), .Y(n2926) );
  MUX2X1 U6410 ( .B(ram[985]), .A(ram[921]), .S(n4282), .Y(n2925) );
  MUX2X1 U6411 ( .B(n2924), .A(n2921), .S(n4165), .Y(n2928) );
  MUX2X1 U6412 ( .B(ram[1113]), .A(ram[1049]), .S(n4282), .Y(n2932) );
  MUX2X1 U6413 ( .B(ram[1241]), .A(ram[1177]), .S(n4282), .Y(n2931) );
  MUX2X1 U6414 ( .B(ram[1369]), .A(ram[1305]), .S(n4282), .Y(n2935) );
  MUX2X1 U6415 ( .B(ram[1497]), .A(ram[1433]), .S(n4282), .Y(n2934) );
  MUX2X1 U6416 ( .B(n2933), .A(n2930), .S(n4165), .Y(n2944) );
  MUX2X1 U6417 ( .B(ram[1625]), .A(ram[1561]), .S(n4283), .Y(n2938) );
  MUX2X1 U6418 ( .B(ram[1753]), .A(ram[1689]), .S(n4283), .Y(n2937) );
  MUX2X1 U6419 ( .B(ram[1881]), .A(ram[1817]), .S(n4283), .Y(n2941) );
  MUX2X1 U6420 ( .B(ram[2009]), .A(ram[1945]), .S(n4283), .Y(n2940) );
  MUX2X1 U6421 ( .B(n2939), .A(n2936), .S(n4165), .Y(n2943) );
  MUX2X1 U6422 ( .B(n2942), .A(n2927), .S(n4152), .Y(n4111) );
  MUX2X1 U6423 ( .B(ram[90]), .A(ram[26]), .S(n4283), .Y(n2947) );
  MUX2X1 U6424 ( .B(ram[218]), .A(ram[154]), .S(n4283), .Y(n2946) );
  MUX2X1 U6425 ( .B(ram[346]), .A(ram[282]), .S(n4283), .Y(n2950) );
  MUX2X1 U6426 ( .B(ram[474]), .A(ram[410]), .S(n4283), .Y(n2949) );
  MUX2X1 U6427 ( .B(n2948), .A(n2945), .S(n4165), .Y(n2959) );
  MUX2X1 U6428 ( .B(ram[602]), .A(ram[538]), .S(n4283), .Y(n2953) );
  MUX2X1 U6429 ( .B(ram[730]), .A(ram[666]), .S(n4283), .Y(n2952) );
  MUX2X1 U6430 ( .B(ram[858]), .A(ram[794]), .S(n4283), .Y(n2956) );
  MUX2X1 U6431 ( .B(ram[986]), .A(ram[922]), .S(n4283), .Y(n2955) );
  MUX2X1 U6432 ( .B(n2954), .A(n2951), .S(n4165), .Y(n2958) );
  MUX2X1 U6433 ( .B(ram[1114]), .A(ram[1050]), .S(n4284), .Y(n2962) );
  MUX2X1 U6434 ( .B(ram[1242]), .A(ram[1178]), .S(n4284), .Y(n2961) );
  MUX2X1 U6435 ( .B(ram[1370]), .A(ram[1306]), .S(n4284), .Y(n2965) );
  MUX2X1 U6436 ( .B(ram[1498]), .A(ram[1434]), .S(n4284), .Y(n2964) );
  MUX2X1 U6437 ( .B(n2963), .A(n2960), .S(n4165), .Y(n2974) );
  MUX2X1 U6438 ( .B(ram[1626]), .A(ram[1562]), .S(n4284), .Y(n2968) );
  MUX2X1 U6439 ( .B(ram[1754]), .A(ram[1690]), .S(n4284), .Y(n2967) );
  MUX2X1 U6440 ( .B(ram[1882]), .A(ram[1818]), .S(n4284), .Y(n2971) );
  MUX2X1 U6441 ( .B(ram[2010]), .A(ram[1946]), .S(n4284), .Y(n2970) );
  MUX2X1 U6442 ( .B(n2969), .A(n2966), .S(n4165), .Y(n2973) );
  MUX2X1 U6443 ( .B(n2972), .A(n2957), .S(n4151), .Y(n4112) );
  MUX2X1 U6444 ( .B(ram[91]), .A(ram[27]), .S(n4284), .Y(n2977) );
  MUX2X1 U6445 ( .B(ram[219]), .A(ram[155]), .S(n4284), .Y(n2976) );
  MUX2X1 U6446 ( .B(ram[347]), .A(ram[283]), .S(n4284), .Y(n2980) );
  MUX2X1 U6447 ( .B(ram[475]), .A(ram[411]), .S(n4284), .Y(n2979) );
  MUX2X1 U6448 ( .B(n2978), .A(n2975), .S(n4165), .Y(n2990) );
  MUX2X1 U6449 ( .B(ram[603]), .A(ram[539]), .S(n4285), .Y(n2983) );
  MUX2X1 U6450 ( .B(ram[731]), .A(ram[667]), .S(n4285), .Y(n2982) );
  MUX2X1 U6451 ( .B(ram[859]), .A(ram[795]), .S(n4285), .Y(n2987) );
  MUX2X1 U6452 ( .B(ram[987]), .A(ram[923]), .S(n4285), .Y(n2985) );
  MUX2X1 U6453 ( .B(n2984), .A(n2981), .S(n4165), .Y(n2989) );
  MUX2X1 U6454 ( .B(ram[1115]), .A(ram[1051]), .S(n4285), .Y(n2993) );
  MUX2X1 U6455 ( .B(ram[1243]), .A(ram[1179]), .S(n4285), .Y(n2992) );
  MUX2X1 U6456 ( .B(ram[1371]), .A(ram[1307]), .S(n4285), .Y(n2996) );
  MUX2X1 U6457 ( .B(ram[1499]), .A(ram[1435]), .S(n4285), .Y(n2995) );
  MUX2X1 U6458 ( .B(n2994), .A(n2991), .S(n4165), .Y(n3005) );
  MUX2X1 U6459 ( .B(ram[1627]), .A(ram[1563]), .S(n4285), .Y(n2999) );
  MUX2X1 U6460 ( .B(ram[1755]), .A(ram[1691]), .S(n4285), .Y(n2998) );
  MUX2X1 U6461 ( .B(ram[1883]), .A(ram[1819]), .S(n4285), .Y(n3002) );
  MUX2X1 U6462 ( .B(ram[2011]), .A(ram[1947]), .S(n4285), .Y(n3001) );
  MUX2X1 U6463 ( .B(n3000), .A(n2997), .S(n4165), .Y(n3004) );
  MUX2X1 U6464 ( .B(n3003), .A(n2988), .S(n4150), .Y(n4113) );
  MUX2X1 U6465 ( .B(ram[92]), .A(ram[28]), .S(n4286), .Y(n3008) );
  MUX2X1 U6466 ( .B(ram[220]), .A(ram[156]), .S(n4286), .Y(n3007) );
  MUX2X1 U6467 ( .B(ram[348]), .A(ram[284]), .S(n4286), .Y(n3011) );
  MUX2X1 U6468 ( .B(ram[476]), .A(ram[412]), .S(n4286), .Y(n3010) );
  MUX2X1 U6469 ( .B(n3009), .A(n3006), .S(n4166), .Y(n3020) );
  MUX2X1 U6470 ( .B(ram[604]), .A(ram[540]), .S(n4286), .Y(n3014) );
  MUX2X1 U6471 ( .B(ram[732]), .A(ram[668]), .S(n4286), .Y(n3013) );
  MUX2X1 U6472 ( .B(ram[860]), .A(ram[796]), .S(n4286), .Y(n3017) );
  MUX2X1 U6473 ( .B(ram[988]), .A(ram[924]), .S(n4286), .Y(n3016) );
  MUX2X1 U6474 ( .B(n3015), .A(n3012), .S(n4166), .Y(n3019) );
  MUX2X1 U6475 ( .B(ram[1116]), .A(ram[1052]), .S(n4286), .Y(n3023) );
  MUX2X1 U6476 ( .B(ram[1244]), .A(ram[1180]), .S(n4286), .Y(n3022) );
  MUX2X1 U6477 ( .B(ram[1372]), .A(ram[1308]), .S(n4286), .Y(n3026) );
  MUX2X1 U6478 ( .B(ram[1500]), .A(ram[1436]), .S(n4286), .Y(n3025) );
  MUX2X1 U6479 ( .B(n3024), .A(n3021), .S(n4166), .Y(n3035) );
  MUX2X1 U6480 ( .B(ram[1628]), .A(ram[1564]), .S(n4287), .Y(n3029) );
  MUX2X1 U6481 ( .B(ram[1756]), .A(ram[1692]), .S(n4287), .Y(n3028) );
  MUX2X1 U6482 ( .B(ram[1884]), .A(ram[1820]), .S(n4287), .Y(n3032) );
  MUX2X1 U6483 ( .B(ram[2012]), .A(ram[1948]), .S(n4287), .Y(n3031) );
  MUX2X1 U6484 ( .B(n3030), .A(n3027), .S(n4166), .Y(n3034) );
  MUX2X1 U6485 ( .B(n3033), .A(n3018), .S(n4151), .Y(n4114) );
  MUX2X1 U6486 ( .B(ram[93]), .A(ram[29]), .S(n4287), .Y(n3038) );
  MUX2X1 U6487 ( .B(ram[221]), .A(ram[157]), .S(n4287), .Y(n3037) );
  MUX2X1 U6488 ( .B(ram[349]), .A(ram[285]), .S(n4287), .Y(n3041) );
  MUX2X1 U6489 ( .B(ram[477]), .A(ram[413]), .S(n4287), .Y(n3040) );
  MUX2X1 U6490 ( .B(n3039), .A(n3036), .S(n4166), .Y(n3050) );
  MUX2X1 U6491 ( .B(ram[605]), .A(ram[541]), .S(n4287), .Y(n3044) );
  MUX2X1 U6492 ( .B(ram[733]), .A(ram[669]), .S(n4287), .Y(n3043) );
  MUX2X1 U6493 ( .B(ram[861]), .A(ram[797]), .S(n4287), .Y(n3047) );
  MUX2X1 U6494 ( .B(ram[989]), .A(ram[925]), .S(n4287), .Y(n3046) );
  MUX2X1 U6495 ( .B(n3045), .A(n3042), .S(n4166), .Y(n3049) );
  MUX2X1 U6496 ( .B(ram[1117]), .A(ram[1053]), .S(n4288), .Y(n3053) );
  MUX2X1 U6497 ( .B(ram[1245]), .A(ram[1181]), .S(n4288), .Y(n3052) );
  MUX2X1 U6498 ( .B(ram[1373]), .A(ram[1309]), .S(n4288), .Y(n3056) );
  MUX2X1 U6499 ( .B(ram[1501]), .A(ram[1437]), .S(n4288), .Y(n3055) );
  MUX2X1 U6500 ( .B(n3054), .A(n3051), .S(n4166), .Y(n3065) );
  MUX2X1 U6501 ( .B(ram[1629]), .A(ram[1565]), .S(n4288), .Y(n3059) );
  MUX2X1 U6502 ( .B(ram[1757]), .A(ram[1693]), .S(n4288), .Y(n3058) );
  MUX2X1 U6503 ( .B(ram[1885]), .A(ram[1821]), .S(n4288), .Y(n3062) );
  MUX2X1 U6504 ( .B(ram[2013]), .A(ram[1949]), .S(n4288), .Y(n3061) );
  MUX2X1 U6505 ( .B(n3060), .A(n3057), .S(n4166), .Y(n3064) );
  MUX2X1 U6506 ( .B(n3063), .A(n3048), .S(n4152), .Y(n4115) );
  MUX2X1 U6507 ( .B(ram[94]), .A(ram[30]), .S(n4288), .Y(n3068) );
  MUX2X1 U6508 ( .B(ram[222]), .A(ram[158]), .S(n4288), .Y(n3067) );
  MUX2X1 U6509 ( .B(ram[350]), .A(ram[286]), .S(n4288), .Y(n3071) );
  MUX2X1 U6510 ( .B(ram[478]), .A(ram[414]), .S(n4288), .Y(n3070) );
  MUX2X1 U6511 ( .B(n3069), .A(n3066), .S(n4166), .Y(n3080) );
  MUX2X1 U6512 ( .B(ram[606]), .A(ram[542]), .S(n4289), .Y(n3074) );
  MUX2X1 U6513 ( .B(ram[734]), .A(ram[670]), .S(n4289), .Y(n3073) );
  MUX2X1 U6514 ( .B(ram[862]), .A(ram[798]), .S(n4289), .Y(n3077) );
  MUX2X1 U6515 ( .B(ram[990]), .A(ram[926]), .S(n4289), .Y(n3076) );
  MUX2X1 U6516 ( .B(n3075), .A(n3072), .S(n4166), .Y(n3079) );
  MUX2X1 U6517 ( .B(ram[1118]), .A(ram[1054]), .S(n4289), .Y(n3083) );
  MUX2X1 U6518 ( .B(ram[1246]), .A(ram[1182]), .S(n4289), .Y(n3082) );
  MUX2X1 U6519 ( .B(ram[1374]), .A(ram[1310]), .S(n4289), .Y(n3086) );
  MUX2X1 U6520 ( .B(ram[1502]), .A(ram[1438]), .S(n4289), .Y(n3085) );
  MUX2X1 U6521 ( .B(n3084), .A(n3081), .S(n4166), .Y(n3095) );
  MUX2X1 U6522 ( .B(ram[1630]), .A(ram[1566]), .S(n4289), .Y(n3089) );
  MUX2X1 U6523 ( .B(ram[1758]), .A(ram[1694]), .S(n4289), .Y(n3088) );
  MUX2X1 U6524 ( .B(ram[1886]), .A(ram[1822]), .S(n4289), .Y(n3092) );
  MUX2X1 U6525 ( .B(ram[2014]), .A(ram[1950]), .S(n4289), .Y(n3091) );
  MUX2X1 U6526 ( .B(n3090), .A(n3087), .S(n4166), .Y(n3094) );
  MUX2X1 U6527 ( .B(n3093), .A(n3078), .S(n4152), .Y(n4116) );
  MUX2X1 U6528 ( .B(ram[95]), .A(ram[31]), .S(n4290), .Y(n3098) );
  MUX2X1 U6529 ( .B(ram[223]), .A(ram[159]), .S(n4290), .Y(n3097) );
  MUX2X1 U6530 ( .B(ram[351]), .A(ram[287]), .S(n4290), .Y(n3101) );
  MUX2X1 U6531 ( .B(ram[479]), .A(ram[415]), .S(n4290), .Y(n3100) );
  MUX2X1 U6532 ( .B(n3099), .A(n3096), .S(n4167), .Y(n3110) );
  MUX2X1 U6533 ( .B(ram[607]), .A(ram[543]), .S(n4290), .Y(n3104) );
  MUX2X1 U6534 ( .B(ram[735]), .A(ram[671]), .S(n4290), .Y(n3103) );
  MUX2X1 U6535 ( .B(ram[863]), .A(ram[799]), .S(n4290), .Y(n3107) );
  MUX2X1 U6536 ( .B(ram[991]), .A(ram[927]), .S(n4290), .Y(n3106) );
  MUX2X1 U6537 ( .B(n3105), .A(n3102), .S(n4167), .Y(n3109) );
  MUX2X1 U6538 ( .B(ram[1119]), .A(ram[1055]), .S(n4290), .Y(n3113) );
  MUX2X1 U6539 ( .B(ram[1247]), .A(ram[1183]), .S(n4290), .Y(n3112) );
  MUX2X1 U6540 ( .B(ram[1375]), .A(ram[1311]), .S(n4290), .Y(n3116) );
  MUX2X1 U6541 ( .B(ram[1503]), .A(ram[1439]), .S(n4290), .Y(n3115) );
  MUX2X1 U6542 ( .B(n3114), .A(n3111), .S(n4167), .Y(n3125) );
  MUX2X1 U6543 ( .B(ram[1631]), .A(ram[1567]), .S(n4291), .Y(n3119) );
  MUX2X1 U6544 ( .B(ram[1759]), .A(ram[1695]), .S(n4291), .Y(n3118) );
  MUX2X1 U6545 ( .B(ram[1887]), .A(ram[1823]), .S(n4291), .Y(n3122) );
  MUX2X1 U6546 ( .B(ram[2015]), .A(ram[1951]), .S(n4291), .Y(n3121) );
  MUX2X1 U6547 ( .B(n3120), .A(n3117), .S(n4167), .Y(n3124) );
  MUX2X1 U6548 ( .B(n3123), .A(n3108), .S(n4150), .Y(n4117) );
  MUX2X1 U6549 ( .B(ram[96]), .A(ram[32]), .S(n4291), .Y(n3128) );
  MUX2X1 U6550 ( .B(ram[224]), .A(ram[160]), .S(n4291), .Y(n3127) );
  MUX2X1 U6551 ( .B(ram[352]), .A(ram[288]), .S(n4291), .Y(n3131) );
  MUX2X1 U6552 ( .B(ram[480]), .A(ram[416]), .S(n4291), .Y(n3130) );
  MUX2X1 U6553 ( .B(n3129), .A(n3126), .S(n4167), .Y(n3140) );
  MUX2X1 U6554 ( .B(ram[608]), .A(ram[544]), .S(n4291), .Y(n3134) );
  MUX2X1 U6555 ( .B(ram[736]), .A(ram[672]), .S(n4291), .Y(n3133) );
  MUX2X1 U6556 ( .B(ram[864]), .A(ram[800]), .S(n4291), .Y(n3137) );
  MUX2X1 U6557 ( .B(ram[992]), .A(ram[928]), .S(n4291), .Y(n3136) );
  MUX2X1 U6558 ( .B(n3135), .A(n3132), .S(n4167), .Y(n3139) );
  MUX2X1 U6559 ( .B(ram[1120]), .A(ram[1056]), .S(n4292), .Y(n3143) );
  MUX2X1 U6560 ( .B(ram[1248]), .A(ram[1184]), .S(n4292), .Y(n3142) );
  MUX2X1 U6561 ( .B(ram[1376]), .A(ram[1312]), .S(n4292), .Y(n3146) );
  MUX2X1 U6562 ( .B(ram[1504]), .A(ram[1440]), .S(n4292), .Y(n3145) );
  MUX2X1 U6563 ( .B(n3144), .A(n3141), .S(n4167), .Y(n3155) );
  MUX2X1 U6564 ( .B(ram[1632]), .A(ram[1568]), .S(n4292), .Y(n3149) );
  MUX2X1 U6565 ( .B(ram[1760]), .A(ram[1696]), .S(n4292), .Y(n3148) );
  MUX2X1 U6566 ( .B(ram[1888]), .A(ram[1824]), .S(n4292), .Y(n3152) );
  MUX2X1 U6567 ( .B(ram[2016]), .A(ram[1952]), .S(n4292), .Y(n3151) );
  MUX2X1 U6568 ( .B(n3150), .A(n3147), .S(n4167), .Y(n3154) );
  MUX2X1 U6569 ( .B(n3153), .A(n3138), .S(n4150), .Y(n4118) );
  MUX2X1 U6570 ( .B(ram[97]), .A(ram[33]), .S(n4292), .Y(n3158) );
  MUX2X1 U6571 ( .B(ram[225]), .A(ram[161]), .S(n4292), .Y(n3157) );
  MUX2X1 U6572 ( .B(ram[353]), .A(ram[289]), .S(n4292), .Y(n3161) );
  MUX2X1 U6573 ( .B(ram[481]), .A(ram[417]), .S(n4292), .Y(n3160) );
  MUX2X1 U6574 ( .B(n3159), .A(n3156), .S(n4167), .Y(n3170) );
  MUX2X1 U6575 ( .B(ram[609]), .A(ram[545]), .S(n4293), .Y(n3164) );
  MUX2X1 U6576 ( .B(ram[737]), .A(ram[673]), .S(n4293), .Y(n3163) );
  MUX2X1 U6577 ( .B(ram[865]), .A(ram[801]), .S(n4293), .Y(n3167) );
  MUX2X1 U6578 ( .B(ram[993]), .A(ram[929]), .S(n4293), .Y(n3166) );
  MUX2X1 U6579 ( .B(n3165), .A(n3162), .S(n4167), .Y(n3169) );
  MUX2X1 U6580 ( .B(ram[1121]), .A(ram[1057]), .S(n4293), .Y(n3173) );
  MUX2X1 U6581 ( .B(ram[1249]), .A(ram[1185]), .S(n4293), .Y(n3172) );
  MUX2X1 U6582 ( .B(ram[1377]), .A(ram[1313]), .S(n4293), .Y(n3176) );
  MUX2X1 U6583 ( .B(ram[1505]), .A(ram[1441]), .S(n4293), .Y(n3175) );
  MUX2X1 U6584 ( .B(n3174), .A(n3171), .S(n4167), .Y(n3185) );
  MUX2X1 U6585 ( .B(ram[1633]), .A(ram[1569]), .S(n4293), .Y(n3179) );
  MUX2X1 U6586 ( .B(ram[1761]), .A(ram[1697]), .S(n4293), .Y(n3178) );
  MUX2X1 U6587 ( .B(ram[1889]), .A(ram[1825]), .S(n4293), .Y(n3182) );
  MUX2X1 U6588 ( .B(ram[2017]), .A(ram[1953]), .S(n4293), .Y(n3181) );
  MUX2X1 U6589 ( .B(n3180), .A(n3177), .S(n4167), .Y(n3184) );
  MUX2X1 U6590 ( .B(n3183), .A(n3168), .S(n4151), .Y(n4119) );
  MUX2X1 U6591 ( .B(ram[98]), .A(ram[34]), .S(n4294), .Y(n3188) );
  MUX2X1 U6592 ( .B(ram[226]), .A(ram[162]), .S(n4294), .Y(n3187) );
  MUX2X1 U6593 ( .B(ram[354]), .A(ram[290]), .S(n4294), .Y(n3191) );
  MUX2X1 U6594 ( .B(ram[482]), .A(ram[418]), .S(n4294), .Y(n3190) );
  MUX2X1 U6595 ( .B(n3189), .A(n3186), .S(n4168), .Y(n3200) );
  MUX2X1 U6596 ( .B(ram[610]), .A(ram[546]), .S(n4294), .Y(n3194) );
  MUX2X1 U6597 ( .B(ram[738]), .A(ram[674]), .S(n4294), .Y(n3193) );
  MUX2X1 U6598 ( .B(ram[866]), .A(ram[802]), .S(n4294), .Y(n3197) );
  MUX2X1 U6599 ( .B(ram[994]), .A(ram[930]), .S(n4294), .Y(n3196) );
  MUX2X1 U6600 ( .B(n3195), .A(n3192), .S(n4168), .Y(n3199) );
  MUX2X1 U6601 ( .B(ram[1122]), .A(ram[1058]), .S(n4294), .Y(n3203) );
  MUX2X1 U6602 ( .B(ram[1250]), .A(ram[1186]), .S(n4294), .Y(n3202) );
  MUX2X1 U6603 ( .B(ram[1378]), .A(ram[1314]), .S(n4294), .Y(n3206) );
  MUX2X1 U6604 ( .B(ram[1506]), .A(ram[1442]), .S(n4294), .Y(n3205) );
  MUX2X1 U6605 ( .B(n3204), .A(n3201), .S(n4168), .Y(n3215) );
  MUX2X1 U6606 ( .B(ram[1634]), .A(ram[1570]), .S(n4295), .Y(n3209) );
  MUX2X1 U6607 ( .B(ram[1762]), .A(ram[1698]), .S(n4295), .Y(n3208) );
  MUX2X1 U6608 ( .B(ram[1890]), .A(ram[1826]), .S(n4295), .Y(n3212) );
  MUX2X1 U6609 ( .B(ram[2018]), .A(ram[1954]), .S(n4295), .Y(n3211) );
  MUX2X1 U6610 ( .B(n3210), .A(n3207), .S(n4168), .Y(n3214) );
  MUX2X1 U6611 ( .B(n3213), .A(n3198), .S(n4152), .Y(n4120) );
  MUX2X1 U6612 ( .B(ram[99]), .A(ram[35]), .S(n4295), .Y(n3218) );
  MUX2X1 U6613 ( .B(ram[227]), .A(ram[163]), .S(n4295), .Y(n3217) );
  MUX2X1 U6614 ( .B(ram[355]), .A(ram[291]), .S(n4295), .Y(n3221) );
  MUX2X1 U6615 ( .B(ram[483]), .A(ram[419]), .S(n4295), .Y(n3220) );
  MUX2X1 U6616 ( .B(n3219), .A(n3216), .S(n4168), .Y(n3230) );
  MUX2X1 U6617 ( .B(ram[611]), .A(ram[547]), .S(n4295), .Y(n3224) );
  MUX2X1 U6618 ( .B(ram[739]), .A(ram[675]), .S(n4295), .Y(n3223) );
  MUX2X1 U6619 ( .B(ram[867]), .A(ram[803]), .S(n4295), .Y(n3227) );
  MUX2X1 U6620 ( .B(ram[995]), .A(ram[931]), .S(n4295), .Y(n3226) );
  MUX2X1 U6621 ( .B(n3225), .A(n3222), .S(n4168), .Y(n3229) );
  MUX2X1 U6622 ( .B(ram[1123]), .A(ram[1059]), .S(n4296), .Y(n3233) );
  MUX2X1 U6623 ( .B(ram[1251]), .A(ram[1187]), .S(n4296), .Y(n3232) );
  MUX2X1 U6624 ( .B(ram[1379]), .A(ram[1315]), .S(n4296), .Y(n3236) );
  MUX2X1 U6625 ( .B(ram[1507]), .A(ram[1443]), .S(n4296), .Y(n3235) );
  MUX2X1 U6626 ( .B(n3234), .A(n3231), .S(n4168), .Y(n3245) );
  MUX2X1 U6627 ( .B(ram[1635]), .A(ram[1571]), .S(n4296), .Y(n3239) );
  MUX2X1 U6628 ( .B(ram[1763]), .A(ram[1699]), .S(n4296), .Y(n3238) );
  MUX2X1 U6629 ( .B(ram[1891]), .A(ram[1827]), .S(n4296), .Y(n3242) );
  MUX2X1 U6630 ( .B(ram[2019]), .A(ram[1955]), .S(n4296), .Y(n3241) );
  MUX2X1 U6631 ( .B(n3240), .A(n3237), .S(n4168), .Y(n3244) );
  MUX2X1 U6632 ( .B(n3243), .A(n3228), .S(n4151), .Y(n4121) );
  MUX2X1 U6633 ( .B(ram[100]), .A(ram[36]), .S(n4296), .Y(n3248) );
  MUX2X1 U6634 ( .B(ram[228]), .A(ram[164]), .S(n4296), .Y(n3247) );
  MUX2X1 U6635 ( .B(ram[356]), .A(ram[292]), .S(n4296), .Y(n3251) );
  MUX2X1 U6636 ( .B(ram[484]), .A(ram[420]), .S(n4296), .Y(n3250) );
  MUX2X1 U6637 ( .B(n3249), .A(n3246), .S(n4168), .Y(n3260) );
  MUX2X1 U6638 ( .B(ram[612]), .A(ram[548]), .S(n4297), .Y(n3254) );
  MUX2X1 U6639 ( .B(ram[740]), .A(ram[676]), .S(n4297), .Y(n3253) );
  MUX2X1 U6640 ( .B(ram[868]), .A(ram[804]), .S(n4297), .Y(n3257) );
  MUX2X1 U6641 ( .B(ram[996]), .A(ram[932]), .S(n4297), .Y(n3256) );
  MUX2X1 U6642 ( .B(n3255), .A(n3252), .S(n4168), .Y(n3259) );
  MUX2X1 U6643 ( .B(ram[1124]), .A(ram[1060]), .S(n4297), .Y(n3263) );
  MUX2X1 U6644 ( .B(ram[1252]), .A(ram[1188]), .S(n4297), .Y(n3262) );
  MUX2X1 U6645 ( .B(ram[1380]), .A(ram[1316]), .S(n4297), .Y(n3266) );
  MUX2X1 U6646 ( .B(ram[1508]), .A(ram[1444]), .S(n4297), .Y(n3265) );
  MUX2X1 U6647 ( .B(n3264), .A(n3261), .S(n4168), .Y(n3275) );
  MUX2X1 U6648 ( .B(ram[1636]), .A(ram[1572]), .S(n4297), .Y(n3269) );
  MUX2X1 U6649 ( .B(ram[1764]), .A(ram[1700]), .S(n4297), .Y(n3268) );
  MUX2X1 U6650 ( .B(ram[1892]), .A(ram[1828]), .S(n4297), .Y(n3272) );
  MUX2X1 U6651 ( .B(ram[2020]), .A(ram[1956]), .S(n4297), .Y(n3271) );
  MUX2X1 U6652 ( .B(n3270), .A(n3267), .S(n4168), .Y(n3274) );
  MUX2X1 U6653 ( .B(n3273), .A(n3258), .S(n4151), .Y(n4122) );
  MUX2X1 U6654 ( .B(ram[101]), .A(ram[37]), .S(n4298), .Y(n3278) );
  MUX2X1 U6655 ( .B(ram[229]), .A(ram[165]), .S(n4298), .Y(n3277) );
  MUX2X1 U6656 ( .B(ram[357]), .A(ram[293]), .S(n4298), .Y(n3281) );
  MUX2X1 U6657 ( .B(ram[485]), .A(ram[421]), .S(n4298), .Y(n3280) );
  MUX2X1 U6658 ( .B(n3279), .A(n3276), .S(n4169), .Y(n3290) );
  MUX2X1 U6659 ( .B(ram[613]), .A(ram[549]), .S(n4298), .Y(n3284) );
  MUX2X1 U6660 ( .B(ram[741]), .A(ram[677]), .S(n4298), .Y(n3283) );
  MUX2X1 U6661 ( .B(ram[869]), .A(ram[805]), .S(n4298), .Y(n3287) );
  MUX2X1 U6662 ( .B(ram[997]), .A(ram[933]), .S(n4298), .Y(n3286) );
  MUX2X1 U6663 ( .B(n3285), .A(n3282), .S(n4169), .Y(n3289) );
  MUX2X1 U6664 ( .B(ram[1125]), .A(ram[1061]), .S(n4298), .Y(n3293) );
  MUX2X1 U6665 ( .B(ram[1253]), .A(ram[1189]), .S(n4298), .Y(n3292) );
  MUX2X1 U6666 ( .B(ram[1381]), .A(ram[1317]), .S(n4298), .Y(n3296) );
  MUX2X1 U6667 ( .B(ram[1509]), .A(ram[1445]), .S(n4298), .Y(n3295) );
  MUX2X1 U6668 ( .B(n3294), .A(n3291), .S(n4169), .Y(n3305) );
  MUX2X1 U6669 ( .B(ram[1637]), .A(ram[1573]), .S(n4299), .Y(n3299) );
  MUX2X1 U6670 ( .B(ram[1765]), .A(ram[1701]), .S(n4299), .Y(n3298) );
  MUX2X1 U6671 ( .B(ram[1893]), .A(ram[1829]), .S(n4299), .Y(n3302) );
  MUX2X1 U6672 ( .B(ram[2021]), .A(ram[1957]), .S(n4299), .Y(n3301) );
  MUX2X1 U6673 ( .B(n3300), .A(n3297), .S(n4169), .Y(n3304) );
  MUX2X1 U6674 ( .B(n3303), .A(n3288), .S(n4151), .Y(n4123) );
  MUX2X1 U6675 ( .B(ram[102]), .A(ram[38]), .S(n4299), .Y(n3308) );
  MUX2X1 U6676 ( .B(ram[230]), .A(ram[166]), .S(n4299), .Y(n3307) );
  MUX2X1 U6677 ( .B(ram[358]), .A(ram[294]), .S(n4299), .Y(n3311) );
  MUX2X1 U6678 ( .B(ram[486]), .A(ram[422]), .S(n4299), .Y(n3310) );
  MUX2X1 U6679 ( .B(n3309), .A(n3306), .S(n4169), .Y(n3320) );
  MUX2X1 U6680 ( .B(ram[614]), .A(ram[550]), .S(n4299), .Y(n3314) );
  MUX2X1 U6681 ( .B(ram[742]), .A(ram[678]), .S(n4299), .Y(n3313) );
  MUX2X1 U6682 ( .B(ram[870]), .A(ram[806]), .S(n4299), .Y(n3317) );
  MUX2X1 U6683 ( .B(ram[998]), .A(ram[934]), .S(n4299), .Y(n3316) );
  MUX2X1 U6684 ( .B(n3315), .A(n3312), .S(n4169), .Y(n3319) );
  MUX2X1 U6685 ( .B(ram[1126]), .A(ram[1062]), .S(n4300), .Y(n3323) );
  MUX2X1 U6686 ( .B(ram[1254]), .A(ram[1190]), .S(n4300), .Y(n3322) );
  MUX2X1 U6687 ( .B(ram[1382]), .A(ram[1318]), .S(n4300), .Y(n3326) );
  MUX2X1 U6688 ( .B(ram[1510]), .A(ram[1446]), .S(n4300), .Y(n3325) );
  MUX2X1 U6689 ( .B(n3324), .A(n3321), .S(n4169), .Y(n3335) );
  MUX2X1 U6690 ( .B(ram[1638]), .A(ram[1574]), .S(n4300), .Y(n3329) );
  MUX2X1 U6691 ( .B(ram[1766]), .A(ram[1702]), .S(n4300), .Y(n3328) );
  MUX2X1 U6692 ( .B(ram[1894]), .A(ram[1830]), .S(n4300), .Y(n3332) );
  MUX2X1 U6693 ( .B(ram[2022]), .A(ram[1958]), .S(n4300), .Y(n3331) );
  MUX2X1 U6694 ( .B(n3330), .A(n3327), .S(n4169), .Y(n3334) );
  MUX2X1 U6695 ( .B(n3333), .A(n3318), .S(n4151), .Y(n4124) );
  MUX2X1 U6696 ( .B(ram[103]), .A(ram[39]), .S(n4300), .Y(n3338) );
  MUX2X1 U6697 ( .B(ram[231]), .A(ram[167]), .S(n4300), .Y(n3337) );
  MUX2X1 U6698 ( .B(ram[359]), .A(ram[295]), .S(n4300), .Y(n3341) );
  MUX2X1 U6699 ( .B(ram[487]), .A(ram[423]), .S(n4300), .Y(n3340) );
  MUX2X1 U6700 ( .B(n3339), .A(n3336), .S(n4169), .Y(n3350) );
  MUX2X1 U6701 ( .B(ram[615]), .A(ram[551]), .S(n4301), .Y(n3344) );
  MUX2X1 U6702 ( .B(ram[743]), .A(ram[679]), .S(n4301), .Y(n3343) );
  MUX2X1 U6703 ( .B(ram[871]), .A(ram[807]), .S(n4301), .Y(n3347) );
  MUX2X1 U6704 ( .B(ram[999]), .A(ram[935]), .S(n4301), .Y(n3346) );
  MUX2X1 U6705 ( .B(n3345), .A(n3342), .S(n4169), .Y(n3349) );
  MUX2X1 U6706 ( .B(ram[1127]), .A(ram[1063]), .S(n4301), .Y(n3353) );
  MUX2X1 U6707 ( .B(ram[1255]), .A(ram[1191]), .S(n4301), .Y(n3352) );
  MUX2X1 U6708 ( .B(ram[1383]), .A(ram[1319]), .S(n4301), .Y(n3356) );
  MUX2X1 U6709 ( .B(ram[1511]), .A(ram[1447]), .S(n4301), .Y(n3355) );
  MUX2X1 U6710 ( .B(n3354), .A(n3351), .S(n4169), .Y(n3365) );
  MUX2X1 U6711 ( .B(ram[1639]), .A(ram[1575]), .S(n4301), .Y(n3359) );
  MUX2X1 U6712 ( .B(ram[1767]), .A(ram[1703]), .S(n4301), .Y(n3358) );
  MUX2X1 U6713 ( .B(ram[1895]), .A(ram[1831]), .S(n4301), .Y(n3362) );
  MUX2X1 U6714 ( .B(ram[2023]), .A(ram[1959]), .S(n4301), .Y(n3361) );
  MUX2X1 U6715 ( .B(n3360), .A(n3357), .S(n4169), .Y(n3364) );
  MUX2X1 U6716 ( .B(n3363), .A(n3348), .S(n4151), .Y(n4125) );
  MUX2X1 U6717 ( .B(ram[104]), .A(ram[40]), .S(n4302), .Y(n3368) );
  MUX2X1 U6718 ( .B(ram[232]), .A(ram[168]), .S(n4302), .Y(n3367) );
  MUX2X1 U6719 ( .B(ram[360]), .A(ram[296]), .S(n4302), .Y(n3371) );
  MUX2X1 U6720 ( .B(ram[488]), .A(ram[424]), .S(n4302), .Y(n3370) );
  MUX2X1 U6721 ( .B(n3369), .A(n3366), .S(n4170), .Y(n3380) );
  MUX2X1 U6722 ( .B(ram[616]), .A(ram[552]), .S(n4302), .Y(n3374) );
  MUX2X1 U6723 ( .B(ram[744]), .A(ram[680]), .S(n4302), .Y(n3373) );
  MUX2X1 U6724 ( .B(ram[872]), .A(ram[808]), .S(n4302), .Y(n3377) );
  MUX2X1 U6725 ( .B(ram[1000]), .A(ram[936]), .S(n4302), .Y(n3376) );
  MUX2X1 U6726 ( .B(n3375), .A(n3372), .S(n4170), .Y(n3379) );
  MUX2X1 U6727 ( .B(ram[1128]), .A(ram[1064]), .S(n4302), .Y(n3383) );
  MUX2X1 U6728 ( .B(ram[1256]), .A(ram[1192]), .S(n4302), .Y(n3382) );
  MUX2X1 U6729 ( .B(ram[1384]), .A(ram[1320]), .S(n4302), .Y(n3386) );
  MUX2X1 U6730 ( .B(ram[1512]), .A(ram[1448]), .S(n4302), .Y(n3385) );
  MUX2X1 U6731 ( .B(n3384), .A(n3381), .S(n4170), .Y(n3395) );
  MUX2X1 U6732 ( .B(ram[1640]), .A(ram[1576]), .S(n4303), .Y(n3389) );
  MUX2X1 U6733 ( .B(ram[1768]), .A(ram[1704]), .S(n4303), .Y(n3388) );
  MUX2X1 U6734 ( .B(ram[1896]), .A(ram[1832]), .S(n4303), .Y(n3392) );
  MUX2X1 U6735 ( .B(ram[2024]), .A(ram[1960]), .S(n4303), .Y(n3391) );
  MUX2X1 U6736 ( .B(n3390), .A(n3387), .S(n4170), .Y(n3394) );
  MUX2X1 U6737 ( .B(n3393), .A(n3378), .S(n4151), .Y(n4126) );
  MUX2X1 U6738 ( .B(ram[105]), .A(ram[41]), .S(n4303), .Y(n3398) );
  MUX2X1 U6739 ( .B(ram[233]), .A(ram[169]), .S(n4303), .Y(n3397) );
  MUX2X1 U6740 ( .B(ram[361]), .A(ram[297]), .S(n4303), .Y(n3401) );
  MUX2X1 U6741 ( .B(ram[489]), .A(ram[425]), .S(n4303), .Y(n3400) );
  MUX2X1 U6742 ( .B(n3399), .A(n3396), .S(n4170), .Y(n3410) );
  MUX2X1 U6743 ( .B(ram[617]), .A(ram[553]), .S(n4303), .Y(n3404) );
  MUX2X1 U6744 ( .B(ram[745]), .A(ram[681]), .S(n4303), .Y(n3403) );
  MUX2X1 U6745 ( .B(ram[873]), .A(ram[809]), .S(n4303), .Y(n3407) );
  MUX2X1 U6746 ( .B(ram[1001]), .A(ram[937]), .S(n4303), .Y(n3406) );
  MUX2X1 U6747 ( .B(n3405), .A(n3402), .S(n4170), .Y(n3409) );
  MUX2X1 U6748 ( .B(ram[1129]), .A(ram[1065]), .S(n4304), .Y(n3413) );
  MUX2X1 U6749 ( .B(ram[1257]), .A(ram[1193]), .S(n4304), .Y(n3412) );
  MUX2X1 U6750 ( .B(ram[1385]), .A(ram[1321]), .S(n4304), .Y(n3416) );
  MUX2X1 U6751 ( .B(ram[1513]), .A(ram[1449]), .S(n4304), .Y(n3415) );
  MUX2X1 U6752 ( .B(n3414), .A(n3411), .S(n4170), .Y(n3425) );
  MUX2X1 U6753 ( .B(ram[1641]), .A(ram[1577]), .S(n4304), .Y(n3419) );
  MUX2X1 U6754 ( .B(ram[1769]), .A(ram[1705]), .S(n4304), .Y(n3418) );
  MUX2X1 U6755 ( .B(ram[1897]), .A(ram[1833]), .S(n4304), .Y(n3422) );
  MUX2X1 U6756 ( .B(ram[2025]), .A(ram[1961]), .S(n4304), .Y(n3421) );
  MUX2X1 U6757 ( .B(n3420), .A(n3417), .S(n4170), .Y(n3424) );
  MUX2X1 U6758 ( .B(n3423), .A(n3408), .S(n4151), .Y(n4127) );
  MUX2X1 U6759 ( .B(ram[106]), .A(ram[42]), .S(n4304), .Y(n3428) );
  MUX2X1 U6760 ( .B(ram[234]), .A(ram[170]), .S(n4304), .Y(n3427) );
  MUX2X1 U6761 ( .B(ram[362]), .A(ram[298]), .S(n4304), .Y(n3431) );
  MUX2X1 U6762 ( .B(ram[490]), .A(ram[426]), .S(n4304), .Y(n3430) );
  MUX2X1 U6763 ( .B(n3429), .A(n3426), .S(n4170), .Y(n3440) );
  MUX2X1 U6764 ( .B(ram[618]), .A(ram[554]), .S(n4305), .Y(n3434) );
  MUX2X1 U6765 ( .B(ram[746]), .A(ram[682]), .S(n4305), .Y(n3433) );
  MUX2X1 U6766 ( .B(ram[874]), .A(ram[810]), .S(n4305), .Y(n3437) );
  MUX2X1 U6767 ( .B(ram[1002]), .A(ram[938]), .S(n4305), .Y(n3436) );
  MUX2X1 U6768 ( .B(n3435), .A(n3432), .S(n4170), .Y(n3439) );
  MUX2X1 U6769 ( .B(ram[1130]), .A(ram[1066]), .S(n4305), .Y(n3443) );
  MUX2X1 U6770 ( .B(ram[1258]), .A(ram[1194]), .S(n4305), .Y(n3442) );
  MUX2X1 U6771 ( .B(ram[1386]), .A(ram[1322]), .S(n4305), .Y(n3446) );
  MUX2X1 U6772 ( .B(ram[1514]), .A(ram[1450]), .S(n4305), .Y(n3445) );
  MUX2X1 U6773 ( .B(n3444), .A(n3441), .S(n4170), .Y(n3455) );
  MUX2X1 U6774 ( .B(ram[1642]), .A(ram[1578]), .S(n4305), .Y(n3449) );
  MUX2X1 U6775 ( .B(ram[1770]), .A(ram[1706]), .S(n4305), .Y(n3448) );
  MUX2X1 U6776 ( .B(ram[1898]), .A(ram[1834]), .S(n4305), .Y(n3452) );
  MUX2X1 U6777 ( .B(ram[2026]), .A(ram[1962]), .S(n4305), .Y(n3451) );
  MUX2X1 U6778 ( .B(n3450), .A(n3447), .S(n4170), .Y(n3454) );
  MUX2X1 U6779 ( .B(n3453), .A(n3438), .S(n4151), .Y(n4128) );
  MUX2X1 U6780 ( .B(ram[107]), .A(ram[43]), .S(n4305), .Y(n3458) );
  MUX2X1 U6781 ( .B(ram[235]), .A(ram[171]), .S(n4269), .Y(n3457) );
  MUX2X1 U6782 ( .B(ram[363]), .A(ram[299]), .S(n4306), .Y(n3461) );
  MUX2X1 U6783 ( .B(ram[491]), .A(ram[427]), .S(n4300), .Y(n3460) );
  MUX2X1 U6784 ( .B(n3459), .A(n3456), .S(n4171), .Y(n3470) );
  MUX2X1 U6785 ( .B(ram[619]), .A(ram[555]), .S(n4301), .Y(n3464) );
  MUX2X1 U6786 ( .B(ram[747]), .A(ram[683]), .S(n4328), .Y(n3463) );
  MUX2X1 U6787 ( .B(ram[875]), .A(ram[811]), .S(n4326), .Y(n3467) );
  MUX2X1 U6788 ( .B(ram[1003]), .A(ram[939]), .S(n4295), .Y(n3466) );
  MUX2X1 U6789 ( .B(n3465), .A(n3462), .S(n4171), .Y(n3469) );
  MUX2X1 U6790 ( .B(ram[1131]), .A(ram[1067]), .S(n4290), .Y(n3473) );
  MUX2X1 U6791 ( .B(ram[1259]), .A(ram[1195]), .S(n4268), .Y(n3472) );
  MUX2X1 U6792 ( .B(ram[1387]), .A(ram[1323]), .S(n4306), .Y(n3476) );
  MUX2X1 U6793 ( .B(ram[1515]), .A(ram[1451]), .S(n4298), .Y(n3475) );
  MUX2X1 U6794 ( .B(n3474), .A(n3471), .S(n4171), .Y(n3485) );
  MUX2X1 U6795 ( .B(ram[1643]), .A(ram[1579]), .S(n4306), .Y(n3479) );
  MUX2X1 U6796 ( .B(ram[1771]), .A(ram[1707]), .S(n4306), .Y(n3478) );
  MUX2X1 U6797 ( .B(ram[1899]), .A(ram[1835]), .S(n4306), .Y(n3482) );
  MUX2X1 U6798 ( .B(ram[2027]), .A(ram[1963]), .S(n4306), .Y(n3481) );
  MUX2X1 U6799 ( .B(n3480), .A(n3477), .S(n4171), .Y(n3484) );
  MUX2X1 U6800 ( .B(n3483), .A(n3468), .S(n4151), .Y(n4129) );
  MUX2X1 U6801 ( .B(ram[108]), .A(ram[44]), .S(n4306), .Y(n3488) );
  MUX2X1 U6802 ( .B(ram[236]), .A(ram[172]), .S(n4306), .Y(n3487) );
  MUX2X1 U6803 ( .B(ram[364]), .A(ram[300]), .S(n4306), .Y(n3491) );
  MUX2X1 U6804 ( .B(ram[492]), .A(ram[428]), .S(n4306), .Y(n3490) );
  MUX2X1 U6805 ( .B(n3489), .A(n3486), .S(n4171), .Y(n3500) );
  MUX2X1 U6806 ( .B(ram[620]), .A(ram[556]), .S(n4306), .Y(n3494) );
  MUX2X1 U6807 ( .B(ram[748]), .A(ram[684]), .S(n4306), .Y(n3493) );
  MUX2X1 U6808 ( .B(ram[876]), .A(ram[812]), .S(n4306), .Y(n3497) );
  MUX2X1 U6809 ( .B(ram[1004]), .A(ram[940]), .S(n4306), .Y(n3496) );
  MUX2X1 U6810 ( .B(n3495), .A(n3492), .S(n4171), .Y(n3499) );
  MUX2X1 U6811 ( .B(ram[1132]), .A(ram[1068]), .S(n4307), .Y(n3503) );
  MUX2X1 U6812 ( .B(ram[1260]), .A(ram[1196]), .S(n4307), .Y(n3502) );
  MUX2X1 U6813 ( .B(ram[1388]), .A(ram[1324]), .S(n4307), .Y(n3506) );
  MUX2X1 U6814 ( .B(ram[1516]), .A(ram[1452]), .S(n4307), .Y(n3505) );
  MUX2X1 U6815 ( .B(n3504), .A(n3501), .S(n4171), .Y(n3515) );
  MUX2X1 U6816 ( .B(ram[1644]), .A(ram[1580]), .S(n4307), .Y(n3509) );
  MUX2X1 U6817 ( .B(ram[1772]), .A(ram[1708]), .S(n4307), .Y(n3508) );
  MUX2X1 U6818 ( .B(ram[1900]), .A(ram[1836]), .S(n4307), .Y(n3512) );
  MUX2X1 U6819 ( .B(ram[2028]), .A(ram[1964]), .S(n4307), .Y(n3511) );
  MUX2X1 U6820 ( .B(n3510), .A(n3507), .S(n4171), .Y(n3514) );
  MUX2X1 U6821 ( .B(n3513), .A(n3498), .S(n4151), .Y(n4130) );
  MUX2X1 U6822 ( .B(ram[109]), .A(ram[45]), .S(n4307), .Y(n3518) );
  MUX2X1 U6823 ( .B(ram[237]), .A(ram[173]), .S(n4307), .Y(n3517) );
  MUX2X1 U6824 ( .B(ram[365]), .A(ram[301]), .S(n4307), .Y(n3521) );
  MUX2X1 U6825 ( .B(ram[493]), .A(ram[429]), .S(n4307), .Y(n3520) );
  MUX2X1 U6826 ( .B(n3519), .A(n3516), .S(n4171), .Y(n3530) );
  MUX2X1 U6827 ( .B(ram[621]), .A(ram[557]), .S(n4308), .Y(n3524) );
  MUX2X1 U6828 ( .B(ram[749]), .A(ram[685]), .S(n4308), .Y(n3523) );
  MUX2X1 U6829 ( .B(ram[877]), .A(ram[813]), .S(n4308), .Y(n3527) );
  MUX2X1 U6830 ( .B(ram[1005]), .A(ram[941]), .S(n4308), .Y(n3526) );
  MUX2X1 U6831 ( .B(n3525), .A(n3522), .S(n4171), .Y(n3529) );
  MUX2X1 U6832 ( .B(ram[1133]), .A(ram[1069]), .S(n4308), .Y(n3533) );
  MUX2X1 U6833 ( .B(ram[1261]), .A(ram[1197]), .S(n4308), .Y(n3532) );
  MUX2X1 U6834 ( .B(ram[1389]), .A(ram[1325]), .S(n4308), .Y(n3536) );
  MUX2X1 U6835 ( .B(ram[1517]), .A(ram[1453]), .S(n4308), .Y(n3535) );
  MUX2X1 U6836 ( .B(n3534), .A(n3531), .S(n4171), .Y(n3545) );
  MUX2X1 U6837 ( .B(ram[1645]), .A(ram[1581]), .S(n4308), .Y(n3539) );
  MUX2X1 U6838 ( .B(ram[1773]), .A(ram[1709]), .S(n4308), .Y(n3538) );
  MUX2X1 U6839 ( .B(ram[1901]), .A(ram[1837]), .S(n4308), .Y(n3542) );
  MUX2X1 U6840 ( .B(ram[2029]), .A(ram[1965]), .S(n4308), .Y(n3541) );
  MUX2X1 U6841 ( .B(n3540), .A(n3537), .S(n4171), .Y(n3544) );
  MUX2X1 U6842 ( .B(n3543), .A(n3528), .S(n4151), .Y(n4131) );
  MUX2X1 U6843 ( .B(ram[110]), .A(ram[46]), .S(n4305), .Y(n3548) );
  MUX2X1 U6844 ( .B(ram[238]), .A(ram[174]), .S(n4323), .Y(n3547) );
  MUX2X1 U6845 ( .B(ram[366]), .A(ram[302]), .S(n4305), .Y(n3551) );
  MUX2X1 U6846 ( .B(ram[494]), .A(ram[430]), .S(n4309), .Y(n3550) );
  MUX2X1 U6847 ( .B(n3549), .A(n3546), .S(n4172), .Y(n3560) );
  MUX2X1 U6848 ( .B(ram[622]), .A(ram[558]), .S(n4315), .Y(n3554) );
  MUX2X1 U6849 ( .B(ram[750]), .A(ram[686]), .S(n4318), .Y(n3553) );
  MUX2X1 U6850 ( .B(ram[878]), .A(ram[814]), .S(n4328), .Y(n3557) );
  MUX2X1 U6851 ( .B(ram[1006]), .A(ram[942]), .S(n4329), .Y(n3556) );
  MUX2X1 U6852 ( .B(n3555), .A(n3552), .S(n4172), .Y(n3559) );
  MUX2X1 U6853 ( .B(ram[1134]), .A(ram[1070]), .S(n4329), .Y(n3563) );
  MUX2X1 U6854 ( .B(ram[1262]), .A(ram[1198]), .S(n4323), .Y(n3562) );
  MUX2X1 U6855 ( .B(ram[1390]), .A(ram[1326]), .S(n4309), .Y(n3566) );
  MUX2X1 U6856 ( .B(ram[1518]), .A(ram[1454]), .S(n4328), .Y(n3565) );
  MUX2X1 U6857 ( .B(n3564), .A(n3561), .S(n4172), .Y(n3575) );
  MUX2X1 U6858 ( .B(ram[1646]), .A(ram[1582]), .S(n4309), .Y(n3569) );
  MUX2X1 U6859 ( .B(ram[1774]), .A(ram[1710]), .S(n4309), .Y(n3568) );
  MUX2X1 U6860 ( .B(ram[1902]), .A(ram[1838]), .S(n4309), .Y(n3572) );
  MUX2X1 U6861 ( .B(ram[2030]), .A(ram[1966]), .S(n4309), .Y(n3571) );
  MUX2X1 U6862 ( .B(n3570), .A(n3567), .S(n4172), .Y(n3574) );
  MUX2X1 U6863 ( .B(n3573), .A(n3558), .S(n4151), .Y(n4132) );
  MUX2X1 U6864 ( .B(ram[111]), .A(ram[47]), .S(n4309), .Y(n3578) );
  MUX2X1 U6865 ( .B(ram[239]), .A(ram[175]), .S(n4309), .Y(n3577) );
  MUX2X1 U6866 ( .B(ram[367]), .A(ram[303]), .S(n4309), .Y(n3581) );
  MUX2X1 U6867 ( .B(ram[495]), .A(ram[431]), .S(n4309), .Y(n3580) );
  MUX2X1 U6868 ( .B(n3579), .A(n3576), .S(n4172), .Y(n3590) );
  MUX2X1 U6869 ( .B(ram[623]), .A(ram[559]), .S(n4309), .Y(n3584) );
  MUX2X1 U6870 ( .B(ram[751]), .A(ram[687]), .S(n4309), .Y(n3583) );
  MUX2X1 U6871 ( .B(ram[879]), .A(ram[815]), .S(n4309), .Y(n3587) );
  MUX2X1 U6872 ( .B(ram[1007]), .A(ram[943]), .S(n4309), .Y(n3586) );
  MUX2X1 U6873 ( .B(n3585), .A(n3582), .S(n4172), .Y(n3589) );
  MUX2X1 U6874 ( .B(ram[1135]), .A(ram[1071]), .S(n4310), .Y(n3593) );
  MUX2X1 U6875 ( .B(ram[1263]), .A(ram[1199]), .S(n4310), .Y(n3592) );
  MUX2X1 U6876 ( .B(ram[1391]), .A(ram[1327]), .S(n4310), .Y(n3596) );
  MUX2X1 U6877 ( .B(ram[1519]), .A(ram[1455]), .S(n4310), .Y(n3595) );
  MUX2X1 U6878 ( .B(n3594), .A(n3591), .S(n4172), .Y(n3605) );
  MUX2X1 U6879 ( .B(ram[1647]), .A(ram[1583]), .S(n4310), .Y(n3599) );
  MUX2X1 U6880 ( .B(ram[1775]), .A(ram[1711]), .S(n4310), .Y(n3598) );
  MUX2X1 U6881 ( .B(ram[1903]), .A(ram[1839]), .S(n4310), .Y(n3602) );
  MUX2X1 U6882 ( .B(ram[2031]), .A(ram[1967]), .S(n4310), .Y(n3601) );
  MUX2X1 U6883 ( .B(n3600), .A(n3597), .S(n4172), .Y(n3604) );
  MUX2X1 U6884 ( .B(n3603), .A(n3588), .S(n4151), .Y(n4133) );
  MUX2X1 U6885 ( .B(ram[112]), .A(ram[48]), .S(n4310), .Y(n3608) );
  MUX2X1 U6886 ( .B(ram[240]), .A(ram[176]), .S(n4310), .Y(n3607) );
  MUX2X1 U6887 ( .B(ram[368]), .A(ram[304]), .S(n4310), .Y(n3611) );
  MUX2X1 U6888 ( .B(ram[496]), .A(ram[432]), .S(n4310), .Y(n3610) );
  MUX2X1 U6889 ( .B(n3609), .A(n3606), .S(n4172), .Y(n3620) );
  MUX2X1 U6890 ( .B(ram[624]), .A(ram[560]), .S(n4311), .Y(n3614) );
  MUX2X1 U6891 ( .B(ram[752]), .A(ram[688]), .S(n4311), .Y(n3613) );
  MUX2X1 U6892 ( .B(ram[880]), .A(ram[816]), .S(n4311), .Y(n3617) );
  MUX2X1 U6893 ( .B(ram[1008]), .A(ram[944]), .S(n4311), .Y(n3616) );
  MUX2X1 U6894 ( .B(n3615), .A(n3612), .S(n4172), .Y(n3619) );
  MUX2X1 U6895 ( .B(ram[1136]), .A(ram[1072]), .S(n4311), .Y(n3623) );
  MUX2X1 U6896 ( .B(ram[1264]), .A(ram[1200]), .S(n4311), .Y(n3622) );
  MUX2X1 U6897 ( .B(ram[1392]), .A(ram[1328]), .S(n4311), .Y(n3626) );
  MUX2X1 U6898 ( .B(ram[1520]), .A(ram[1456]), .S(n4311), .Y(n3625) );
  MUX2X1 U6899 ( .B(n3624), .A(n3621), .S(n4172), .Y(n3635) );
  MUX2X1 U6900 ( .B(ram[1648]), .A(ram[1584]), .S(n4311), .Y(n3629) );
  MUX2X1 U6901 ( .B(ram[1776]), .A(ram[1712]), .S(n4311), .Y(n3628) );
  MUX2X1 U6902 ( .B(ram[1904]), .A(ram[1840]), .S(n4311), .Y(n3632) );
  MUX2X1 U6903 ( .B(ram[2032]), .A(ram[1968]), .S(n4311), .Y(n3631) );
  MUX2X1 U6904 ( .B(n3630), .A(n3627), .S(n4172), .Y(n3634) );
  MUX2X1 U6905 ( .B(n3633), .A(n3618), .S(n4150), .Y(n4134) );
  MUX2X1 U6906 ( .B(ram[113]), .A(ram[49]), .S(n4312), .Y(n3638) );
  MUX2X1 U6907 ( .B(ram[241]), .A(ram[177]), .S(n4312), .Y(n3637) );
  MUX2X1 U6908 ( .B(ram[369]), .A(ram[305]), .S(n4312), .Y(n3641) );
  MUX2X1 U6909 ( .B(ram[497]), .A(ram[433]), .S(n4312), .Y(n3640) );
  MUX2X1 U6910 ( .B(n3639), .A(n3636), .S(n4173), .Y(n3650) );
  MUX2X1 U6911 ( .B(ram[625]), .A(ram[561]), .S(n4312), .Y(n3644) );
  MUX2X1 U6912 ( .B(ram[753]), .A(ram[689]), .S(n4312), .Y(n3643) );
  MUX2X1 U6913 ( .B(ram[881]), .A(ram[817]), .S(n4312), .Y(n3647) );
  MUX2X1 U6914 ( .B(ram[1009]), .A(ram[945]), .S(n4312), .Y(n3646) );
  MUX2X1 U6915 ( .B(n3645), .A(n3642), .S(n4173), .Y(n3649) );
  MUX2X1 U6916 ( .B(ram[1137]), .A(ram[1073]), .S(n4312), .Y(n3653) );
  MUX2X1 U6917 ( .B(ram[1265]), .A(ram[1201]), .S(n4312), .Y(n3652) );
  MUX2X1 U6918 ( .B(ram[1393]), .A(ram[1329]), .S(n4312), .Y(n3656) );
  MUX2X1 U6919 ( .B(ram[1521]), .A(ram[1457]), .S(n4312), .Y(n3655) );
  MUX2X1 U6920 ( .B(n3654), .A(n3651), .S(n4173), .Y(n3665) );
  MUX2X1 U6921 ( .B(ram[1649]), .A(ram[1585]), .S(n4313), .Y(n3659) );
  MUX2X1 U6922 ( .B(ram[1777]), .A(ram[1713]), .S(n4313), .Y(n3658) );
  MUX2X1 U6923 ( .B(ram[1905]), .A(ram[1841]), .S(n4313), .Y(n3662) );
  MUX2X1 U6924 ( .B(ram[2033]), .A(ram[1969]), .S(n4313), .Y(n3661) );
  MUX2X1 U6925 ( .B(n3660), .A(n3657), .S(n4173), .Y(n3664) );
  MUX2X1 U6926 ( .B(n3663), .A(n3648), .S(n4150), .Y(n4135) );
  MUX2X1 U6927 ( .B(ram[114]), .A(ram[50]), .S(n4313), .Y(n3668) );
  MUX2X1 U6928 ( .B(ram[242]), .A(ram[178]), .S(n4313), .Y(n3667) );
  MUX2X1 U6929 ( .B(ram[370]), .A(ram[306]), .S(n4313), .Y(n3671) );
  MUX2X1 U6930 ( .B(ram[498]), .A(ram[434]), .S(n4313), .Y(n3670) );
  MUX2X1 U6931 ( .B(n3669), .A(n3666), .S(n4173), .Y(n3680) );
  MUX2X1 U6932 ( .B(ram[626]), .A(ram[562]), .S(n4313), .Y(n3674) );
  MUX2X1 U6933 ( .B(ram[754]), .A(ram[690]), .S(n4313), .Y(n3673) );
  MUX2X1 U6934 ( .B(ram[882]), .A(ram[818]), .S(n4313), .Y(n3677) );
  MUX2X1 U6935 ( .B(ram[1010]), .A(ram[946]), .S(n4313), .Y(n3676) );
  MUX2X1 U6936 ( .B(n3675), .A(n3672), .S(n4173), .Y(n3679) );
  MUX2X1 U6937 ( .B(ram[1138]), .A(ram[1074]), .S(n4314), .Y(n3683) );
  MUX2X1 U6938 ( .B(ram[1266]), .A(ram[1202]), .S(n4314), .Y(n3682) );
  MUX2X1 U6939 ( .B(ram[1394]), .A(ram[1330]), .S(n4314), .Y(n3686) );
  MUX2X1 U6940 ( .B(ram[1522]), .A(ram[1458]), .S(n4314), .Y(n3685) );
  MUX2X1 U6941 ( .B(n3684), .A(n3681), .S(n4173), .Y(n3695) );
  MUX2X1 U6942 ( .B(ram[1650]), .A(ram[1586]), .S(n4314), .Y(n3689) );
  MUX2X1 U6943 ( .B(ram[1778]), .A(ram[1714]), .S(n4314), .Y(n3688) );
  MUX2X1 U6944 ( .B(ram[1906]), .A(ram[1842]), .S(n4314), .Y(n3692) );
  MUX2X1 U6945 ( .B(ram[2034]), .A(ram[1970]), .S(n4314), .Y(n3691) );
  MUX2X1 U6946 ( .B(n3690), .A(n3687), .S(n4173), .Y(n3694) );
  MUX2X1 U6947 ( .B(n3693), .A(n3678), .S(n4150), .Y(n4136) );
  MUX2X1 U6948 ( .B(ram[115]), .A(ram[51]), .S(n4314), .Y(n3698) );
  MUX2X1 U6949 ( .B(ram[243]), .A(ram[179]), .S(n4314), .Y(n3697) );
  MUX2X1 U6950 ( .B(ram[371]), .A(ram[307]), .S(n4314), .Y(n3701) );
  MUX2X1 U6951 ( .B(ram[499]), .A(ram[435]), .S(n4314), .Y(n3700) );
  MUX2X1 U6952 ( .B(n3699), .A(n3696), .S(n4173), .Y(n3710) );
  MUX2X1 U6953 ( .B(ram[627]), .A(ram[563]), .S(n4315), .Y(n3704) );
  MUX2X1 U6954 ( .B(ram[755]), .A(ram[691]), .S(n4299), .Y(n3703) );
  MUX2X1 U6955 ( .B(ram[883]), .A(ram[819]), .S(n4314), .Y(n3707) );
  MUX2X1 U6956 ( .B(ram[1011]), .A(ram[947]), .S(n4305), .Y(n3706) );
  MUX2X1 U6957 ( .B(n3705), .A(n3702), .S(n4173), .Y(n3709) );
  MUX2X1 U6958 ( .B(ram[1139]), .A(ram[1075]), .S(n4319), .Y(n3713) );
  MUX2X1 U6959 ( .B(ram[1267]), .A(ram[1203]), .S(n4301), .Y(n3712) );
  MUX2X1 U6960 ( .B(ram[1395]), .A(ram[1331]), .S(n4316), .Y(n3716) );
  MUX2X1 U6961 ( .B(ram[1523]), .A(ram[1459]), .S(n4322), .Y(n3715) );
  MUX2X1 U6962 ( .B(n3714), .A(n3711), .S(n4173), .Y(n3725) );
  MUX2X1 U6963 ( .B(ram[1651]), .A(ram[1587]), .S(n4316), .Y(n3719) );
  MUX2X1 U6964 ( .B(ram[1779]), .A(ram[1715]), .S(n4320), .Y(n3718) );
  MUX2X1 U6965 ( .B(ram[1907]), .A(ram[1843]), .S(n4314), .Y(n3722) );
  MUX2X1 U6966 ( .B(ram[2035]), .A(ram[1971]), .S(n4317), .Y(n3721) );
  MUX2X1 U6967 ( .B(n3720), .A(n3717), .S(n4173), .Y(n3724) );
  MUX2X1 U6968 ( .B(n3723), .A(n3708), .S(n4150), .Y(n4137) );
  MUX2X1 U6969 ( .B(ram[116]), .A(ram[52]), .S(n4315), .Y(n3728) );
  MUX2X1 U6970 ( .B(ram[244]), .A(ram[180]), .S(n4315), .Y(n3727) );
  MUX2X1 U6971 ( .B(ram[372]), .A(ram[308]), .S(n4315), .Y(n3731) );
  MUX2X1 U6972 ( .B(ram[500]), .A(ram[436]), .S(n4315), .Y(n3730) );
  MUX2X1 U6973 ( .B(n3729), .A(n3726), .S(n4174), .Y(n3740) );
  MUX2X1 U6974 ( .B(ram[628]), .A(ram[564]), .S(n4315), .Y(n3734) );
  MUX2X1 U6975 ( .B(ram[756]), .A(ram[692]), .S(n4315), .Y(n3733) );
  MUX2X1 U6976 ( .B(ram[884]), .A(ram[820]), .S(n4315), .Y(n3737) );
  MUX2X1 U6977 ( .B(ram[1012]), .A(ram[948]), .S(n4315), .Y(n3736) );
  MUX2X1 U6978 ( .B(n3735), .A(n3732), .S(n4174), .Y(n3739) );
  MUX2X1 U6979 ( .B(ram[1140]), .A(ram[1076]), .S(n4315), .Y(n3743) );
  MUX2X1 U6980 ( .B(ram[1268]), .A(ram[1204]), .S(n4315), .Y(n3742) );
  MUX2X1 U6981 ( .B(ram[1396]), .A(ram[1332]), .S(n4315), .Y(n3746) );
  MUX2X1 U6982 ( .B(ram[1524]), .A(ram[1460]), .S(n4315), .Y(n3745) );
  MUX2X1 U6983 ( .B(n3744), .A(n3741), .S(n4174), .Y(n3755) );
  MUX2X1 U6984 ( .B(ram[1652]), .A(ram[1588]), .S(n4316), .Y(n3749) );
  MUX2X1 U6985 ( .B(ram[1780]), .A(ram[1716]), .S(n4316), .Y(n3748) );
  MUX2X1 U6986 ( .B(ram[1908]), .A(ram[1844]), .S(n4316), .Y(n3752) );
  MUX2X1 U6987 ( .B(ram[2036]), .A(ram[1972]), .S(n4316), .Y(n3751) );
  MUX2X1 U6988 ( .B(n3750), .A(n3747), .S(n4174), .Y(n3754) );
  MUX2X1 U6989 ( .B(n3753), .A(n3738), .S(n4150), .Y(n4138) );
  MUX2X1 U6990 ( .B(ram[117]), .A(ram[53]), .S(n4316), .Y(n3758) );
  MUX2X1 U6991 ( .B(ram[245]), .A(ram[181]), .S(n4316), .Y(n3757) );
  MUX2X1 U6992 ( .B(ram[373]), .A(ram[309]), .S(n4316), .Y(n3761) );
  MUX2X1 U6993 ( .B(ram[501]), .A(ram[437]), .S(n4316), .Y(n3760) );
  MUX2X1 U6994 ( .B(n3759), .A(n3756), .S(n4174), .Y(n3770) );
  MUX2X1 U6995 ( .B(ram[629]), .A(ram[565]), .S(n4316), .Y(n3764) );
  MUX2X1 U6996 ( .B(ram[757]), .A(ram[693]), .S(n4316), .Y(n3763) );
  MUX2X1 U6997 ( .B(ram[885]), .A(ram[821]), .S(n4316), .Y(n3767) );
  MUX2X1 U6998 ( .B(ram[1013]), .A(ram[949]), .S(n4316), .Y(n3766) );
  MUX2X1 U6999 ( .B(n3765), .A(n3762), .S(n4174), .Y(n3769) );
  MUX2X1 U7000 ( .B(ram[1141]), .A(ram[1077]), .S(n4317), .Y(n3773) );
  MUX2X1 U7001 ( .B(ram[1269]), .A(ram[1205]), .S(n4317), .Y(n3772) );
  MUX2X1 U7002 ( .B(ram[1397]), .A(ram[1333]), .S(n4317), .Y(n3776) );
  MUX2X1 U7003 ( .B(ram[1525]), .A(ram[1461]), .S(n4317), .Y(n3775) );
  MUX2X1 U7004 ( .B(n3774), .A(n3771), .S(n4174), .Y(n3785) );
  MUX2X1 U7005 ( .B(ram[1653]), .A(ram[1589]), .S(n4317), .Y(n3779) );
  MUX2X1 U7006 ( .B(ram[1781]), .A(ram[1717]), .S(n4317), .Y(n3778) );
  MUX2X1 U7007 ( .B(ram[1909]), .A(ram[1845]), .S(n4317), .Y(n3782) );
  MUX2X1 U7008 ( .B(ram[2037]), .A(ram[1973]), .S(n4317), .Y(n3781) );
  MUX2X1 U7009 ( .B(n3780), .A(n3777), .S(n4174), .Y(n3784) );
  MUX2X1 U7010 ( .B(n3783), .A(n3768), .S(n4150), .Y(n4139) );
  MUX2X1 U7011 ( .B(ram[118]), .A(ram[54]), .S(n4317), .Y(n3788) );
  MUX2X1 U7012 ( .B(ram[246]), .A(ram[182]), .S(n4317), .Y(n3787) );
  MUX2X1 U7013 ( .B(ram[374]), .A(ram[310]), .S(n4317), .Y(n3791) );
  MUX2X1 U7014 ( .B(ram[502]), .A(ram[438]), .S(n4317), .Y(n3790) );
  MUX2X1 U7015 ( .B(n3789), .A(n3786), .S(n4174), .Y(n3800) );
  MUX2X1 U7016 ( .B(ram[630]), .A(ram[566]), .S(n4318), .Y(n3794) );
  MUX2X1 U7017 ( .B(ram[758]), .A(ram[694]), .S(n4318), .Y(n3793) );
  MUX2X1 U7018 ( .B(ram[886]), .A(ram[822]), .S(n4318), .Y(n3797) );
  MUX2X1 U7019 ( .B(ram[1014]), .A(ram[950]), .S(n4318), .Y(n3796) );
  MUX2X1 U7020 ( .B(n3795), .A(n3792), .S(n4174), .Y(n3799) );
  MUX2X1 U7021 ( .B(ram[1142]), .A(ram[1078]), .S(n4318), .Y(n3803) );
  MUX2X1 U7022 ( .B(ram[1270]), .A(ram[1206]), .S(n4318), .Y(n3802) );
  MUX2X1 U7023 ( .B(ram[1398]), .A(ram[1334]), .S(n4318), .Y(n3806) );
  MUX2X1 U7024 ( .B(ram[1526]), .A(ram[1462]), .S(n4318), .Y(n3805) );
  MUX2X1 U7025 ( .B(n3804), .A(n3801), .S(n4174), .Y(n3815) );
  MUX2X1 U7026 ( .B(ram[1654]), .A(ram[1590]), .S(n4318), .Y(n3809) );
  MUX2X1 U7027 ( .B(ram[1782]), .A(ram[1718]), .S(n4318), .Y(n3808) );
  MUX2X1 U7028 ( .B(ram[1910]), .A(ram[1846]), .S(n4318), .Y(n3812) );
  MUX2X1 U7029 ( .B(ram[2038]), .A(ram[1974]), .S(n4318), .Y(n3811) );
  MUX2X1 U7030 ( .B(n3810), .A(n3807), .S(n4174), .Y(n3814) );
  MUX2X1 U7031 ( .B(n3813), .A(n3798), .S(n4150), .Y(n4140) );
  MUX2X1 U7032 ( .B(ram[119]), .A(ram[55]), .S(n4319), .Y(n3818) );
  MUX2X1 U7033 ( .B(ram[247]), .A(ram[183]), .S(n4319), .Y(n3817) );
  MUX2X1 U7034 ( .B(ram[375]), .A(ram[311]), .S(n4319), .Y(n3821) );
  MUX2X1 U7035 ( .B(ram[503]), .A(ram[439]), .S(n4319), .Y(n3820) );
  MUX2X1 U7036 ( .B(n3819), .A(n3816), .S(n4175), .Y(n3830) );
  MUX2X1 U7037 ( .B(ram[631]), .A(ram[567]), .S(n4319), .Y(n3824) );
  MUX2X1 U7038 ( .B(ram[759]), .A(ram[695]), .S(n4319), .Y(n3823) );
  MUX2X1 U7039 ( .B(ram[887]), .A(ram[823]), .S(n4319), .Y(n3827) );
  MUX2X1 U7040 ( .B(ram[1015]), .A(ram[951]), .S(n4319), .Y(n3826) );
  MUX2X1 U7041 ( .B(n3825), .A(n3822), .S(n4175), .Y(n3829) );
  MUX2X1 U7042 ( .B(ram[1143]), .A(ram[1079]), .S(n4319), .Y(n3833) );
  MUX2X1 U7043 ( .B(ram[1271]), .A(ram[1207]), .S(n4319), .Y(n3832) );
  MUX2X1 U7044 ( .B(ram[1399]), .A(ram[1335]), .S(n4319), .Y(n3836) );
  MUX2X1 U7045 ( .B(ram[1527]), .A(ram[1463]), .S(n4319), .Y(n3835) );
  MUX2X1 U7046 ( .B(n3834), .A(n3831), .S(n4175), .Y(n3845) );
  MUX2X1 U7047 ( .B(ram[1655]), .A(ram[1591]), .S(n4320), .Y(n3839) );
  MUX2X1 U7048 ( .B(ram[1783]), .A(ram[1719]), .S(n4320), .Y(n3838) );
  MUX2X1 U7049 ( .B(ram[1911]), .A(ram[1847]), .S(n4320), .Y(n3842) );
  MUX2X1 U7050 ( .B(ram[2039]), .A(ram[1975]), .S(n4320), .Y(n3841) );
  MUX2X1 U7051 ( .B(n3840), .A(n3837), .S(n4175), .Y(n3844) );
  MUX2X1 U7052 ( .B(n3843), .A(n3828), .S(n4150), .Y(n4141) );
  MUX2X1 U7053 ( .B(ram[120]), .A(ram[56]), .S(n4320), .Y(n3848) );
  MUX2X1 U7054 ( .B(ram[248]), .A(ram[184]), .S(n4320), .Y(n3847) );
  MUX2X1 U7055 ( .B(ram[376]), .A(ram[312]), .S(n4320), .Y(n3851) );
  MUX2X1 U7056 ( .B(ram[504]), .A(ram[440]), .S(n4320), .Y(n3850) );
  MUX2X1 U7057 ( .B(n3849), .A(n3846), .S(n4175), .Y(n3860) );
  MUX2X1 U7058 ( .B(ram[632]), .A(ram[568]), .S(n4320), .Y(n3854) );
  MUX2X1 U7059 ( .B(ram[760]), .A(ram[696]), .S(n4320), .Y(n3853) );
  MUX2X1 U7060 ( .B(ram[888]), .A(ram[824]), .S(n4320), .Y(n3857) );
  MUX2X1 U7061 ( .B(ram[1016]), .A(ram[952]), .S(n4320), .Y(n3856) );
  MUX2X1 U7062 ( .B(n3855), .A(n3852), .S(n4175), .Y(n3859) );
  MUX2X1 U7063 ( .B(ram[1144]), .A(ram[1080]), .S(n4321), .Y(n3863) );
  MUX2X1 U7064 ( .B(ram[1272]), .A(ram[1208]), .S(n4321), .Y(n3862) );
  MUX2X1 U7065 ( .B(ram[1400]), .A(ram[1336]), .S(n4321), .Y(n3866) );
  MUX2X1 U7066 ( .B(ram[1528]), .A(ram[1464]), .S(n4321), .Y(n3865) );
  MUX2X1 U7067 ( .B(n3864), .A(n3861), .S(n4175), .Y(n3875) );
  MUX2X1 U7068 ( .B(ram[1656]), .A(ram[1592]), .S(n4321), .Y(n3869) );
  MUX2X1 U7069 ( .B(ram[1784]), .A(ram[1720]), .S(n4321), .Y(n3868) );
  MUX2X1 U7070 ( .B(ram[1912]), .A(ram[1848]), .S(n4321), .Y(n3872) );
  MUX2X1 U7071 ( .B(ram[2040]), .A(ram[1976]), .S(n4321), .Y(n3871) );
  MUX2X1 U7072 ( .B(n3870), .A(n3867), .S(n4175), .Y(n3874) );
  MUX2X1 U7073 ( .B(n3873), .A(n3858), .S(n4150), .Y(n4142) );
  MUX2X1 U7074 ( .B(ram[121]), .A(ram[57]), .S(n4321), .Y(n3878) );
  MUX2X1 U7075 ( .B(ram[249]), .A(ram[185]), .S(n4321), .Y(n3877) );
  MUX2X1 U7076 ( .B(ram[377]), .A(ram[313]), .S(n4321), .Y(n3881) );
  MUX2X1 U7077 ( .B(ram[505]), .A(ram[441]), .S(n4321), .Y(n3880) );
  MUX2X1 U7078 ( .B(n3879), .A(n3876), .S(n4175), .Y(n3890) );
  MUX2X1 U7079 ( .B(ram[633]), .A(ram[569]), .S(n4322), .Y(n3884) );
  MUX2X1 U7080 ( .B(ram[761]), .A(ram[697]), .S(n4322), .Y(n3883) );
  MUX2X1 U7081 ( .B(ram[889]), .A(ram[825]), .S(n4322), .Y(n3887) );
  MUX2X1 U7082 ( .B(ram[1017]), .A(ram[953]), .S(n4322), .Y(n3886) );
  MUX2X1 U7083 ( .B(n3885), .A(n3882), .S(n4175), .Y(n3889) );
  MUX2X1 U7084 ( .B(ram[1145]), .A(ram[1081]), .S(n4322), .Y(n3893) );
  MUX2X1 U7085 ( .B(ram[1273]), .A(ram[1209]), .S(n4322), .Y(n3892) );
  MUX2X1 U7086 ( .B(ram[1401]), .A(ram[1337]), .S(n4322), .Y(n3896) );
  MUX2X1 U7087 ( .B(ram[1529]), .A(ram[1465]), .S(n4322), .Y(n3895) );
  MUX2X1 U7088 ( .B(n3894), .A(n3891), .S(n4175), .Y(n3905) );
  MUX2X1 U7089 ( .B(ram[1657]), .A(ram[1593]), .S(n4322), .Y(n3899) );
  MUX2X1 U7090 ( .B(ram[1785]), .A(ram[1721]), .S(n4322), .Y(n3898) );
  MUX2X1 U7091 ( .B(ram[1913]), .A(ram[1849]), .S(n4322), .Y(n3902) );
  MUX2X1 U7092 ( .B(ram[2041]), .A(ram[1977]), .S(n4322), .Y(n3901) );
  MUX2X1 U7093 ( .B(n3900), .A(n3897), .S(n4175), .Y(n3904) );
  MUX2X1 U7094 ( .B(n3903), .A(n3888), .S(n4150), .Y(n4143) );
  MUX2X1 U7095 ( .B(ram[122]), .A(ram[58]), .S(n4323), .Y(n3908) );
  MUX2X1 U7096 ( .B(ram[250]), .A(ram[186]), .S(n4323), .Y(n3907) );
  MUX2X1 U7097 ( .B(ram[378]), .A(ram[314]), .S(n4323), .Y(n3911) );
  MUX2X1 U7098 ( .B(ram[506]), .A(ram[442]), .S(n4323), .Y(n3910) );
  MUX2X1 U7099 ( .B(n3909), .A(n3906), .S(n4174), .Y(n3920) );
  MUX2X1 U7100 ( .B(ram[634]), .A(ram[570]), .S(n4323), .Y(n3914) );
  MUX2X1 U7101 ( .B(ram[762]), .A(ram[698]), .S(n4323), .Y(n3913) );
  MUX2X1 U7102 ( .B(ram[890]), .A(ram[826]), .S(n4323), .Y(n3917) );
  MUX2X1 U7103 ( .B(ram[1018]), .A(ram[954]), .S(n4323), .Y(n3916) );
  MUX2X1 U7104 ( .B(n3915), .A(n3912), .S(n4171), .Y(n3919) );
  MUX2X1 U7105 ( .B(ram[1146]), .A(ram[1082]), .S(n4323), .Y(n3923) );
  MUX2X1 U7106 ( .B(ram[1274]), .A(ram[1210]), .S(n4323), .Y(n3922) );
  MUX2X1 U7107 ( .B(ram[1402]), .A(ram[1338]), .S(n4323), .Y(n3926) );
  MUX2X1 U7108 ( .B(ram[1530]), .A(ram[1466]), .S(n4323), .Y(n3925) );
  MUX2X1 U7109 ( .B(n3924), .A(n3921), .S(n4175), .Y(n3935) );
  MUX2X1 U7110 ( .B(ram[1658]), .A(ram[1594]), .S(n4328), .Y(n3929) );
  MUX2X1 U7111 ( .B(ram[1786]), .A(ram[1722]), .S(n4327), .Y(n3928) );
  MUX2X1 U7112 ( .B(ram[1914]), .A(ram[1850]), .S(n4323), .Y(n3932) );
  MUX2X1 U7113 ( .B(ram[2042]), .A(ram[1978]), .S(n4329), .Y(n3931) );
  MUX2X1 U7114 ( .B(n3930), .A(n3927), .S(n4168), .Y(n3934) );
  MUX2X1 U7115 ( .B(n3933), .A(n3918), .S(n4150), .Y(n4144) );
  MUX2X1 U7116 ( .B(ram[123]), .A(ram[59]), .S(n4329), .Y(n3938) );
  MUX2X1 U7117 ( .B(ram[251]), .A(ram[187]), .S(n4309), .Y(n3937) );
  MUX2X1 U7118 ( .B(ram[379]), .A(ram[315]), .S(n4323), .Y(n3941) );
  MUX2X1 U7119 ( .B(ram[507]), .A(ram[443]), .S(n4294), .Y(n3940) );
  MUX2X1 U7120 ( .B(n3939), .A(n3936), .S(n4173), .Y(n3950) );
  MUX2X1 U7121 ( .B(ram[635]), .A(ram[571]), .S(n4298), .Y(n3944) );
  MUX2X1 U7122 ( .B(ram[763]), .A(ram[699]), .S(n4305), .Y(n3943) );
  MUX2X1 U7123 ( .B(ram[891]), .A(ram[827]), .S(n4309), .Y(n3947) );
  MUX2X1 U7124 ( .B(ram[1019]), .A(ram[955]), .S(n4323), .Y(n3946) );
  MUX2X1 U7125 ( .B(n3945), .A(n3942), .S(n4172), .Y(n3949) );
  MUX2X1 U7126 ( .B(ram[1147]), .A(ram[1083]), .S(n4324), .Y(n3953) );
  MUX2X1 U7127 ( .B(ram[1275]), .A(ram[1211]), .S(n4324), .Y(n3952) );
  MUX2X1 U7128 ( .B(ram[1403]), .A(ram[1339]), .S(n4324), .Y(n3956) );
  MUX2X1 U7129 ( .B(ram[1531]), .A(ram[1467]), .S(n4324), .Y(n3955) );
  MUX2X1 U7130 ( .B(n3954), .A(n3951), .S(n4169), .Y(n3965) );
  MUX2X1 U7131 ( .B(ram[1659]), .A(ram[1595]), .S(n4324), .Y(n3959) );
  MUX2X1 U7132 ( .B(ram[1787]), .A(ram[1723]), .S(n4324), .Y(n3958) );
  MUX2X1 U7133 ( .B(ram[1915]), .A(ram[1851]), .S(n4324), .Y(n3962) );
  MUX2X1 U7134 ( .B(ram[2043]), .A(ram[1979]), .S(n4324), .Y(n3961) );
  MUX2X1 U7135 ( .B(n3960), .A(n3957), .S(n4170), .Y(n3964) );
  MUX2X1 U7136 ( .B(n3963), .A(n3948), .S(n4150), .Y(n4145) );
  MUX2X1 U7137 ( .B(ram[124]), .A(ram[60]), .S(n4324), .Y(n3968) );
  MUX2X1 U7138 ( .B(ram[252]), .A(ram[188]), .S(n4324), .Y(n3967) );
  MUX2X1 U7139 ( .B(ram[380]), .A(ram[316]), .S(n4324), .Y(n3971) );
  MUX2X1 U7140 ( .B(ram[508]), .A(ram[444]), .S(n4324), .Y(n3970) );
  MUX2X1 U7141 ( .B(n3969), .A(n3966), .S(n4174), .Y(n3980) );
  MUX2X1 U7142 ( .B(ram[636]), .A(ram[572]), .S(n4325), .Y(n3974) );
  MUX2X1 U7143 ( .B(ram[764]), .A(ram[700]), .S(n4325), .Y(n3973) );
  MUX2X1 U7144 ( .B(ram[892]), .A(ram[828]), .S(n4325), .Y(n3977) );
  MUX2X1 U7145 ( .B(ram[1020]), .A(ram[956]), .S(n4325), .Y(n3976) );
  MUX2X1 U7146 ( .B(n3975), .A(n3972), .S(n4169), .Y(n3979) );
  MUX2X1 U7147 ( .B(ram[1148]), .A(ram[1084]), .S(n4325), .Y(n3983) );
  MUX2X1 U7148 ( .B(ram[1276]), .A(ram[1212]), .S(n4325), .Y(n3982) );
  MUX2X1 U7149 ( .B(ram[1404]), .A(ram[1340]), .S(n4325), .Y(n3986) );
  MUX2X1 U7150 ( .B(ram[1532]), .A(ram[1468]), .S(n4325), .Y(n3985) );
  MUX2X1 U7151 ( .B(n3984), .A(n3981), .S(n4175), .Y(n3995) );
  MUX2X1 U7152 ( .B(ram[1660]), .A(ram[1596]), .S(n4325), .Y(n3989) );
  MUX2X1 U7153 ( .B(ram[1788]), .A(ram[1724]), .S(n4325), .Y(n3988) );
  MUX2X1 U7154 ( .B(ram[1916]), .A(ram[1852]), .S(n4325), .Y(n3992) );
  MUX2X1 U7155 ( .B(ram[2044]), .A(ram[1980]), .S(n4325), .Y(n3991) );
  MUX2X1 U7156 ( .B(n3990), .A(n3987), .S(n4168), .Y(n3994) );
  MUX2X1 U7157 ( .B(n3993), .A(n3978), .S(n4151), .Y(n4146) );
  MUX2X1 U7158 ( .B(ram[125]), .A(ram[61]), .S(n4326), .Y(n3998) );
  MUX2X1 U7159 ( .B(ram[253]), .A(ram[189]), .S(n4326), .Y(n3997) );
  MUX2X1 U7160 ( .B(ram[381]), .A(ram[317]), .S(n4326), .Y(n4001) );
  MUX2X1 U7161 ( .B(ram[509]), .A(ram[445]), .S(n4326), .Y(n4000) );
  MUX2X1 U7162 ( .B(n3999), .A(n3996), .S(n4170), .Y(n4010) );
  MUX2X1 U7163 ( .B(ram[637]), .A(ram[573]), .S(n4326), .Y(n4004) );
  MUX2X1 U7164 ( .B(ram[765]), .A(ram[701]), .S(n4326), .Y(n4003) );
  MUX2X1 U7165 ( .B(ram[893]), .A(ram[829]), .S(n4326), .Y(n4007) );
  MUX2X1 U7166 ( .B(ram[1021]), .A(ram[957]), .S(n4326), .Y(n4006) );
  MUX2X1 U7167 ( .B(n4005), .A(n4002), .S(n4173), .Y(n4009) );
  MUX2X1 U7168 ( .B(ram[1149]), .A(ram[1085]), .S(n4326), .Y(n4013) );
  MUX2X1 U7169 ( .B(ram[1277]), .A(ram[1213]), .S(n4326), .Y(n4012) );
  MUX2X1 U7170 ( .B(ram[1405]), .A(ram[1341]), .S(n4326), .Y(n4016) );
  MUX2X1 U7171 ( .B(ram[1533]), .A(ram[1469]), .S(n4326), .Y(n4015) );
  MUX2X1 U7172 ( .B(n4014), .A(n4011), .S(n4175), .Y(n4025) );
  MUX2X1 U7173 ( .B(ram[1661]), .A(ram[1597]), .S(n4327), .Y(n4019) );
  MUX2X1 U7174 ( .B(ram[1789]), .A(ram[1725]), .S(n4327), .Y(n4018) );
  MUX2X1 U7175 ( .B(ram[1917]), .A(ram[1853]), .S(n4327), .Y(n4022) );
  MUX2X1 U7176 ( .B(ram[2045]), .A(ram[1981]), .S(n4327), .Y(n4021) );
  MUX2X1 U7177 ( .B(n4020), .A(n4017), .S(n4168), .Y(n4024) );
  MUX2X1 U7178 ( .B(n4023), .A(n4008), .S(n4150), .Y(n4147) );
  MUX2X1 U7179 ( .B(ram[126]), .A(ram[62]), .S(n4327), .Y(n4028) );
  MUX2X1 U7180 ( .B(ram[254]), .A(ram[190]), .S(n4327), .Y(n4027) );
  MUX2X1 U7181 ( .B(ram[382]), .A(ram[318]), .S(n4327), .Y(n4031) );
  MUX2X1 U7182 ( .B(ram[510]), .A(ram[446]), .S(n4327), .Y(n4030) );
  MUX2X1 U7183 ( .B(n4029), .A(n4026), .S(n4169), .Y(n4040) );
  MUX2X1 U7184 ( .B(ram[638]), .A(ram[574]), .S(n4327), .Y(n4034) );
  MUX2X1 U7185 ( .B(ram[766]), .A(ram[702]), .S(n4327), .Y(n4033) );
  MUX2X1 U7186 ( .B(ram[894]), .A(ram[830]), .S(n4327), .Y(n4037) );
  MUX2X1 U7187 ( .B(ram[1022]), .A(ram[958]), .S(n4327), .Y(n4036) );
  MUX2X1 U7188 ( .B(n4035), .A(n4032), .S(n4171), .Y(n4039) );
  MUX2X1 U7189 ( .B(ram[1150]), .A(ram[1086]), .S(n4328), .Y(n4043) );
  MUX2X1 U7190 ( .B(ram[1278]), .A(ram[1214]), .S(n4328), .Y(n4042) );
  MUX2X1 U7191 ( .B(ram[1406]), .A(ram[1342]), .S(n4328), .Y(n4046) );
  MUX2X1 U7192 ( .B(ram[1534]), .A(ram[1470]), .S(n4328), .Y(n4045) );
  MUX2X1 U7193 ( .B(n4044), .A(n4041), .S(n4172), .Y(n4055) );
  MUX2X1 U7194 ( .B(ram[1662]), .A(ram[1598]), .S(n4328), .Y(n4049) );
  MUX2X1 U7195 ( .B(ram[1790]), .A(ram[1726]), .S(n4328), .Y(n4048) );
  MUX2X1 U7196 ( .B(ram[1918]), .A(ram[1854]), .S(n4328), .Y(n4052) );
  MUX2X1 U7197 ( .B(ram[2046]), .A(ram[1982]), .S(n4328), .Y(n4051) );
  MUX2X1 U7198 ( .B(n4050), .A(n4047), .S(n4174), .Y(n4054) );
  MUX2X1 U7199 ( .B(n4053), .A(n4038), .S(n4151), .Y(n4148) );
  MUX2X1 U7200 ( .B(ram[127]), .A(ram[63]), .S(n4328), .Y(n4058) );
  MUX2X1 U7201 ( .B(ram[255]), .A(ram[191]), .S(n4328), .Y(n4057) );
  MUX2X1 U7202 ( .B(ram[383]), .A(ram[319]), .S(n4328), .Y(n4061) );
  MUX2X1 U7203 ( .B(ram[511]), .A(ram[447]), .S(n4328), .Y(n4060) );
  MUX2X1 U7204 ( .B(n4059), .A(n4056), .S(n4170), .Y(n4070) );
  MUX2X1 U7205 ( .B(ram[639]), .A(ram[575]), .S(n4329), .Y(n4064) );
  MUX2X1 U7206 ( .B(ram[767]), .A(ram[703]), .S(n4329), .Y(n4063) );
  MUX2X1 U7207 ( .B(ram[895]), .A(ram[831]), .S(n4329), .Y(n4067) );
  MUX2X1 U7208 ( .B(ram[1023]), .A(ram[959]), .S(n4329), .Y(n4066) );
  MUX2X1 U7209 ( .B(n4065), .A(n4062), .S(n4173), .Y(n4069) );
  MUX2X1 U7210 ( .B(ram[1151]), .A(ram[1087]), .S(n4329), .Y(n4073) );
  MUX2X1 U7211 ( .B(ram[1279]), .A(ram[1215]), .S(n4329), .Y(n4072) );
  MUX2X1 U7212 ( .B(ram[1407]), .A(ram[1343]), .S(n4329), .Y(n4076) );
  MUX2X1 U7213 ( .B(ram[1535]), .A(ram[1471]), .S(n4329), .Y(n4075) );
  MUX2X1 U7214 ( .B(n4074), .A(n4071), .S(n4175), .Y(n4085) );
  MUX2X1 U7215 ( .B(ram[1663]), .A(ram[1599]), .S(n4329), .Y(n4079) );
  MUX2X1 U7216 ( .B(ram[1791]), .A(ram[1727]), .S(n4329), .Y(n4078) );
  MUX2X1 U7217 ( .B(ram[1919]), .A(ram[1855]), .S(n4329), .Y(n4082) );
  MUX2X1 U7218 ( .B(ram[2047]), .A(ram[1983]), .S(n4329), .Y(n4081) );
  MUX2X1 U7219 ( .B(n4080), .A(n4077), .S(n4168), .Y(n4084) );
  MUX2X1 U7220 ( .B(n4083), .A(n4068), .S(n4150), .Y(n4149) );
  MUX2X1 U7221 ( .B(n4340), .A(n4341), .S(n8416), .Y(n4339) );
  MUX2X1 U7222 ( .B(n4343), .A(n4344), .S(n8416), .Y(n4342) );
  MUX2X1 U7223 ( .B(n4346), .A(n4347), .S(n8416), .Y(n4345) );
  MUX2X1 U7224 ( .B(n4349), .A(n4350), .S(n8416), .Y(n4348) );
  MUX2X1 U7225 ( .B(n4352), .A(n4353), .S(n8389), .Y(n4351) );
  MUX2X1 U7226 ( .B(n4355), .A(n4356), .S(n8416), .Y(n4354) );
  MUX2X1 U7227 ( .B(n4358), .A(n4359), .S(n8416), .Y(n4357) );
  MUX2X1 U7228 ( .B(n4361), .A(n4362), .S(n8416), .Y(n4360) );
  MUX2X1 U7229 ( .B(n4364), .A(n4365), .S(n8416), .Y(n4363) );
  MUX2X1 U7230 ( .B(n4367), .A(n4368), .S(n8393), .Y(n4366) );
  MUX2X1 U7231 ( .B(n4370), .A(n4371), .S(n8417), .Y(n4369) );
  MUX2X1 U7232 ( .B(n4373), .A(n4374), .S(n8417), .Y(n4372) );
  MUX2X1 U7233 ( .B(n4376), .A(n4377), .S(n8417), .Y(n4375) );
  MUX2X1 U7234 ( .B(n4379), .A(n4380), .S(n8417), .Y(n4378) );
  MUX2X1 U7235 ( .B(n4382), .A(n4383), .S(n8393), .Y(n4381) );
  MUX2X1 U7236 ( .B(n4385), .A(n4386), .S(n8417), .Y(n4384) );
  MUX2X1 U7237 ( .B(n4388), .A(n4389), .S(n8417), .Y(n4387) );
  MUX2X1 U7238 ( .B(n4391), .A(n4392), .S(n8417), .Y(n4390) );
  MUX2X1 U7239 ( .B(n4394), .A(n4395), .S(n8417), .Y(n4393) );
  MUX2X1 U7240 ( .B(n4397), .A(n4398), .S(n8390), .Y(n4396) );
  MUX2X1 U7241 ( .B(n4400), .A(n4401), .S(n8417), .Y(n4399) );
  MUX2X1 U7242 ( .B(n4403), .A(n4404), .S(n8417), .Y(n4402) );
  MUX2X1 U7243 ( .B(n4406), .A(n4407), .S(n8417), .Y(n4405) );
  MUX2X1 U7244 ( .B(n4409), .A(n4410), .S(n8417), .Y(n4408) );
  MUX2X1 U7245 ( .B(n4412), .A(n4413), .S(n8392), .Y(n4411) );
  MUX2X1 U7246 ( .B(n4415), .A(n4416), .S(n8418), .Y(n4414) );
  MUX2X1 U7247 ( .B(n4418), .A(n4419), .S(n8418), .Y(n4417) );
  MUX2X1 U7248 ( .B(n4421), .A(n4422), .S(n8418), .Y(n4420) );
  MUX2X1 U7249 ( .B(n4424), .A(n4425), .S(n8418), .Y(n4423) );
  MUX2X1 U7250 ( .B(n4427), .A(n4428), .S(n8389), .Y(n4426) );
  MUX2X1 U7251 ( .B(n4430), .A(n4431), .S(n8418), .Y(n4429) );
  MUX2X1 U7252 ( .B(n4433), .A(n4434), .S(n8418), .Y(n4432) );
  MUX2X1 U7253 ( .B(n4436), .A(n4437), .S(n8418), .Y(n4435) );
  MUX2X1 U7254 ( .B(n4439), .A(n4440), .S(n8418), .Y(n4438) );
  MUX2X1 U7255 ( .B(n4442), .A(n4443), .S(n8394), .Y(n4441) );
  MUX2X1 U7256 ( .B(n4445), .A(n4446), .S(n8418), .Y(n4444) );
  MUX2X1 U7257 ( .B(n4448), .A(n4449), .S(n8418), .Y(n4447) );
  MUX2X1 U7258 ( .B(n4451), .A(n4452), .S(n8418), .Y(n4450) );
  MUX2X1 U7259 ( .B(n4454), .A(n4455), .S(n8418), .Y(n4453) );
  MUX2X1 U7260 ( .B(n4457), .A(n4458), .S(n8391), .Y(n4456) );
  MUX2X1 U7261 ( .B(n4460), .A(n4461), .S(n8419), .Y(n4459) );
  MUX2X1 U7262 ( .B(n4463), .A(n4464), .S(n8419), .Y(n4462) );
  MUX2X1 U7263 ( .B(n4466), .A(n4467), .S(n8419), .Y(n4465) );
  MUX2X1 U7264 ( .B(n4469), .A(n4470), .S(n8419), .Y(n4468) );
  MUX2X1 U7265 ( .B(n4472), .A(n4473), .S(n8390), .Y(n4471) );
  MUX2X1 U7266 ( .B(n4475), .A(n4476), .S(n8419), .Y(n4474) );
  MUX2X1 U7267 ( .B(n4478), .A(n4479), .S(n8419), .Y(n4477) );
  MUX2X1 U7268 ( .B(n4481), .A(n4482), .S(n8419), .Y(n4480) );
  MUX2X1 U7269 ( .B(n4484), .A(n4485), .S(n8419), .Y(n4483) );
  MUX2X1 U7270 ( .B(n4487), .A(n4488), .S(n8393), .Y(n4486) );
  MUX2X1 U7271 ( .B(n4490), .A(n4491), .S(n8419), .Y(n4489) );
  MUX2X1 U7272 ( .B(n4493), .A(n4494), .S(n8419), .Y(n4492) );
  MUX2X1 U7273 ( .B(n4496), .A(n4497), .S(n8419), .Y(n4495) );
  MUX2X1 U7274 ( .B(n4499), .A(n4500), .S(n8419), .Y(n4498) );
  MUX2X1 U7275 ( .B(n4502), .A(n4503), .S(n8389), .Y(n4501) );
  MUX2X1 U7276 ( .B(n4505), .A(n4506), .S(n8420), .Y(n4504) );
  MUX2X1 U7277 ( .B(n4509), .A(n4510), .S(n8420), .Y(n4507) );
  MUX2X1 U7278 ( .B(n4512), .A(n4513), .S(n8420), .Y(n4511) );
  MUX2X1 U7279 ( .B(n4515), .A(n4516), .S(n8420), .Y(n4514) );
  MUX2X1 U7280 ( .B(n4518), .A(n4519), .S(n8390), .Y(n4517) );
  MUX2X1 U7281 ( .B(n4521), .A(n4522), .S(n8420), .Y(n4520) );
  MUX2X1 U7282 ( .B(n4524), .A(n4525), .S(n8420), .Y(n4523) );
  MUX2X1 U7283 ( .B(n4527), .A(n4528), .S(n8420), .Y(n4526) );
  MUX2X1 U7284 ( .B(n4530), .A(n4531), .S(n8420), .Y(n4529) );
  MUX2X1 U7285 ( .B(n4533), .A(n4534), .S(n8392), .Y(n4532) );
  MUX2X1 U7286 ( .B(n4536), .A(n4537), .S(n8420), .Y(n4535) );
  MUX2X1 U7287 ( .B(n4539), .A(n4540), .S(n8420), .Y(n4538) );
  MUX2X1 U7288 ( .B(n4542), .A(n4543), .S(n8420), .Y(n4541) );
  MUX2X1 U7289 ( .B(n4545), .A(n4546), .S(n8420), .Y(n4544) );
  MUX2X1 U7290 ( .B(n4548), .A(n4549), .S(n8391), .Y(n4547) );
  MUX2X1 U7291 ( .B(n4551), .A(n4552), .S(n8421), .Y(n4550) );
  MUX2X1 U7292 ( .B(n4554), .A(n4555), .S(n8421), .Y(n4553) );
  MUX2X1 U7293 ( .B(n4557), .A(n4558), .S(n8421), .Y(n4556) );
  MUX2X1 U7294 ( .B(n4560), .A(n4561), .S(n8421), .Y(n4559) );
  MUX2X1 U7295 ( .B(n4563), .A(n4564), .S(n8391), .Y(n4562) );
  MUX2X1 U7296 ( .B(n4566), .A(n4567), .S(n8421), .Y(n4565) );
  MUX2X1 U7297 ( .B(n4569), .A(n4570), .S(n8421), .Y(n4568) );
  MUX2X1 U7298 ( .B(n4572), .A(n4573), .S(n8421), .Y(n4571) );
  MUX2X1 U7299 ( .B(n4575), .A(n4581), .S(n8421), .Y(n4574) );
  MUX2X1 U7300 ( .B(n4583), .A(n4584), .S(n8391), .Y(n4582) );
  MUX2X1 U7301 ( .B(n4586), .A(n4587), .S(n8421), .Y(n4585) );
  MUX2X1 U7302 ( .B(n4589), .A(n4590), .S(n8421), .Y(n4588) );
  MUX2X1 U7303 ( .B(n4592), .A(n4593), .S(n8421), .Y(n4591) );
  MUX2X1 U7304 ( .B(n4595), .A(n4596), .S(n8421), .Y(n4594) );
  MUX2X1 U7305 ( .B(n4598), .A(n4599), .S(n8392), .Y(n4597) );
  MUX2X1 U7306 ( .B(n4601), .A(n4602), .S(n8422), .Y(n4600) );
  MUX2X1 U7307 ( .B(n4604), .A(n4605), .S(n8422), .Y(n4603) );
  MUX2X1 U7308 ( .B(n4607), .A(n4608), .S(n8422), .Y(n4606) );
  MUX2X1 U7309 ( .B(n4610), .A(n4611), .S(n8422), .Y(n4609) );
  MUX2X1 U7310 ( .B(n4613), .A(n4614), .S(n8394), .Y(n4612) );
  MUX2X1 U7311 ( .B(n4616), .A(n4617), .S(n8422), .Y(n4615) );
  MUX2X1 U7312 ( .B(n4619), .A(n4620), .S(n8422), .Y(n4618) );
  MUX2X1 U7313 ( .B(n4622), .A(n4623), .S(n8422), .Y(n4621) );
  MUX2X1 U7314 ( .B(n4625), .A(n4626), .S(n8422), .Y(n4624) );
  MUX2X1 U7315 ( .B(n4628), .A(n4629), .S(n8392), .Y(n4627) );
  MUX2X1 U7316 ( .B(n4631), .A(n4632), .S(n8422), .Y(n4630) );
  MUX2X1 U7317 ( .B(n4634), .A(n4635), .S(n8422), .Y(n4633) );
  MUX2X1 U7318 ( .B(n4637), .A(n4638), .S(n8422), .Y(n4636) );
  MUX2X1 U7319 ( .B(n4640), .A(n4641), .S(n8422), .Y(n4639) );
  MUX2X1 U7320 ( .B(n4643), .A(n4644), .S(n8394), .Y(n4642) );
  MUX2X1 U7321 ( .B(n4646), .A(n4647), .S(n8423), .Y(n4645) );
  MUX2X1 U7322 ( .B(n4649), .A(n4650), .S(n8423), .Y(n4648) );
  MUX2X1 U7323 ( .B(n4652), .A(n4653), .S(n8423), .Y(n4651) );
  MUX2X1 U7324 ( .B(n4655), .A(n4656), .S(n8423), .Y(n4654) );
  MUX2X1 U7325 ( .B(n4658), .A(n4659), .S(n8389), .Y(n4657) );
  MUX2X1 U7326 ( .B(n4661), .A(n6717), .S(n8423), .Y(n4660) );
  MUX2X1 U7327 ( .B(n6719), .A(n6720), .S(n8423), .Y(n6718) );
  MUX2X1 U7328 ( .B(n6722), .A(n6723), .S(n8423), .Y(n6721) );
  MUX2X1 U7329 ( .B(n6725), .A(n6726), .S(n8423), .Y(n6724) );
  MUX2X1 U7330 ( .B(n6728), .A(n6729), .S(n8389), .Y(n6727) );
  MUX2X1 U7331 ( .B(n6731), .A(n6732), .S(n8423), .Y(n6730) );
  MUX2X1 U7332 ( .B(n6734), .A(n6735), .S(n8423), .Y(n6733) );
  MUX2X1 U7333 ( .B(n6737), .A(n6738), .S(n8423), .Y(n6736) );
  MUX2X1 U7334 ( .B(n6740), .A(n6741), .S(n8423), .Y(n6739) );
  MUX2X1 U7335 ( .B(n6743), .A(n6744), .S(n8389), .Y(n6742) );
  MUX2X1 U7336 ( .B(n6746), .A(n6747), .S(n8424), .Y(n6745) );
  MUX2X1 U7337 ( .B(n6749), .A(n6750), .S(n8424), .Y(n6748) );
  MUX2X1 U7338 ( .B(n6752), .A(n6753), .S(n8424), .Y(n6751) );
  MUX2X1 U7339 ( .B(n6755), .A(n6756), .S(n8424), .Y(n6754) );
  MUX2X1 U7340 ( .B(n6758), .A(n6759), .S(n8389), .Y(n6757) );
  MUX2X1 U7341 ( .B(n6761), .A(n6762), .S(n8424), .Y(n6760) );
  MUX2X1 U7342 ( .B(n6764), .A(n6765), .S(n8424), .Y(n6763) );
  MUX2X1 U7343 ( .B(n6767), .A(n6768), .S(n8424), .Y(n6766) );
  MUX2X1 U7344 ( .B(n6770), .A(n6771), .S(n8424), .Y(n6769) );
  MUX2X1 U7345 ( .B(n6773), .A(n6774), .S(n8389), .Y(n6772) );
  MUX2X1 U7346 ( .B(n6776), .A(n6777), .S(n8424), .Y(n6775) );
  MUX2X1 U7347 ( .B(n6779), .A(n6780), .S(n8424), .Y(n6778) );
  MUX2X1 U7348 ( .B(n6782), .A(n6783), .S(n8424), .Y(n6781) );
  MUX2X1 U7349 ( .B(n6785), .A(n6786), .S(n8424), .Y(n6784) );
  MUX2X1 U7350 ( .B(n6788), .A(n6789), .S(n8389), .Y(n6787) );
  MUX2X1 U7351 ( .B(n6791), .A(n6792), .S(n8425), .Y(n6790) );
  MUX2X1 U7352 ( .B(n6794), .A(n6795), .S(n8425), .Y(n6793) );
  MUX2X1 U7353 ( .B(n6797), .A(n6798), .S(n8425), .Y(n6796) );
  MUX2X1 U7354 ( .B(n6800), .A(n6801), .S(n8425), .Y(n6799) );
  MUX2X1 U7355 ( .B(n6803), .A(n6804), .S(n8389), .Y(n6802) );
  MUX2X1 U7356 ( .B(n6806), .A(n6807), .S(n8425), .Y(n6805) );
  MUX2X1 U7357 ( .B(n6809), .A(n6810), .S(n8425), .Y(n6808) );
  MUX2X1 U7358 ( .B(n6812), .A(n6813), .S(n8425), .Y(n6811) );
  MUX2X1 U7359 ( .B(n6815), .A(n6816), .S(n8425), .Y(n6814) );
  MUX2X1 U7360 ( .B(n6818), .A(n6819), .S(n8389), .Y(n6817) );
  MUX2X1 U7361 ( .B(n6821), .A(n6822), .S(n8425), .Y(n6820) );
  MUX2X1 U7362 ( .B(n6824), .A(n6825), .S(n8425), .Y(n6823) );
  MUX2X1 U7363 ( .B(n6827), .A(n6828), .S(n8425), .Y(n6826) );
  MUX2X1 U7364 ( .B(n6830), .A(n6831), .S(n8425), .Y(n6829) );
  MUX2X1 U7365 ( .B(n6833), .A(n6834), .S(n8389), .Y(n6832) );
  MUX2X1 U7366 ( .B(n6836), .A(n6837), .S(n8426), .Y(n6835) );
  MUX2X1 U7367 ( .B(n6839), .A(n6840), .S(n8426), .Y(n6838) );
  MUX2X1 U7368 ( .B(n6842), .A(n6843), .S(n8426), .Y(n6841) );
  MUX2X1 U7369 ( .B(n6845), .A(n6846), .S(n8426), .Y(n6844) );
  MUX2X1 U7370 ( .B(n6848), .A(n6849), .S(n8389), .Y(n6847) );
  MUX2X1 U7371 ( .B(n6851), .A(n6852), .S(n8426), .Y(n6850) );
  MUX2X1 U7372 ( .B(n6854), .A(n6855), .S(n8426), .Y(n6853) );
  MUX2X1 U7373 ( .B(n6857), .A(n6858), .S(n8426), .Y(n6856) );
  MUX2X1 U7374 ( .B(n6860), .A(n6861), .S(n8426), .Y(n6859) );
  MUX2X1 U7375 ( .B(n6863), .A(n6864), .S(n8389), .Y(n6862) );
  MUX2X1 U7376 ( .B(n6866), .A(n6867), .S(n8426), .Y(n6865) );
  MUX2X1 U7377 ( .B(n6869), .A(n6870), .S(n8426), .Y(n6868) );
  MUX2X1 U7378 ( .B(n6872), .A(n6873), .S(n8426), .Y(n6871) );
  MUX2X1 U7379 ( .B(n6875), .A(n6876), .S(n8426), .Y(n6874) );
  MUX2X1 U7380 ( .B(n6878), .A(n6879), .S(n8389), .Y(n6877) );
  MUX2X1 U7381 ( .B(n6881), .A(n6882), .S(n8427), .Y(n6880) );
  MUX2X1 U7382 ( .B(n6884), .A(n6885), .S(n8427), .Y(n6883) );
  MUX2X1 U7383 ( .B(n6887), .A(n6888), .S(n8427), .Y(n6886) );
  MUX2X1 U7384 ( .B(n6890), .A(n6891), .S(n8427), .Y(n6889) );
  MUX2X1 U7385 ( .B(n6893), .A(n6894), .S(n8390), .Y(n6892) );
  MUX2X1 U7386 ( .B(n6896), .A(n6897), .S(n8427), .Y(n6895) );
  MUX2X1 U7387 ( .B(n6899), .A(n6900), .S(n8427), .Y(n6898) );
  MUX2X1 U7388 ( .B(n6902), .A(n6903), .S(n8427), .Y(n6901) );
  MUX2X1 U7389 ( .B(n6905), .A(n6906), .S(n8427), .Y(n6904) );
  MUX2X1 U7390 ( .B(n6908), .A(n6909), .S(n8394), .Y(n6907) );
  MUX2X1 U7391 ( .B(n6911), .A(n6912), .S(n8427), .Y(n6910) );
  MUX2X1 U7392 ( .B(n6914), .A(n6915), .S(n8427), .Y(n6913) );
  MUX2X1 U7393 ( .B(n6917), .A(n6918), .S(n8427), .Y(n6916) );
  MUX2X1 U7394 ( .B(n6920), .A(n6921), .S(n8427), .Y(n6919) );
  MUX2X1 U7395 ( .B(n6923), .A(n6924), .S(n8393), .Y(n6922) );
  MUX2X1 U7396 ( .B(n6926), .A(n6927), .S(n8428), .Y(n6925) );
  MUX2X1 U7397 ( .B(n6929), .A(n6930), .S(n8428), .Y(n6928) );
  MUX2X1 U7398 ( .B(n6932), .A(n6933), .S(n8428), .Y(n6931) );
  MUX2X1 U7399 ( .B(n6935), .A(n6936), .S(n8428), .Y(n6934) );
  MUX2X1 U7400 ( .B(n6938), .A(n6939), .S(n8390), .Y(n6937) );
  MUX2X1 U7401 ( .B(n6941), .A(n6942), .S(n8428), .Y(n6940) );
  MUX2X1 U7402 ( .B(n6944), .A(n6945), .S(n8428), .Y(n6943) );
  MUX2X1 U7403 ( .B(n6947), .A(n6948), .S(n8428), .Y(n6946) );
  MUX2X1 U7404 ( .B(n6950), .A(n6951), .S(n8428), .Y(n6949) );
  MUX2X1 U7405 ( .B(n6953), .A(n6954), .S(n8390), .Y(n6952) );
  MUX2X1 U7406 ( .B(n6956), .A(n6957), .S(n8428), .Y(n6955) );
  MUX2X1 U7407 ( .B(n6959), .A(n6960), .S(n8428), .Y(n6958) );
  MUX2X1 U7408 ( .B(n6962), .A(n6963), .S(n8428), .Y(n6961) );
  MUX2X1 U7409 ( .B(n6965), .A(n6966), .S(n8428), .Y(n6964) );
  MUX2X1 U7410 ( .B(n6968), .A(n6969), .S(n8391), .Y(n6967) );
  MUX2X1 U7411 ( .B(n6971), .A(n6972), .S(n8429), .Y(n6970) );
  MUX2X1 U7412 ( .B(n6974), .A(n6975), .S(n8429), .Y(n6973) );
  MUX2X1 U7413 ( .B(n6977), .A(n6978), .S(n8429), .Y(n6976) );
  MUX2X1 U7414 ( .B(n6980), .A(n6981), .S(n8429), .Y(n6979) );
  MUX2X1 U7415 ( .B(n6983), .A(n6984), .S(n8394), .Y(n6982) );
  MUX2X1 U7416 ( .B(n6986), .A(n6987), .S(n8429), .Y(n6985) );
  MUX2X1 U7417 ( .B(n6989), .A(n6990), .S(n8429), .Y(n6988) );
  MUX2X1 U7418 ( .B(n6992), .A(n6993), .S(n8429), .Y(n6991) );
  MUX2X1 U7419 ( .B(n6995), .A(n6996), .S(n8429), .Y(n6994) );
  MUX2X1 U7420 ( .B(n6998), .A(n6999), .S(n8389), .Y(n6997) );
  MUX2X1 U7421 ( .B(n7001), .A(n7002), .S(n8429), .Y(n7000) );
  MUX2X1 U7422 ( .B(n7004), .A(n7005), .S(n8429), .Y(n7003) );
  MUX2X1 U7423 ( .B(n7007), .A(n7008), .S(n8429), .Y(n7006) );
  MUX2X1 U7424 ( .B(n7010), .A(n7011), .S(n8429), .Y(n7009) );
  MUX2X1 U7425 ( .B(n7013), .A(n7014), .S(n8394), .Y(n7012) );
  MUX2X1 U7426 ( .B(n7016), .A(n7017), .S(n8430), .Y(n7015) );
  MUX2X1 U7427 ( .B(n7019), .A(n7020), .S(n8430), .Y(n7018) );
  MUX2X1 U7428 ( .B(n7022), .A(n7023), .S(n8430), .Y(n7021) );
  MUX2X1 U7429 ( .B(n7025), .A(n7026), .S(n8430), .Y(n7024) );
  MUX2X1 U7430 ( .B(n7028), .A(n7029), .S(n8393), .Y(n7027) );
  MUX2X1 U7431 ( .B(n7031), .A(n7032), .S(n8430), .Y(n7030) );
  MUX2X1 U7432 ( .B(n7034), .A(n7035), .S(n8430), .Y(n7033) );
  MUX2X1 U7433 ( .B(n7037), .A(n7038), .S(n8430), .Y(n7036) );
  MUX2X1 U7434 ( .B(n7040), .A(n7041), .S(n8430), .Y(n7039) );
  MUX2X1 U7435 ( .B(n7043), .A(n7044), .S(n8393), .Y(n7042) );
  MUX2X1 U7436 ( .B(n7046), .A(n7047), .S(n8430), .Y(n7045) );
  MUX2X1 U7437 ( .B(n7049), .A(n7050), .S(n8430), .Y(n7048) );
  MUX2X1 U7438 ( .B(n7052), .A(n7053), .S(n8430), .Y(n7051) );
  MUX2X1 U7439 ( .B(n7055), .A(n7056), .S(n8430), .Y(n7054) );
  MUX2X1 U7440 ( .B(n7058), .A(n7059), .S(n8392), .Y(n7057) );
  MUX2X1 U7441 ( .B(n7061), .A(n7062), .S(n8431), .Y(n7060) );
  MUX2X1 U7442 ( .B(n7064), .A(n7065), .S(n8431), .Y(n7063) );
  MUX2X1 U7443 ( .B(n7067), .A(n7068), .S(n8431), .Y(n7066) );
  MUX2X1 U7444 ( .B(n7070), .A(n7071), .S(n8431), .Y(n7069) );
  MUX2X1 U7445 ( .B(n7073), .A(n7074), .S(n8393), .Y(n7072) );
  MUX2X1 U7446 ( .B(n7076), .A(n7077), .S(n8431), .Y(n7075) );
  MUX2X1 U7447 ( .B(n7079), .A(n7080), .S(n8431), .Y(n7078) );
  MUX2X1 U7448 ( .B(n7082), .A(n7083), .S(n8431), .Y(n7081) );
  MUX2X1 U7449 ( .B(n7085), .A(n7086), .S(n8431), .Y(n7084) );
  MUX2X1 U7450 ( .B(n7088), .A(n7089), .S(n8389), .Y(n7087) );
  MUX2X1 U7451 ( .B(n7091), .A(n7092), .S(n8431), .Y(n7090) );
  MUX2X1 U7452 ( .B(n7094), .A(n7095), .S(n8431), .Y(n7093) );
  MUX2X1 U7453 ( .B(n7097), .A(n7098), .S(n8431), .Y(n7096) );
  MUX2X1 U7454 ( .B(n7100), .A(n7101), .S(n8431), .Y(n7099) );
  MUX2X1 U7455 ( .B(n7103), .A(n7104), .S(n8391), .Y(n7102) );
  MUX2X1 U7456 ( .B(n7106), .A(n7107), .S(n8432), .Y(n7105) );
  MUX2X1 U7457 ( .B(n7109), .A(n7110), .S(n8432), .Y(n7108) );
  MUX2X1 U7458 ( .B(n7112), .A(n7113), .S(n8432), .Y(n7111) );
  MUX2X1 U7459 ( .B(n7115), .A(n7116), .S(n8432), .Y(n7114) );
  MUX2X1 U7460 ( .B(n7118), .A(n7119), .S(n8394), .Y(n7117) );
  MUX2X1 U7461 ( .B(n7121), .A(n7122), .S(n8432), .Y(n7120) );
  MUX2X1 U7462 ( .B(n7124), .A(n7125), .S(n8432), .Y(n7123) );
  MUX2X1 U7463 ( .B(n7127), .A(n7128), .S(n8432), .Y(n7126) );
  MUX2X1 U7464 ( .B(n7130), .A(n7131), .S(n8432), .Y(n7129) );
  MUX2X1 U7465 ( .B(n7133), .A(n7134), .S(n8391), .Y(n7132) );
  MUX2X1 U7466 ( .B(n7136), .A(n7137), .S(n8432), .Y(n7135) );
  MUX2X1 U7467 ( .B(n7139), .A(n7140), .S(n8432), .Y(n7138) );
  MUX2X1 U7468 ( .B(n7142), .A(n7143), .S(n8432), .Y(n7141) );
  MUX2X1 U7469 ( .B(n7145), .A(n7146), .S(n8432), .Y(n7144) );
  MUX2X1 U7470 ( .B(n7148), .A(n7149), .S(n8392), .Y(n7147) );
  MUX2X1 U7471 ( .B(n7151), .A(n7152), .S(n8433), .Y(n7150) );
  MUX2X1 U7472 ( .B(n7154), .A(n7155), .S(n8433), .Y(n7153) );
  MUX2X1 U7473 ( .B(n7157), .A(n7158), .S(n8433), .Y(n7156) );
  MUX2X1 U7474 ( .B(n7160), .A(n7161), .S(n8433), .Y(n7159) );
  MUX2X1 U7475 ( .B(n7163), .A(n7164), .S(n8394), .Y(n7162) );
  MUX2X1 U7476 ( .B(n7166), .A(n7167), .S(n8433), .Y(n7165) );
  MUX2X1 U7477 ( .B(n7169), .A(n7170), .S(n8433), .Y(n7168) );
  MUX2X1 U7478 ( .B(n7172), .A(n7173), .S(n8433), .Y(n7171) );
  MUX2X1 U7479 ( .B(n7175), .A(n7176), .S(n8433), .Y(n7174) );
  MUX2X1 U7480 ( .B(n7178), .A(n7179), .S(n8391), .Y(n7177) );
  MUX2X1 U7481 ( .B(n7181), .A(n7182), .S(n8433), .Y(n7180) );
  MUX2X1 U7482 ( .B(n7184), .A(n7185), .S(n8433), .Y(n7183) );
  MUX2X1 U7483 ( .B(n7187), .A(n7188), .S(n8433), .Y(n7186) );
  MUX2X1 U7484 ( .B(n7190), .A(n7191), .S(n8433), .Y(n7189) );
  MUX2X1 U7485 ( .B(n7193), .A(n7194), .S(n8390), .Y(n7192) );
  MUX2X1 U7486 ( .B(n7196), .A(n7197), .S(n8434), .Y(n7195) );
  MUX2X1 U7487 ( .B(n7199), .A(n7200), .S(n8434), .Y(n7198) );
  MUX2X1 U7488 ( .B(n7202), .A(n7203), .S(n8434), .Y(n7201) );
  MUX2X1 U7489 ( .B(n7205), .A(n7206), .S(n8434), .Y(n7204) );
  MUX2X1 U7490 ( .B(n7208), .A(n7209), .S(n8391), .Y(n7207) );
  MUX2X1 U7491 ( .B(n7211), .A(n7212), .S(n8434), .Y(n7210) );
  MUX2X1 U7492 ( .B(n7214), .A(n7215), .S(n8434), .Y(n7213) );
  MUX2X1 U7493 ( .B(n7217), .A(n7218), .S(n8434), .Y(n7216) );
  MUX2X1 U7494 ( .B(n7220), .A(n7221), .S(n8434), .Y(n7219) );
  MUX2X1 U7495 ( .B(n7223), .A(n7224), .S(n8392), .Y(n7222) );
  MUX2X1 U7496 ( .B(n7226), .A(n7227), .S(n8434), .Y(n7225) );
  MUX2X1 U7497 ( .B(n7229), .A(n7230), .S(n8434), .Y(n7228) );
  MUX2X1 U7498 ( .B(n7232), .A(n7233), .S(n8434), .Y(n7231) );
  MUX2X1 U7499 ( .B(n7235), .A(n7236), .S(n8434), .Y(n7234) );
  MUX2X1 U7500 ( .B(n7238), .A(n7239), .S(n8392), .Y(n7237) );
  MUX2X1 U7501 ( .B(n7241), .A(n7242), .S(n8435), .Y(n7240) );
  MUX2X1 U7502 ( .B(n7244), .A(n7245), .S(n8435), .Y(n7243) );
  MUX2X1 U7503 ( .B(n7247), .A(n7248), .S(n8435), .Y(n7246) );
  MUX2X1 U7504 ( .B(n7250), .A(n7251), .S(n8435), .Y(n7249) );
  MUX2X1 U7505 ( .B(n7253), .A(n7254), .S(n8390), .Y(n7252) );
  MUX2X1 U7506 ( .B(n7256), .A(n7257), .S(n8435), .Y(n7255) );
  MUX2X1 U7507 ( .B(n7259), .A(n7260), .S(n8435), .Y(n7258) );
  MUX2X1 U7508 ( .B(n7262), .A(n7263), .S(n8435), .Y(n7261) );
  MUX2X1 U7509 ( .B(n7265), .A(n7266), .S(n8435), .Y(n7264) );
  MUX2X1 U7510 ( .B(n7268), .A(n7269), .S(n8390), .Y(n7267) );
  MUX2X1 U7511 ( .B(n7271), .A(n7272), .S(n8435), .Y(n7270) );
  MUX2X1 U7512 ( .B(n7274), .A(n7275), .S(n8435), .Y(n7273) );
  MUX2X1 U7513 ( .B(n7277), .A(n7278), .S(n8435), .Y(n7276) );
  MUX2X1 U7514 ( .B(n7280), .A(n7281), .S(n8435), .Y(n7279) );
  MUX2X1 U7515 ( .B(n7283), .A(n7284), .S(n8390), .Y(n7282) );
  MUX2X1 U7516 ( .B(n7286), .A(n7287), .S(n8436), .Y(n7285) );
  MUX2X1 U7517 ( .B(n7289), .A(n7290), .S(n8436), .Y(n7288) );
  MUX2X1 U7518 ( .B(n7292), .A(n7293), .S(n8436), .Y(n7291) );
  MUX2X1 U7519 ( .B(n7295), .A(n7296), .S(n8436), .Y(n7294) );
  MUX2X1 U7520 ( .B(n7298), .A(n7299), .S(n8390), .Y(n7297) );
  MUX2X1 U7521 ( .B(n7301), .A(n7302), .S(n8436), .Y(n7300) );
  MUX2X1 U7522 ( .B(n7304), .A(n7305), .S(n8436), .Y(n7303) );
  MUX2X1 U7523 ( .B(n7307), .A(n7308), .S(n8436), .Y(n7306) );
  MUX2X1 U7524 ( .B(n7310), .A(n7311), .S(n8436), .Y(n7309) );
  MUX2X1 U7525 ( .B(n7313), .A(n7314), .S(n8390), .Y(n7312) );
  MUX2X1 U7526 ( .B(n7316), .A(n7317), .S(n8436), .Y(n7315) );
  MUX2X1 U7527 ( .B(n7319), .A(n7320), .S(n8436), .Y(n7318) );
  MUX2X1 U7528 ( .B(n7322), .A(n7323), .S(n8436), .Y(n7321) );
  MUX2X1 U7529 ( .B(n7325), .A(n7326), .S(n8436), .Y(n7324) );
  MUX2X1 U7530 ( .B(n7328), .A(n7329), .S(n8390), .Y(n7327) );
  MUX2X1 U7531 ( .B(n7331), .A(n7332), .S(n8437), .Y(n7330) );
  MUX2X1 U7532 ( .B(n7334), .A(n7335), .S(n8437), .Y(n7333) );
  MUX2X1 U7533 ( .B(n7337), .A(n7338), .S(n8437), .Y(n7336) );
  MUX2X1 U7534 ( .B(n7340), .A(n7341), .S(n8437), .Y(n7339) );
  MUX2X1 U7535 ( .B(n7343), .A(n7344), .S(n8390), .Y(n7342) );
  MUX2X1 U7536 ( .B(n7346), .A(n7347), .S(n8437), .Y(n7345) );
  MUX2X1 U7537 ( .B(n7349), .A(n7350), .S(n8437), .Y(n7348) );
  MUX2X1 U7538 ( .B(n7352), .A(n7353), .S(n8437), .Y(n7351) );
  MUX2X1 U7539 ( .B(n7355), .A(n7356), .S(n8437), .Y(n7354) );
  MUX2X1 U7540 ( .B(n7358), .A(n7359), .S(n8390), .Y(n7357) );
  MUX2X1 U7541 ( .B(n7361), .A(n7362), .S(n8437), .Y(n7360) );
  MUX2X1 U7542 ( .B(n7364), .A(n7365), .S(n8437), .Y(n7363) );
  MUX2X1 U7543 ( .B(n7367), .A(n7368), .S(n8437), .Y(n7366) );
  MUX2X1 U7544 ( .B(n7370), .A(n7371), .S(n8437), .Y(n7369) );
  MUX2X1 U7545 ( .B(n7373), .A(n7374), .S(n8390), .Y(n7372) );
  MUX2X1 U7546 ( .B(n7376), .A(n7377), .S(n8438), .Y(n7375) );
  MUX2X1 U7547 ( .B(n7379), .A(n7380), .S(n8438), .Y(n7378) );
  MUX2X1 U7548 ( .B(n7382), .A(n7383), .S(n8438), .Y(n7381) );
  MUX2X1 U7549 ( .B(n7385), .A(n7386), .S(n8438), .Y(n7384) );
  MUX2X1 U7550 ( .B(n7388), .A(n7389), .S(n8390), .Y(n7387) );
  MUX2X1 U7551 ( .B(n7391), .A(n7392), .S(n8438), .Y(n7390) );
  MUX2X1 U7552 ( .B(n7394), .A(n7395), .S(n8438), .Y(n7393) );
  MUX2X1 U7553 ( .B(n7397), .A(n7398), .S(n8438), .Y(n7396) );
  MUX2X1 U7554 ( .B(n7400), .A(n7401), .S(n8438), .Y(n7399) );
  MUX2X1 U7555 ( .B(n7403), .A(n7404), .S(n8390), .Y(n7402) );
  MUX2X1 U7556 ( .B(n7406), .A(n7407), .S(n8438), .Y(n7405) );
  MUX2X1 U7557 ( .B(n7409), .A(n7410), .S(n8438), .Y(n7408) );
  MUX2X1 U7558 ( .B(n7412), .A(n7413), .S(n8438), .Y(n7411) );
  MUX2X1 U7559 ( .B(n7415), .A(n7416), .S(n8438), .Y(n7414) );
  MUX2X1 U7560 ( .B(n7418), .A(n7419), .S(n8390), .Y(n7417) );
  MUX2X1 U7561 ( .B(n7421), .A(n7422), .S(n8439), .Y(n7420) );
  MUX2X1 U7562 ( .B(n7424), .A(n7425), .S(n8439), .Y(n7423) );
  MUX2X1 U7563 ( .B(n7427), .A(n7428), .S(n8439), .Y(n7426) );
  MUX2X1 U7564 ( .B(n7430), .A(n7431), .S(n8439), .Y(n7429) );
  MUX2X1 U7565 ( .B(n7433), .A(n7434), .S(n8391), .Y(n7432) );
  MUX2X1 U7566 ( .B(n7436), .A(n7437), .S(n8439), .Y(n7435) );
  MUX2X1 U7567 ( .B(n7439), .A(n7440), .S(n8439), .Y(n7438) );
  MUX2X1 U7568 ( .B(n7442), .A(n7443), .S(n8439), .Y(n7441) );
  MUX2X1 U7569 ( .B(n7445), .A(n7446), .S(n8439), .Y(n7444) );
  MUX2X1 U7570 ( .B(n7448), .A(n7449), .S(n8391), .Y(n7447) );
  MUX2X1 U7571 ( .B(n7451), .A(n7452), .S(n8439), .Y(n7450) );
  MUX2X1 U7572 ( .B(n7454), .A(n7455), .S(n8439), .Y(n7453) );
  MUX2X1 U7573 ( .B(n7457), .A(n7458), .S(n8439), .Y(n7456) );
  MUX2X1 U7574 ( .B(n7460), .A(n7461), .S(n8439), .Y(n7459) );
  MUX2X1 U7575 ( .B(n7463), .A(n7464), .S(n8391), .Y(n7462) );
  MUX2X1 U7576 ( .B(n7466), .A(n7467), .S(n8440), .Y(n7465) );
  MUX2X1 U7577 ( .B(n7469), .A(n7470), .S(n8440), .Y(n7468) );
  MUX2X1 U7578 ( .B(n7472), .A(n7473), .S(n8440), .Y(n7471) );
  MUX2X1 U7579 ( .B(n7475), .A(n7476), .S(n8440), .Y(n7474) );
  MUX2X1 U7580 ( .B(n7478), .A(n7479), .S(n8391), .Y(n7477) );
  MUX2X1 U7581 ( .B(n7481), .A(n7482), .S(n8440), .Y(n7480) );
  MUX2X1 U7582 ( .B(n7484), .A(n7485), .S(n8440), .Y(n7483) );
  MUX2X1 U7583 ( .B(n7487), .A(n7488), .S(n8440), .Y(n7486) );
  MUX2X1 U7584 ( .B(n7490), .A(n7491), .S(n8440), .Y(n7489) );
  MUX2X1 U7585 ( .B(n7493), .A(n7494), .S(n8391), .Y(n7492) );
  MUX2X1 U7586 ( .B(n7496), .A(n7497), .S(n8440), .Y(n7495) );
  MUX2X1 U7587 ( .B(n7499), .A(n7500), .S(n8440), .Y(n7498) );
  MUX2X1 U7588 ( .B(n7502), .A(n7503), .S(n8440), .Y(n7501) );
  MUX2X1 U7589 ( .B(n7505), .A(n7506), .S(n8440), .Y(n7504) );
  MUX2X1 U7590 ( .B(n7508), .A(n7509), .S(n8391), .Y(n7507) );
  MUX2X1 U7591 ( .B(n7511), .A(n7512), .S(n8441), .Y(n7510) );
  MUX2X1 U7592 ( .B(n7514), .A(n7515), .S(n8441), .Y(n7513) );
  MUX2X1 U7593 ( .B(n7517), .A(n7518), .S(n8441), .Y(n7516) );
  MUX2X1 U7594 ( .B(n7520), .A(n7521), .S(n8441), .Y(n7519) );
  MUX2X1 U7595 ( .B(n7523), .A(n7524), .S(n8391), .Y(n7522) );
  MUX2X1 U7596 ( .B(n7526), .A(n7527), .S(n8441), .Y(n7525) );
  MUX2X1 U7597 ( .B(n7529), .A(n7530), .S(n8441), .Y(n7528) );
  MUX2X1 U7598 ( .B(n7532), .A(n7533), .S(n8441), .Y(n7531) );
  MUX2X1 U7599 ( .B(n7535), .A(n7536), .S(n8441), .Y(n7534) );
  MUX2X1 U7600 ( .B(n7538), .A(n7539), .S(n8391), .Y(n7537) );
  MUX2X1 U7601 ( .B(n7541), .A(n7542), .S(n8441), .Y(n7540) );
  MUX2X1 U7602 ( .B(n7544), .A(n7545), .S(n8441), .Y(n7543) );
  MUX2X1 U7603 ( .B(n7547), .A(n7548), .S(n8441), .Y(n7546) );
  MUX2X1 U7604 ( .B(n7550), .A(n7551), .S(n8441), .Y(n7549) );
  MUX2X1 U7605 ( .B(n7553), .A(n7554), .S(n8391), .Y(n7552) );
  MUX2X1 U7606 ( .B(n7556), .A(n7557), .S(n8442), .Y(n7555) );
  MUX2X1 U7607 ( .B(n7559), .A(n7560), .S(n8442), .Y(n7558) );
  MUX2X1 U7608 ( .B(n7562), .A(n7563), .S(n8442), .Y(n7561) );
  MUX2X1 U7609 ( .B(n7565), .A(n7566), .S(n8442), .Y(n7564) );
  MUX2X1 U7610 ( .B(n7568), .A(n7569), .S(n8391), .Y(n7567) );
  MUX2X1 U7611 ( .B(n7571), .A(n7572), .S(n8442), .Y(n7570) );
  MUX2X1 U7612 ( .B(n7574), .A(n7575), .S(n8442), .Y(n7573) );
  MUX2X1 U7613 ( .B(n7577), .A(n7578), .S(n8442), .Y(n7576) );
  MUX2X1 U7614 ( .B(n7580), .A(n7581), .S(n8442), .Y(n7579) );
  MUX2X1 U7615 ( .B(n7583), .A(n7584), .S(n8391), .Y(n7582) );
  MUX2X1 U7616 ( .B(n7586), .A(n7587), .S(n8442), .Y(n7585) );
  MUX2X1 U7617 ( .B(n7589), .A(n7590), .S(n8442), .Y(n7588) );
  MUX2X1 U7618 ( .B(n7592), .A(n7593), .S(n8442), .Y(n7591) );
  MUX2X1 U7619 ( .B(n7595), .A(n7596), .S(n8442), .Y(n7594) );
  MUX2X1 U7620 ( .B(n7598), .A(n7599), .S(n8391), .Y(n7597) );
  MUX2X1 U7621 ( .B(n7601), .A(n7602), .S(n8443), .Y(n7600) );
  MUX2X1 U7622 ( .B(n7604), .A(n7605), .S(n8443), .Y(n7603) );
  MUX2X1 U7623 ( .B(n7607), .A(n7608), .S(n8443), .Y(n7606) );
  MUX2X1 U7624 ( .B(n7610), .A(n7611), .S(n8443), .Y(n7609) );
  MUX2X1 U7625 ( .B(n7613), .A(n7614), .S(n8392), .Y(n7612) );
  MUX2X1 U7626 ( .B(n7616), .A(n7617), .S(n8443), .Y(n7615) );
  MUX2X1 U7627 ( .B(n7619), .A(n7620), .S(n8443), .Y(n7618) );
  MUX2X1 U7628 ( .B(n7622), .A(n7623), .S(n8443), .Y(n7621) );
  MUX2X1 U7629 ( .B(n7625), .A(n7626), .S(n8443), .Y(n7624) );
  MUX2X1 U7630 ( .B(n7628), .A(n7629), .S(n8392), .Y(n7627) );
  MUX2X1 U7631 ( .B(n7631), .A(n7632), .S(n8443), .Y(n7630) );
  MUX2X1 U7632 ( .B(n7634), .A(n7635), .S(n8443), .Y(n7633) );
  MUX2X1 U7633 ( .B(n7637), .A(n7638), .S(n8443), .Y(n7636) );
  MUX2X1 U7634 ( .B(n7640), .A(n7641), .S(n8443), .Y(n7639) );
  MUX2X1 U7635 ( .B(n7643), .A(n7644), .S(n8392), .Y(n7642) );
  MUX2X1 U7636 ( .B(n7646), .A(n7647), .S(n8444), .Y(n7645) );
  MUX2X1 U7637 ( .B(n7649), .A(n7650), .S(n8444), .Y(n7648) );
  MUX2X1 U7638 ( .B(n7652), .A(n7653), .S(n8444), .Y(n7651) );
  MUX2X1 U7639 ( .B(n7655), .A(n7656), .S(n8444), .Y(n7654) );
  MUX2X1 U7640 ( .B(n7658), .A(n7659), .S(n8392), .Y(n7657) );
  MUX2X1 U7641 ( .B(n7661), .A(n7662), .S(n8444), .Y(n7660) );
  MUX2X1 U7642 ( .B(n7664), .A(n7665), .S(n8444), .Y(n7663) );
  MUX2X1 U7643 ( .B(n7667), .A(n7668), .S(n8444), .Y(n7666) );
  MUX2X1 U7644 ( .B(n7670), .A(n7671), .S(n8444), .Y(n7669) );
  MUX2X1 U7645 ( .B(n7673), .A(n7674), .S(n8392), .Y(n7672) );
  MUX2X1 U7646 ( .B(n7676), .A(n7677), .S(n8444), .Y(n7675) );
  MUX2X1 U7647 ( .B(n7679), .A(n7680), .S(n8444), .Y(n7678) );
  MUX2X1 U7648 ( .B(n7682), .A(n7683), .S(n8444), .Y(n7681) );
  MUX2X1 U7649 ( .B(n7685), .A(n7686), .S(n8444), .Y(n7684) );
  MUX2X1 U7650 ( .B(n7688), .A(n7689), .S(n8392), .Y(n7687) );
  MUX2X1 U7651 ( .B(n7691), .A(n7692), .S(n8445), .Y(n7690) );
  MUX2X1 U7652 ( .B(n7694), .A(n7695), .S(n8445), .Y(n7693) );
  MUX2X1 U7653 ( .B(n7697), .A(n7698), .S(n8445), .Y(n7696) );
  MUX2X1 U7654 ( .B(n7700), .A(n7701), .S(n8445), .Y(n7699) );
  MUX2X1 U7655 ( .B(n7703), .A(n7704), .S(n8392), .Y(n7702) );
  MUX2X1 U7656 ( .B(n7706), .A(n7707), .S(n8445), .Y(n7705) );
  MUX2X1 U7657 ( .B(n7709), .A(n7710), .S(n8445), .Y(n7708) );
  MUX2X1 U7658 ( .B(n7712), .A(n7713), .S(n8445), .Y(n7711) );
  MUX2X1 U7659 ( .B(n7715), .A(n7716), .S(n8445), .Y(n7714) );
  MUX2X1 U7660 ( .B(n7718), .A(n7719), .S(n8392), .Y(n7717) );
  MUX2X1 U7661 ( .B(n7721), .A(n7722), .S(n8445), .Y(n7720) );
  MUX2X1 U7662 ( .B(n7724), .A(n7725), .S(n8445), .Y(n7723) );
  MUX2X1 U7663 ( .B(n7727), .A(n7728), .S(n8445), .Y(n7726) );
  MUX2X1 U7664 ( .B(n7730), .A(n7731), .S(n8445), .Y(n7729) );
  MUX2X1 U7665 ( .B(n7733), .A(n7734), .S(n8392), .Y(n7732) );
  MUX2X1 U7666 ( .B(n7736), .A(n7737), .S(n8446), .Y(n7735) );
  MUX2X1 U7667 ( .B(n7739), .A(n7740), .S(n8446), .Y(n7738) );
  MUX2X1 U7668 ( .B(n7742), .A(n7743), .S(n8446), .Y(n7741) );
  MUX2X1 U7669 ( .B(n7745), .A(n7746), .S(n8446), .Y(n7744) );
  MUX2X1 U7670 ( .B(n7748), .A(n7749), .S(n8392), .Y(n7747) );
  MUX2X1 U7671 ( .B(n7751), .A(n7752), .S(n8446), .Y(n7750) );
  MUX2X1 U7672 ( .B(n7754), .A(n7755), .S(n8446), .Y(n7753) );
  MUX2X1 U7673 ( .B(n7757), .A(n7758), .S(n8446), .Y(n7756) );
  MUX2X1 U7674 ( .B(n7760), .A(n7761), .S(n8446), .Y(n7759) );
  MUX2X1 U7675 ( .B(n7763), .A(n7764), .S(n8392), .Y(n7762) );
  MUX2X1 U7676 ( .B(n7766), .A(n7767), .S(n8446), .Y(n7765) );
  MUX2X1 U7677 ( .B(n7769), .A(n7770), .S(n8446), .Y(n7768) );
  MUX2X1 U7678 ( .B(n7772), .A(n7773), .S(n8446), .Y(n7771) );
  MUX2X1 U7679 ( .B(n7775), .A(n7776), .S(n8446), .Y(n7774) );
  MUX2X1 U7680 ( .B(n7778), .A(n7779), .S(n8392), .Y(n7777) );
  MUX2X1 U7681 ( .B(n7781), .A(n7782), .S(n8447), .Y(n7780) );
  MUX2X1 U7682 ( .B(n7784), .A(n7785), .S(n8447), .Y(n7783) );
  MUX2X1 U7683 ( .B(n7787), .A(n7788), .S(n8447), .Y(n7786) );
  MUX2X1 U7684 ( .B(n7790), .A(n7791), .S(n8447), .Y(n7789) );
  MUX2X1 U7685 ( .B(n7793), .A(n7794), .S(n8393), .Y(n7792) );
  MUX2X1 U7686 ( .B(n7796), .A(n7797), .S(n8447), .Y(n7795) );
  MUX2X1 U7687 ( .B(n7799), .A(n7800), .S(n8447), .Y(n7798) );
  MUX2X1 U7688 ( .B(n7802), .A(n7803), .S(n8447), .Y(n7801) );
  MUX2X1 U7689 ( .B(n7805), .A(n7806), .S(n8447), .Y(n7804) );
  MUX2X1 U7690 ( .B(n7808), .A(n7809), .S(n8393), .Y(n7807) );
  MUX2X1 U7691 ( .B(n7811), .A(n7812), .S(n8447), .Y(n7810) );
  MUX2X1 U7692 ( .B(n7814), .A(n7815), .S(n8447), .Y(n7813) );
  MUX2X1 U7693 ( .B(n7817), .A(n7818), .S(n8447), .Y(n7816) );
  MUX2X1 U7694 ( .B(n7820), .A(n7821), .S(n8447), .Y(n7819) );
  MUX2X1 U7695 ( .B(n7823), .A(n7824), .S(n8393), .Y(n7822) );
  MUX2X1 U7696 ( .B(n7826), .A(n7827), .S(n8448), .Y(n7825) );
  MUX2X1 U7697 ( .B(n7829), .A(n7830), .S(n8448), .Y(n7828) );
  MUX2X1 U7698 ( .B(n7832), .A(n7833), .S(n8448), .Y(n7831) );
  MUX2X1 U7699 ( .B(n7835), .A(n7836), .S(n8448), .Y(n7834) );
  MUX2X1 U7700 ( .B(n7838), .A(n7839), .S(n8393), .Y(n7837) );
  MUX2X1 U7701 ( .B(n7841), .A(n7842), .S(n8448), .Y(n7840) );
  MUX2X1 U7702 ( .B(n7844), .A(n7845), .S(n8448), .Y(n7843) );
  MUX2X1 U7703 ( .B(n7847), .A(n7848), .S(n8448), .Y(n7846) );
  MUX2X1 U7704 ( .B(n7850), .A(n7851), .S(n8448), .Y(n7849) );
  MUX2X1 U7705 ( .B(n7853), .A(n7854), .S(n8393), .Y(n7852) );
  MUX2X1 U7706 ( .B(n7856), .A(n7857), .S(n8448), .Y(n7855) );
  MUX2X1 U7707 ( .B(n7859), .A(n7860), .S(n8448), .Y(n7858) );
  MUX2X1 U7708 ( .B(n7862), .A(n7863), .S(n8448), .Y(n7861) );
  MUX2X1 U7709 ( .B(n7865), .A(n7866), .S(n8448), .Y(n7864) );
  MUX2X1 U7710 ( .B(n7868), .A(n7869), .S(n8393), .Y(n7867) );
  MUX2X1 U7711 ( .B(n7871), .A(n7872), .S(n8449), .Y(n7870) );
  MUX2X1 U7712 ( .B(n7874), .A(n7875), .S(n8449), .Y(n7873) );
  MUX2X1 U7713 ( .B(n7877), .A(n7878), .S(n8449), .Y(n7876) );
  MUX2X1 U7714 ( .B(n7880), .A(n7881), .S(n8449), .Y(n7879) );
  MUX2X1 U7715 ( .B(n7883), .A(n7884), .S(n8393), .Y(n7882) );
  MUX2X1 U7716 ( .B(n7886), .A(n7887), .S(n8449), .Y(n7885) );
  MUX2X1 U7717 ( .B(n7889), .A(n7890), .S(n8449), .Y(n7888) );
  MUX2X1 U7718 ( .B(n7892), .A(n7893), .S(n8449), .Y(n7891) );
  MUX2X1 U7719 ( .B(n7895), .A(n7896), .S(n8449), .Y(n7894) );
  MUX2X1 U7720 ( .B(n7898), .A(n7899), .S(n8393), .Y(n7897) );
  MUX2X1 U7721 ( .B(n7901), .A(n7902), .S(n8449), .Y(n7900) );
  MUX2X1 U7722 ( .B(n7904), .A(n7905), .S(n8449), .Y(n7903) );
  MUX2X1 U7723 ( .B(n7907), .A(n7908), .S(n8449), .Y(n7906) );
  MUX2X1 U7724 ( .B(n7910), .A(n7911), .S(n8449), .Y(n7909) );
  MUX2X1 U7725 ( .B(n7913), .A(n7914), .S(n8393), .Y(n7912) );
  MUX2X1 U7726 ( .B(n7916), .A(n7917), .S(n8450), .Y(n7915) );
  MUX2X1 U7727 ( .B(n7919), .A(n7920), .S(n8450), .Y(n7918) );
  MUX2X1 U7728 ( .B(n7922), .A(n7923), .S(n8450), .Y(n7921) );
  MUX2X1 U7729 ( .B(n7925), .A(n7926), .S(n8450), .Y(n7924) );
  MUX2X1 U7730 ( .B(n7928), .A(n7929), .S(n8393), .Y(n7927) );
  MUX2X1 U7731 ( .B(n7931), .A(n7932), .S(n8450), .Y(n7930) );
  MUX2X1 U7732 ( .B(n7934), .A(n7935), .S(n8450), .Y(n7933) );
  MUX2X1 U7733 ( .B(n7937), .A(n7938), .S(n8450), .Y(n7936) );
  MUX2X1 U7734 ( .B(n7940), .A(n7941), .S(n8450), .Y(n7939) );
  MUX2X1 U7735 ( .B(n7943), .A(n7944), .S(n8393), .Y(n7942) );
  MUX2X1 U7736 ( .B(n7946), .A(n7947), .S(n8450), .Y(n7945) );
  MUX2X1 U7737 ( .B(n7949), .A(n7950), .S(n8450), .Y(n7948) );
  MUX2X1 U7738 ( .B(n7952), .A(n7953), .S(n8450), .Y(n7951) );
  MUX2X1 U7739 ( .B(n7955), .A(n7956), .S(n8450), .Y(n7954) );
  MUX2X1 U7740 ( .B(n7958), .A(n7959), .S(n8393), .Y(n7957) );
  MUX2X1 U7741 ( .B(n7961), .A(n7962), .S(n8451), .Y(n7960) );
  MUX2X1 U7742 ( .B(n7964), .A(n7965), .S(n8451), .Y(n7963) );
  MUX2X1 U7743 ( .B(n7967), .A(n7968), .S(n8451), .Y(n7966) );
  MUX2X1 U7744 ( .B(n7970), .A(n7971), .S(n8451), .Y(n7969) );
  MUX2X1 U7745 ( .B(n7973), .A(n7974), .S(n8394), .Y(n7972) );
  MUX2X1 U7746 ( .B(n7976), .A(n7977), .S(n8451), .Y(n7975) );
  MUX2X1 U7747 ( .B(n7979), .A(n7980), .S(n8451), .Y(n7978) );
  MUX2X1 U7748 ( .B(n7982), .A(n7983), .S(n8451), .Y(n7981) );
  MUX2X1 U7749 ( .B(n7985), .A(n7986), .S(n8451), .Y(n7984) );
  MUX2X1 U7750 ( .B(n7988), .A(n7989), .S(n8394), .Y(n7987) );
  MUX2X1 U7751 ( .B(n7991), .A(n7992), .S(n8451), .Y(n7990) );
  MUX2X1 U7752 ( .B(n7994), .A(n7995), .S(n8451), .Y(n7993) );
  MUX2X1 U7753 ( .B(n7997), .A(n7998), .S(n8451), .Y(n7996) );
  MUX2X1 U7754 ( .B(n8000), .A(n8001), .S(n8451), .Y(n7999) );
  MUX2X1 U7755 ( .B(n8003), .A(n8004), .S(n8394), .Y(n8002) );
  MUX2X1 U7756 ( .B(n8006), .A(n8007), .S(n8452), .Y(n8005) );
  MUX2X1 U7757 ( .B(n8009), .A(n8010), .S(n8452), .Y(n8008) );
  MUX2X1 U7758 ( .B(n8012), .A(n8013), .S(n8452), .Y(n8011) );
  MUX2X1 U7759 ( .B(n8015), .A(n8016), .S(n8452), .Y(n8014) );
  MUX2X1 U7760 ( .B(n8018), .A(n8019), .S(n8394), .Y(n8017) );
  MUX2X1 U7761 ( .B(n8021), .A(n8022), .S(n8452), .Y(n8020) );
  MUX2X1 U7762 ( .B(n8024), .A(n8025), .S(n8452), .Y(n8023) );
  MUX2X1 U7763 ( .B(n8027), .A(n8028), .S(n8452), .Y(n8026) );
  MUX2X1 U7764 ( .B(n8030), .A(n8031), .S(n8452), .Y(n8029) );
  MUX2X1 U7765 ( .B(n8033), .A(n8034), .S(n8394), .Y(n8032) );
  MUX2X1 U7766 ( .B(n8036), .A(n8037), .S(n8452), .Y(n8035) );
  MUX2X1 U7767 ( .B(n8039), .A(n8040), .S(n8452), .Y(n8038) );
  MUX2X1 U7768 ( .B(n8042), .A(n8043), .S(n8452), .Y(n8041) );
  MUX2X1 U7769 ( .B(n8045), .A(n8046), .S(n8452), .Y(n8044) );
  MUX2X1 U7770 ( .B(n8048), .A(n8049), .S(n8394), .Y(n8047) );
  MUX2X1 U7771 ( .B(n8051), .A(n8052), .S(n8453), .Y(n8050) );
  MUX2X1 U7772 ( .B(n8054), .A(n8055), .S(n8453), .Y(n8053) );
  MUX2X1 U7773 ( .B(n8057), .A(n8058), .S(n8453), .Y(n8056) );
  MUX2X1 U7774 ( .B(n8060), .A(n8061), .S(n8453), .Y(n8059) );
  MUX2X1 U7775 ( .B(n8063), .A(n8064), .S(n8394), .Y(n8062) );
  MUX2X1 U7776 ( .B(n8066), .A(n8067), .S(n8453), .Y(n8065) );
  MUX2X1 U7777 ( .B(n8069), .A(n8070), .S(n8453), .Y(n8068) );
  MUX2X1 U7778 ( .B(n8072), .A(n8073), .S(n8453), .Y(n8071) );
  MUX2X1 U7779 ( .B(n8075), .A(n8076), .S(n8453), .Y(n8074) );
  MUX2X1 U7780 ( .B(n8078), .A(n8079), .S(n8394), .Y(n8077) );
  MUX2X1 U7781 ( .B(n8081), .A(n8082), .S(n8453), .Y(n8080) );
  MUX2X1 U7782 ( .B(n8084), .A(n8085), .S(n8453), .Y(n8083) );
  MUX2X1 U7783 ( .B(n8087), .A(n8088), .S(n8453), .Y(n8086) );
  MUX2X1 U7784 ( .B(n8090), .A(n8091), .S(n8453), .Y(n8089) );
  MUX2X1 U7785 ( .B(n8093), .A(n8094), .S(n8394), .Y(n8092) );
  MUX2X1 U7786 ( .B(n8096), .A(n8097), .S(n8454), .Y(n8095) );
  MUX2X1 U7787 ( .B(n8099), .A(n8100), .S(n8454), .Y(n8098) );
  MUX2X1 U7788 ( .B(n8102), .A(n8103), .S(n8454), .Y(n8101) );
  MUX2X1 U7789 ( .B(n8105), .A(n8106), .S(n8454), .Y(n8104) );
  MUX2X1 U7790 ( .B(n8108), .A(n8109), .S(n8394), .Y(n8107) );
  MUX2X1 U7791 ( .B(n8111), .A(n8112), .S(n8454), .Y(n8110) );
  MUX2X1 U7792 ( .B(n8114), .A(n8115), .S(n8454), .Y(n8113) );
  MUX2X1 U7793 ( .B(n8117), .A(n8118), .S(n8454), .Y(n8116) );
  MUX2X1 U7794 ( .B(n8120), .A(n8121), .S(n8454), .Y(n8119) );
  MUX2X1 U7795 ( .B(n8123), .A(n8124), .S(n8394), .Y(n8122) );
  MUX2X1 U7796 ( .B(n8126), .A(n8127), .S(n8454), .Y(n8125) );
  MUX2X1 U7797 ( .B(n8129), .A(n8130), .S(n8454), .Y(n8128) );
  MUX2X1 U7798 ( .B(n8132), .A(n8133), .S(n8454), .Y(n8131) );
  MUX2X1 U7799 ( .B(n8135), .A(n8136), .S(n8454), .Y(n8134) );
  MUX2X1 U7800 ( .B(n8138), .A(n8139), .S(n8394), .Y(n8137) );
  MUX2X1 U7801 ( .B(n8141), .A(n8142), .S(n8455), .Y(n8140) );
  MUX2X1 U7802 ( .B(n8144), .A(n8145), .S(n8455), .Y(n8143) );
  MUX2X1 U7803 ( .B(n8147), .A(n8148), .S(n8455), .Y(n8146) );
  MUX2X1 U7804 ( .B(n8150), .A(n8151), .S(n8455), .Y(n8149) );
  MUX2X1 U7805 ( .B(n8153), .A(n8154), .S(n8394), .Y(n8152) );
  MUX2X1 U7806 ( .B(n8156), .A(n8157), .S(n8455), .Y(n8155) );
  MUX2X1 U7807 ( .B(n8159), .A(n8160), .S(n8455), .Y(n8158) );
  MUX2X1 U7808 ( .B(n8162), .A(n8163), .S(n8455), .Y(n8161) );
  MUX2X1 U7809 ( .B(n8165), .A(n8166), .S(n8455), .Y(n8164) );
  MUX2X1 U7810 ( .B(n8168), .A(n8169), .S(n8391), .Y(n8167) );
  MUX2X1 U7811 ( .B(n8171), .A(n8172), .S(n8455), .Y(n8170) );
  MUX2X1 U7812 ( .B(n8174), .A(n8175), .S(n8455), .Y(n8173) );
  MUX2X1 U7813 ( .B(n8177), .A(n8178), .S(n8455), .Y(n8176) );
  MUX2X1 U7814 ( .B(n8180), .A(n8181), .S(n8455), .Y(n8179) );
  MUX2X1 U7815 ( .B(n8183), .A(n8184), .S(n8392), .Y(n8182) );
  MUX2X1 U7816 ( .B(n8186), .A(n8187), .S(n8456), .Y(n8185) );
  MUX2X1 U7817 ( .B(n8189), .A(n8190), .S(n8456), .Y(n8188) );
  MUX2X1 U7818 ( .B(n8192), .A(n8193), .S(n8456), .Y(n8191) );
  MUX2X1 U7819 ( .B(n8195), .A(n8196), .S(n8456), .Y(n8194) );
  MUX2X1 U7820 ( .B(n8198), .A(n8199), .S(n8389), .Y(n8197) );
  MUX2X1 U7821 ( .B(n8201), .A(n8202), .S(n8456), .Y(n8200) );
  MUX2X1 U7822 ( .B(n8204), .A(n8205), .S(n8456), .Y(n8203) );
  MUX2X1 U7823 ( .B(n8207), .A(n8208), .S(n8456), .Y(n8206) );
  MUX2X1 U7824 ( .B(n8210), .A(n8211), .S(n8456), .Y(n8209) );
  MUX2X1 U7825 ( .B(n8213), .A(n8214), .S(n8391), .Y(n8212) );
  MUX2X1 U7826 ( .B(n8216), .A(n8217), .S(n8456), .Y(n8215) );
  MUX2X1 U7827 ( .B(n8219), .A(n8220), .S(n8456), .Y(n8218) );
  MUX2X1 U7828 ( .B(n8222), .A(n8223), .S(n8456), .Y(n8221) );
  MUX2X1 U7829 ( .B(n8225), .A(n8226), .S(n8456), .Y(n8224) );
  MUX2X1 U7830 ( .B(n8228), .A(n8229), .S(n8394), .Y(n8227) );
  MUX2X1 U7831 ( .B(n8231), .A(n8232), .S(n8457), .Y(n8230) );
  MUX2X1 U7832 ( .B(n8234), .A(n8235), .S(n8457), .Y(n8233) );
  MUX2X1 U7833 ( .B(n8237), .A(n8238), .S(n8457), .Y(n8236) );
  MUX2X1 U7834 ( .B(n8240), .A(n8241), .S(n8457), .Y(n8239) );
  MUX2X1 U7835 ( .B(n8243), .A(n8244), .S(n8392), .Y(n8242) );
  MUX2X1 U7836 ( .B(n8246), .A(n8247), .S(n8457), .Y(n8245) );
  MUX2X1 U7837 ( .B(n8249), .A(n8250), .S(n8457), .Y(n8248) );
  MUX2X1 U7838 ( .B(n8252), .A(n8253), .S(n8457), .Y(n8251) );
  MUX2X1 U7839 ( .B(n8255), .A(n8256), .S(n8457), .Y(n8254) );
  MUX2X1 U7840 ( .B(n8258), .A(n8259), .S(n8394), .Y(n8257) );
  MUX2X1 U7841 ( .B(n8261), .A(n8262), .S(n8457), .Y(n8260) );
  MUX2X1 U7842 ( .B(n8264), .A(n8265), .S(n8457), .Y(n8263) );
  MUX2X1 U7843 ( .B(n8267), .A(n8268), .S(n8457), .Y(n8266) );
  MUX2X1 U7844 ( .B(n8270), .A(n8271), .S(n8457), .Y(n8269) );
  MUX2X1 U7845 ( .B(n8273), .A(n8274), .S(n8392), .Y(n8272) );
  MUX2X1 U7846 ( .B(n8276), .A(n8277), .S(n8458), .Y(n8275) );
  MUX2X1 U7847 ( .B(n8279), .A(n8280), .S(n8458), .Y(n8278) );
  MUX2X1 U7848 ( .B(n8282), .A(n8283), .S(n8458), .Y(n8281) );
  MUX2X1 U7849 ( .B(n8285), .A(n8286), .S(n8458), .Y(n8284) );
  MUX2X1 U7850 ( .B(n8288), .A(n8289), .S(n8389), .Y(n8287) );
  MUX2X1 U7851 ( .B(n8291), .A(n8292), .S(n8458), .Y(n8290) );
  MUX2X1 U7852 ( .B(n8294), .A(n8295), .S(n8458), .Y(n8293) );
  MUX2X1 U7853 ( .B(n8297), .A(n8298), .S(n8458), .Y(n8296) );
  MUX2X1 U7854 ( .B(n8300), .A(n8301), .S(n8458), .Y(n8299) );
  MUX2X1 U7855 ( .B(n8303), .A(n8304), .S(n8394), .Y(n8302) );
  MUX2X1 U7856 ( .B(n8306), .A(n8307), .S(n8458), .Y(n8305) );
  MUX2X1 U7857 ( .B(n8309), .A(n8310), .S(n8458), .Y(n8308) );
  MUX2X1 U7858 ( .B(n8312), .A(n8313), .S(n8458), .Y(n8311) );
  MUX2X1 U7859 ( .B(n8315), .A(n8316), .S(n8458), .Y(n8314) );
  MUX2X1 U7860 ( .B(n8318), .A(n8319), .S(n8391), .Y(n8317) );
  MUX2X1 U7861 ( .B(ram[64]), .A(ram[0]), .S(n8482), .Y(n4341) );
  MUX2X1 U7862 ( .B(ram[192]), .A(ram[128]), .S(n8482), .Y(n4340) );
  MUX2X1 U7863 ( .B(ram[320]), .A(ram[256]), .S(n8482), .Y(n4344) );
  MUX2X1 U7864 ( .B(ram[448]), .A(ram[384]), .S(n8482), .Y(n4343) );
  MUX2X1 U7865 ( .B(n4342), .A(n4339), .S(n8396), .Y(n4353) );
  MUX2X1 U7866 ( .B(ram[576]), .A(ram[512]), .S(n8483), .Y(n4347) );
  MUX2X1 U7867 ( .B(ram[704]), .A(ram[640]), .S(n8483), .Y(n4346) );
  MUX2X1 U7868 ( .B(ram[832]), .A(ram[768]), .S(n8483), .Y(n4350) );
  MUX2X1 U7869 ( .B(ram[960]), .A(ram[896]), .S(n8483), .Y(n4349) );
  MUX2X1 U7870 ( .B(n4348), .A(n4345), .S(n8397), .Y(n4352) );
  MUX2X1 U7871 ( .B(ram[1088]), .A(ram[1024]), .S(n8483), .Y(n4356) );
  MUX2X1 U7872 ( .B(ram[1216]), .A(ram[1152]), .S(n8483), .Y(n4355) );
  MUX2X1 U7873 ( .B(ram[1344]), .A(ram[1280]), .S(n8483), .Y(n4359) );
  MUX2X1 U7874 ( .B(ram[1472]), .A(ram[1408]), .S(n8483), .Y(n4358) );
  MUX2X1 U7875 ( .B(n4357), .A(n4354), .S(n8400), .Y(n4368) );
  MUX2X1 U7876 ( .B(ram[1600]), .A(ram[1536]), .S(n8483), .Y(n4362) );
  MUX2X1 U7877 ( .B(ram[1728]), .A(ram[1664]), .S(n8483), .Y(n4361) );
  MUX2X1 U7878 ( .B(ram[1856]), .A(ram[1792]), .S(n8483), .Y(n4365) );
  MUX2X1 U7879 ( .B(ram[1984]), .A(ram[1920]), .S(n8483), .Y(n4364) );
  MUX2X1 U7880 ( .B(n4363), .A(n4360), .S(n8400), .Y(n4367) );
  MUX2X1 U7881 ( .B(n4366), .A(n4351), .S(n8387), .Y(n8320) );
  MUX2X1 U7882 ( .B(ram[65]), .A(ram[1]), .S(n8484), .Y(n4371) );
  MUX2X1 U7883 ( .B(ram[193]), .A(ram[129]), .S(n8484), .Y(n4370) );
  MUX2X1 U7884 ( .B(ram[321]), .A(ram[257]), .S(n8484), .Y(n4374) );
  MUX2X1 U7885 ( .B(ram[449]), .A(ram[385]), .S(n8484), .Y(n4373) );
  MUX2X1 U7886 ( .B(n4372), .A(n4369), .S(n8396), .Y(n4383) );
  MUX2X1 U7887 ( .B(ram[577]), .A(ram[513]), .S(n8484), .Y(n4377) );
  MUX2X1 U7888 ( .B(ram[705]), .A(ram[641]), .S(n8484), .Y(n4376) );
  MUX2X1 U7889 ( .B(ram[833]), .A(ram[769]), .S(n8484), .Y(n4380) );
  MUX2X1 U7890 ( .B(ram[961]), .A(ram[897]), .S(n8484), .Y(n4379) );
  MUX2X1 U7891 ( .B(n4378), .A(n4375), .S(n8396), .Y(n4382) );
  MUX2X1 U7892 ( .B(ram[1089]), .A(ram[1025]), .S(n8484), .Y(n4386) );
  MUX2X1 U7893 ( .B(ram[1217]), .A(ram[1153]), .S(n8484), .Y(n4385) );
  MUX2X1 U7894 ( .B(ram[1345]), .A(ram[1281]), .S(n8484), .Y(n4389) );
  MUX2X1 U7895 ( .B(ram[1473]), .A(ram[1409]), .S(n8484), .Y(n4388) );
  MUX2X1 U7896 ( .B(n4387), .A(n4384), .S(n8396), .Y(n4398) );
  MUX2X1 U7897 ( .B(ram[1601]), .A(ram[1537]), .S(n8485), .Y(n4392) );
  MUX2X1 U7898 ( .B(ram[1729]), .A(ram[1665]), .S(n8485), .Y(n4391) );
  MUX2X1 U7899 ( .B(ram[1857]), .A(ram[1793]), .S(n8485), .Y(n4395) );
  MUX2X1 U7900 ( .B(ram[1985]), .A(ram[1921]), .S(n8485), .Y(n4394) );
  MUX2X1 U7901 ( .B(n4393), .A(n4390), .S(n8396), .Y(n4397) );
  MUX2X1 U7902 ( .B(n4396), .A(n4381), .S(read1_addr[0]), .Y(n8321) );
  MUX2X1 U7903 ( .B(ram[66]), .A(ram[2]), .S(n8485), .Y(n4401) );
  MUX2X1 U7904 ( .B(ram[194]), .A(ram[130]), .S(n8485), .Y(n4400) );
  MUX2X1 U7905 ( .B(ram[322]), .A(ram[258]), .S(n8485), .Y(n4404) );
  MUX2X1 U7906 ( .B(ram[450]), .A(ram[386]), .S(n8485), .Y(n4403) );
  MUX2X1 U7907 ( .B(n4402), .A(n4399), .S(n8396), .Y(n4413) );
  MUX2X1 U7908 ( .B(ram[578]), .A(ram[514]), .S(n8485), .Y(n4407) );
  MUX2X1 U7909 ( .B(ram[706]), .A(ram[642]), .S(n8485), .Y(n4406) );
  MUX2X1 U7910 ( .B(ram[834]), .A(ram[770]), .S(n8485), .Y(n4410) );
  MUX2X1 U7911 ( .B(ram[962]), .A(ram[898]), .S(n8485), .Y(n4409) );
  MUX2X1 U7912 ( .B(n4408), .A(n4405), .S(n8396), .Y(n4412) );
  MUX2X1 U7913 ( .B(ram[1090]), .A(ram[1026]), .S(n8486), .Y(n4416) );
  MUX2X1 U7914 ( .B(ram[1218]), .A(ram[1154]), .S(n8486), .Y(n4415) );
  MUX2X1 U7915 ( .B(ram[1346]), .A(ram[1282]), .S(n8486), .Y(n4419) );
  MUX2X1 U7916 ( .B(ram[1474]), .A(ram[1410]), .S(n8486), .Y(n4418) );
  MUX2X1 U7917 ( .B(n4417), .A(n4414), .S(n8396), .Y(n4428) );
  MUX2X1 U7918 ( .B(ram[1602]), .A(ram[1538]), .S(n8486), .Y(n4422) );
  MUX2X1 U7919 ( .B(ram[1730]), .A(ram[1666]), .S(n8486), .Y(n4421) );
  MUX2X1 U7920 ( .B(ram[1858]), .A(ram[1794]), .S(n8486), .Y(n4425) );
  MUX2X1 U7921 ( .B(ram[1986]), .A(ram[1922]), .S(n8486), .Y(n4424) );
  MUX2X1 U7922 ( .B(n4423), .A(n4420), .S(n8396), .Y(n4427) );
  MUX2X1 U7923 ( .B(n4426), .A(n4411), .S(n8386), .Y(n8322) );
  MUX2X1 U7924 ( .B(ram[67]), .A(ram[3]), .S(n8486), .Y(n4431) );
  MUX2X1 U7925 ( .B(ram[195]), .A(ram[131]), .S(n8486), .Y(n4430) );
  MUX2X1 U7926 ( .B(ram[323]), .A(ram[259]), .S(n8486), .Y(n4434) );
  MUX2X1 U7927 ( .B(ram[451]), .A(ram[387]), .S(n8486), .Y(n4433) );
  MUX2X1 U7928 ( .B(n4432), .A(n4429), .S(n8396), .Y(n4443) );
  MUX2X1 U7929 ( .B(ram[579]), .A(ram[515]), .S(n8487), .Y(n4437) );
  MUX2X1 U7930 ( .B(ram[707]), .A(ram[643]), .S(n8487), .Y(n4436) );
  MUX2X1 U7931 ( .B(ram[835]), .A(ram[771]), .S(n8487), .Y(n4440) );
  MUX2X1 U7932 ( .B(ram[963]), .A(ram[899]), .S(n8487), .Y(n4439) );
  MUX2X1 U7933 ( .B(n4438), .A(n4435), .S(n8396), .Y(n4442) );
  MUX2X1 U7934 ( .B(ram[1091]), .A(ram[1027]), .S(n8487), .Y(n4446) );
  MUX2X1 U7935 ( .B(ram[1219]), .A(ram[1155]), .S(n8487), .Y(n4445) );
  MUX2X1 U7936 ( .B(ram[1347]), .A(ram[1283]), .S(n8487), .Y(n4449) );
  MUX2X1 U7937 ( .B(ram[1475]), .A(ram[1411]), .S(n8487), .Y(n4448) );
  MUX2X1 U7938 ( .B(n4447), .A(n4444), .S(n8396), .Y(n4458) );
  MUX2X1 U7939 ( .B(ram[1603]), .A(ram[1539]), .S(n8487), .Y(n4452) );
  MUX2X1 U7940 ( .B(ram[1731]), .A(ram[1667]), .S(n8487), .Y(n4451) );
  MUX2X1 U7941 ( .B(ram[1859]), .A(ram[1795]), .S(n8487), .Y(n4455) );
  MUX2X1 U7942 ( .B(ram[1987]), .A(ram[1923]), .S(n8487), .Y(n4454) );
  MUX2X1 U7943 ( .B(n4453), .A(n4450), .S(n8396), .Y(n4457) );
  MUX2X1 U7944 ( .B(n4456), .A(n4441), .S(n8386), .Y(n8323) );
  MUX2X1 U7945 ( .B(ram[68]), .A(ram[4]), .S(n8488), .Y(n4461) );
  MUX2X1 U7946 ( .B(ram[196]), .A(ram[132]), .S(n8488), .Y(n4460) );
  MUX2X1 U7947 ( .B(ram[324]), .A(ram[260]), .S(n8488), .Y(n4464) );
  MUX2X1 U7948 ( .B(ram[452]), .A(ram[388]), .S(n8488), .Y(n4463) );
  MUX2X1 U7949 ( .B(n4462), .A(n4459), .S(n8399), .Y(n4473) );
  MUX2X1 U7950 ( .B(ram[580]), .A(ram[516]), .S(n8488), .Y(n4467) );
  MUX2X1 U7951 ( .B(ram[708]), .A(ram[644]), .S(n8488), .Y(n4466) );
  MUX2X1 U7952 ( .B(ram[836]), .A(ram[772]), .S(n8488), .Y(n4470) );
  MUX2X1 U7953 ( .B(ram[964]), .A(ram[900]), .S(n8488), .Y(n4469) );
  MUX2X1 U7954 ( .B(n4468), .A(n4465), .S(n8399), .Y(n4472) );
  MUX2X1 U7955 ( .B(ram[1092]), .A(ram[1028]), .S(n8488), .Y(n4476) );
  MUX2X1 U7956 ( .B(ram[1220]), .A(ram[1156]), .S(n8488), .Y(n4475) );
  MUX2X1 U7957 ( .B(ram[1348]), .A(ram[1284]), .S(n8488), .Y(n4479) );
  MUX2X1 U7958 ( .B(ram[1476]), .A(ram[1412]), .S(n8488), .Y(n4478) );
  MUX2X1 U7959 ( .B(n4477), .A(n4474), .S(n8396), .Y(n4488) );
  MUX2X1 U7960 ( .B(ram[1604]), .A(ram[1540]), .S(n8489), .Y(n4482) );
  MUX2X1 U7961 ( .B(ram[1732]), .A(ram[1668]), .S(n8489), .Y(n4481) );
  MUX2X1 U7962 ( .B(ram[1860]), .A(ram[1796]), .S(n8489), .Y(n4485) );
  MUX2X1 U7963 ( .B(ram[1988]), .A(ram[1924]), .S(n8489), .Y(n4484) );
  MUX2X1 U7964 ( .B(n4483), .A(n4480), .S(n8403), .Y(n4487) );
  MUX2X1 U7965 ( .B(n4486), .A(n4471), .S(read1_addr[0]), .Y(n8324) );
  MUX2X1 U7966 ( .B(ram[69]), .A(ram[5]), .S(n8489), .Y(n4491) );
  MUX2X1 U7967 ( .B(ram[197]), .A(ram[133]), .S(n8489), .Y(n4490) );
  MUX2X1 U7968 ( .B(ram[325]), .A(ram[261]), .S(n8489), .Y(n4494) );
  MUX2X1 U7969 ( .B(ram[453]), .A(ram[389]), .S(n8489), .Y(n4493) );
  MUX2X1 U7970 ( .B(n4492), .A(n4489), .S(n8401), .Y(n4503) );
  MUX2X1 U7971 ( .B(ram[581]), .A(ram[517]), .S(n8489), .Y(n4497) );
  MUX2X1 U7972 ( .B(ram[709]), .A(ram[645]), .S(n8489), .Y(n4496) );
  MUX2X1 U7973 ( .B(ram[837]), .A(ram[773]), .S(n8489), .Y(n4500) );
  MUX2X1 U7974 ( .B(ram[965]), .A(ram[901]), .S(n8489), .Y(n4499) );
  MUX2X1 U7975 ( .B(n4498), .A(n4495), .S(n8404), .Y(n4502) );
  MUX2X1 U7976 ( .B(ram[1093]), .A(ram[1029]), .S(n8490), .Y(n4506) );
  MUX2X1 U7977 ( .B(ram[1221]), .A(ram[1157]), .S(n8490), .Y(n4505) );
  MUX2X1 U7978 ( .B(ram[1349]), .A(ram[1285]), .S(n8490), .Y(n4510) );
  MUX2X1 U7979 ( .B(ram[1477]), .A(ram[1413]), .S(n8490), .Y(n4509) );
  MUX2X1 U7980 ( .B(n4507), .A(n4504), .S(n8406), .Y(n4519) );
  MUX2X1 U7981 ( .B(ram[1605]), .A(ram[1541]), .S(n8490), .Y(n4513) );
  MUX2X1 U7982 ( .B(ram[1733]), .A(ram[1669]), .S(n8490), .Y(n4512) );
  MUX2X1 U7983 ( .B(ram[1861]), .A(ram[1797]), .S(n8490), .Y(n4516) );
  MUX2X1 U7984 ( .B(ram[1989]), .A(ram[1925]), .S(n8490), .Y(n4515) );
  MUX2X1 U7985 ( .B(n4514), .A(n4511), .S(n8402), .Y(n4518) );
  MUX2X1 U7986 ( .B(n4517), .A(n4501), .S(n8385), .Y(n8325) );
  MUX2X1 U7987 ( .B(ram[70]), .A(ram[6]), .S(n8490), .Y(n4522) );
  MUX2X1 U7988 ( .B(ram[198]), .A(ram[134]), .S(n8490), .Y(n4521) );
  MUX2X1 U7989 ( .B(ram[326]), .A(ram[262]), .S(n8490), .Y(n4525) );
  MUX2X1 U7990 ( .B(ram[454]), .A(ram[390]), .S(n8490), .Y(n4524) );
  MUX2X1 U7991 ( .B(n4523), .A(n4520), .S(n8410), .Y(n4534) );
  MUX2X1 U7992 ( .B(ram[582]), .A(ram[518]), .S(n8491), .Y(n4528) );
  MUX2X1 U7993 ( .B(ram[710]), .A(ram[646]), .S(n8491), .Y(n4527) );
  MUX2X1 U7994 ( .B(ram[838]), .A(ram[774]), .S(n8491), .Y(n4531) );
  MUX2X1 U7995 ( .B(ram[966]), .A(ram[902]), .S(n8491), .Y(n4530) );
  MUX2X1 U7996 ( .B(n4529), .A(n4526), .S(n8409), .Y(n4533) );
  MUX2X1 U7997 ( .B(ram[1094]), .A(ram[1030]), .S(n8491), .Y(n4537) );
  MUX2X1 U7998 ( .B(ram[1222]), .A(ram[1158]), .S(n8491), .Y(n4536) );
  MUX2X1 U7999 ( .B(ram[1350]), .A(ram[1286]), .S(n8491), .Y(n4540) );
  MUX2X1 U8000 ( .B(ram[1478]), .A(ram[1414]), .S(n8491), .Y(n4539) );
  MUX2X1 U8001 ( .B(n4538), .A(n4535), .S(n8407), .Y(n4549) );
  MUX2X1 U8002 ( .B(ram[1606]), .A(ram[1542]), .S(n8491), .Y(n4543) );
  MUX2X1 U8003 ( .B(ram[1734]), .A(ram[1670]), .S(n8491), .Y(n4542) );
  MUX2X1 U8004 ( .B(ram[1862]), .A(ram[1798]), .S(n8491), .Y(n4546) );
  MUX2X1 U8005 ( .B(ram[1990]), .A(ram[1926]), .S(n8491), .Y(n4545) );
  MUX2X1 U8006 ( .B(n4544), .A(n4541), .S(n8398), .Y(n4548) );
  MUX2X1 U8007 ( .B(n4547), .A(n4532), .S(n8386), .Y(n8326) );
  MUX2X1 U8008 ( .B(ram[71]), .A(ram[7]), .S(n8492), .Y(n4552) );
  MUX2X1 U8009 ( .B(ram[199]), .A(ram[135]), .S(n8492), .Y(n4551) );
  MUX2X1 U8010 ( .B(ram[327]), .A(ram[263]), .S(n8492), .Y(n4555) );
  MUX2X1 U8011 ( .B(ram[455]), .A(ram[391]), .S(n8492), .Y(n4554) );
  MUX2X1 U8012 ( .B(n4553), .A(n4550), .S(n8397), .Y(n4564) );
  MUX2X1 U8013 ( .B(ram[583]), .A(ram[519]), .S(n8492), .Y(n4558) );
  MUX2X1 U8014 ( .B(ram[711]), .A(ram[647]), .S(n8492), .Y(n4557) );
  MUX2X1 U8015 ( .B(ram[839]), .A(ram[775]), .S(n8492), .Y(n4561) );
  MUX2X1 U8016 ( .B(ram[967]), .A(ram[903]), .S(n8492), .Y(n4560) );
  MUX2X1 U8017 ( .B(n4559), .A(n4556), .S(n8397), .Y(n4563) );
  MUX2X1 U8018 ( .B(ram[1095]), .A(ram[1031]), .S(n8492), .Y(n4567) );
  MUX2X1 U8019 ( .B(ram[1223]), .A(ram[1159]), .S(n8492), .Y(n4566) );
  MUX2X1 U8020 ( .B(ram[1351]), .A(ram[1287]), .S(n8492), .Y(n4570) );
  MUX2X1 U8021 ( .B(ram[1479]), .A(ram[1415]), .S(n8492), .Y(n4569) );
  MUX2X1 U8022 ( .B(n4568), .A(n4565), .S(n8397), .Y(n4584) );
  MUX2X1 U8023 ( .B(ram[1607]), .A(ram[1543]), .S(n8493), .Y(n4573) );
  MUX2X1 U8024 ( .B(ram[1735]), .A(ram[1671]), .S(n8493), .Y(n4572) );
  MUX2X1 U8025 ( .B(ram[1863]), .A(ram[1799]), .S(n8493), .Y(n4581) );
  MUX2X1 U8026 ( .B(ram[1991]), .A(ram[1927]), .S(n8493), .Y(n4575) );
  MUX2X1 U8027 ( .B(n4574), .A(n4571), .S(n8397), .Y(n4583) );
  MUX2X1 U8028 ( .B(n4582), .A(n4562), .S(read1_addr[0]), .Y(n8327) );
  MUX2X1 U8029 ( .B(ram[72]), .A(ram[8]), .S(n8493), .Y(n4587) );
  MUX2X1 U8030 ( .B(ram[200]), .A(ram[136]), .S(n8493), .Y(n4586) );
  MUX2X1 U8031 ( .B(ram[328]), .A(ram[264]), .S(n8493), .Y(n4590) );
  MUX2X1 U8032 ( .B(ram[456]), .A(ram[392]), .S(n8493), .Y(n4589) );
  MUX2X1 U8033 ( .B(n4588), .A(n4585), .S(n8397), .Y(n4599) );
  MUX2X1 U8034 ( .B(ram[584]), .A(ram[520]), .S(n8493), .Y(n4593) );
  MUX2X1 U8035 ( .B(ram[712]), .A(ram[648]), .S(n8493), .Y(n4592) );
  MUX2X1 U8036 ( .B(ram[840]), .A(ram[776]), .S(n8493), .Y(n4596) );
  MUX2X1 U8037 ( .B(ram[968]), .A(ram[904]), .S(n8493), .Y(n4595) );
  MUX2X1 U8038 ( .B(n4594), .A(n4591), .S(n8397), .Y(n4598) );
  MUX2X1 U8039 ( .B(ram[1096]), .A(ram[1032]), .S(n8494), .Y(n4602) );
  MUX2X1 U8040 ( .B(ram[1224]), .A(ram[1160]), .S(n8494), .Y(n4601) );
  MUX2X1 U8041 ( .B(ram[1352]), .A(ram[1288]), .S(n8494), .Y(n4605) );
  MUX2X1 U8042 ( .B(ram[1480]), .A(ram[1416]), .S(n8494), .Y(n4604) );
  MUX2X1 U8043 ( .B(n4603), .A(n4600), .S(n8397), .Y(n4614) );
  MUX2X1 U8044 ( .B(ram[1608]), .A(ram[1544]), .S(n8494), .Y(n4608) );
  MUX2X1 U8045 ( .B(ram[1736]), .A(ram[1672]), .S(n8494), .Y(n4607) );
  MUX2X1 U8046 ( .B(ram[1864]), .A(ram[1800]), .S(n8494), .Y(n4611) );
  MUX2X1 U8047 ( .B(ram[1992]), .A(ram[1928]), .S(n8494), .Y(n4610) );
  MUX2X1 U8048 ( .B(n4609), .A(n4606), .S(n8397), .Y(n4613) );
  MUX2X1 U8049 ( .B(n4612), .A(n4597), .S(read1_addr[0]), .Y(n8328) );
  MUX2X1 U8050 ( .B(ram[73]), .A(ram[9]), .S(n8494), .Y(n4617) );
  MUX2X1 U8051 ( .B(ram[201]), .A(ram[137]), .S(n8494), .Y(n4616) );
  MUX2X1 U8052 ( .B(ram[329]), .A(ram[265]), .S(n8494), .Y(n4620) );
  MUX2X1 U8053 ( .B(ram[457]), .A(ram[393]), .S(n8494), .Y(n4619) );
  MUX2X1 U8054 ( .B(n4618), .A(n4615), .S(n8397), .Y(n4629) );
  MUX2X1 U8055 ( .B(ram[585]), .A(ram[521]), .S(n8495), .Y(n4623) );
  MUX2X1 U8056 ( .B(ram[713]), .A(ram[649]), .S(n8495), .Y(n4622) );
  MUX2X1 U8057 ( .B(ram[841]), .A(ram[777]), .S(n8495), .Y(n4626) );
  MUX2X1 U8058 ( .B(ram[969]), .A(ram[905]), .S(n8495), .Y(n4625) );
  MUX2X1 U8059 ( .B(n4624), .A(n4621), .S(n8397), .Y(n4628) );
  MUX2X1 U8060 ( .B(ram[1097]), .A(ram[1033]), .S(n8495), .Y(n4632) );
  MUX2X1 U8061 ( .B(ram[1225]), .A(ram[1161]), .S(n8495), .Y(n4631) );
  MUX2X1 U8062 ( .B(ram[1353]), .A(ram[1289]), .S(n8495), .Y(n4635) );
  MUX2X1 U8063 ( .B(ram[1481]), .A(ram[1417]), .S(n8495), .Y(n4634) );
  MUX2X1 U8064 ( .B(n4633), .A(n4630), .S(n8397), .Y(n4644) );
  MUX2X1 U8065 ( .B(ram[1609]), .A(ram[1545]), .S(n8495), .Y(n4638) );
  MUX2X1 U8066 ( .B(ram[1737]), .A(ram[1673]), .S(n8495), .Y(n4637) );
  MUX2X1 U8067 ( .B(ram[1865]), .A(ram[1801]), .S(n8495), .Y(n4641) );
  MUX2X1 U8068 ( .B(ram[1993]), .A(ram[1929]), .S(n8495), .Y(n4640) );
  MUX2X1 U8069 ( .B(n4639), .A(n4636), .S(n8397), .Y(n4643) );
  MUX2X1 U8070 ( .B(n4642), .A(n4627), .S(read1_addr[0]), .Y(n8329) );
  MUX2X1 U8071 ( .B(ram[74]), .A(ram[10]), .S(n8496), .Y(n4647) );
  MUX2X1 U8072 ( .B(ram[202]), .A(ram[138]), .S(n8496), .Y(n4646) );
  MUX2X1 U8073 ( .B(ram[330]), .A(ram[266]), .S(n8496), .Y(n4650) );
  MUX2X1 U8074 ( .B(ram[458]), .A(ram[394]), .S(n8496), .Y(n4649) );
  MUX2X1 U8075 ( .B(n4648), .A(n4645), .S(n8398), .Y(n4659) );
  MUX2X1 U8076 ( .B(ram[586]), .A(ram[522]), .S(n8496), .Y(n4653) );
  MUX2X1 U8077 ( .B(ram[714]), .A(ram[650]), .S(n8496), .Y(n4652) );
  MUX2X1 U8078 ( .B(ram[842]), .A(ram[778]), .S(n8496), .Y(n4656) );
  MUX2X1 U8079 ( .B(ram[970]), .A(ram[906]), .S(n8496), .Y(n4655) );
  MUX2X1 U8080 ( .B(n4654), .A(n4651), .S(n8398), .Y(n4658) );
  MUX2X1 U8081 ( .B(ram[1098]), .A(ram[1034]), .S(n8496), .Y(n6717) );
  MUX2X1 U8082 ( .B(ram[1226]), .A(ram[1162]), .S(n8496), .Y(n4661) );
  MUX2X1 U8083 ( .B(ram[1354]), .A(ram[1290]), .S(n8496), .Y(n6720) );
  MUX2X1 U8084 ( .B(ram[1482]), .A(ram[1418]), .S(n8496), .Y(n6719) );
  MUX2X1 U8085 ( .B(n6718), .A(n4660), .S(n8398), .Y(n6729) );
  MUX2X1 U8086 ( .B(ram[1610]), .A(ram[1546]), .S(n8497), .Y(n6723) );
  MUX2X1 U8087 ( .B(ram[1738]), .A(ram[1674]), .S(n8497), .Y(n6722) );
  MUX2X1 U8088 ( .B(ram[1866]), .A(ram[1802]), .S(n8497), .Y(n6726) );
  MUX2X1 U8089 ( .B(ram[1994]), .A(ram[1930]), .S(n8497), .Y(n6725) );
  MUX2X1 U8090 ( .B(n6724), .A(n6721), .S(n8398), .Y(n6728) );
  MUX2X1 U8091 ( .B(n6727), .A(n4657), .S(read1_addr[0]), .Y(n8330) );
  MUX2X1 U8092 ( .B(ram[75]), .A(ram[11]), .S(n8497), .Y(n6732) );
  MUX2X1 U8093 ( .B(ram[203]), .A(ram[139]), .S(n8497), .Y(n6731) );
  MUX2X1 U8094 ( .B(ram[331]), .A(ram[267]), .S(n8497), .Y(n6735) );
  MUX2X1 U8095 ( .B(ram[459]), .A(ram[395]), .S(n8497), .Y(n6734) );
  MUX2X1 U8096 ( .B(n6733), .A(n6730), .S(n8398), .Y(n6744) );
  MUX2X1 U8097 ( .B(ram[587]), .A(ram[523]), .S(n8497), .Y(n6738) );
  MUX2X1 U8098 ( .B(ram[715]), .A(ram[651]), .S(n8497), .Y(n6737) );
  MUX2X1 U8099 ( .B(ram[843]), .A(ram[779]), .S(n8497), .Y(n6741) );
  MUX2X1 U8100 ( .B(ram[971]), .A(ram[907]), .S(n8497), .Y(n6740) );
  MUX2X1 U8101 ( .B(n6739), .A(n6736), .S(n8398), .Y(n6743) );
  MUX2X1 U8102 ( .B(ram[1099]), .A(ram[1035]), .S(n8498), .Y(n6747) );
  MUX2X1 U8103 ( .B(ram[1227]), .A(ram[1163]), .S(n8498), .Y(n6746) );
  MUX2X1 U8104 ( .B(ram[1355]), .A(ram[1291]), .S(n8498), .Y(n6750) );
  MUX2X1 U8105 ( .B(ram[1483]), .A(ram[1419]), .S(n8498), .Y(n6749) );
  MUX2X1 U8106 ( .B(n6748), .A(n6745), .S(n8398), .Y(n6759) );
  MUX2X1 U8107 ( .B(ram[1611]), .A(ram[1547]), .S(n8498), .Y(n6753) );
  MUX2X1 U8108 ( .B(ram[1739]), .A(ram[1675]), .S(n8498), .Y(n6752) );
  MUX2X1 U8109 ( .B(ram[1867]), .A(ram[1803]), .S(n8498), .Y(n6756) );
  MUX2X1 U8110 ( .B(ram[1995]), .A(ram[1931]), .S(n8498), .Y(n6755) );
  MUX2X1 U8111 ( .B(n6754), .A(n6751), .S(n8398), .Y(n6758) );
  MUX2X1 U8112 ( .B(n6757), .A(n6742), .S(read1_addr[0]), .Y(n8331) );
  MUX2X1 U8113 ( .B(ram[76]), .A(ram[12]), .S(n8498), .Y(n6762) );
  MUX2X1 U8114 ( .B(ram[204]), .A(ram[140]), .S(n8498), .Y(n6761) );
  MUX2X1 U8115 ( .B(ram[332]), .A(ram[268]), .S(n8498), .Y(n6765) );
  MUX2X1 U8116 ( .B(ram[460]), .A(ram[396]), .S(n8498), .Y(n6764) );
  MUX2X1 U8117 ( .B(n6763), .A(n6760), .S(n8398), .Y(n6774) );
  MUX2X1 U8118 ( .B(ram[588]), .A(ram[524]), .S(n8499), .Y(n6768) );
  MUX2X1 U8119 ( .B(ram[716]), .A(ram[652]), .S(n8499), .Y(n6767) );
  MUX2X1 U8120 ( .B(ram[844]), .A(ram[780]), .S(n8499), .Y(n6771) );
  MUX2X1 U8121 ( .B(ram[972]), .A(ram[908]), .S(n8499), .Y(n6770) );
  MUX2X1 U8122 ( .B(n6769), .A(n6766), .S(n8398), .Y(n6773) );
  MUX2X1 U8123 ( .B(ram[1100]), .A(ram[1036]), .S(n8499), .Y(n6777) );
  MUX2X1 U8124 ( .B(ram[1228]), .A(ram[1164]), .S(n8499), .Y(n6776) );
  MUX2X1 U8125 ( .B(ram[1356]), .A(ram[1292]), .S(n8499), .Y(n6780) );
  MUX2X1 U8126 ( .B(ram[1484]), .A(ram[1420]), .S(n8499), .Y(n6779) );
  MUX2X1 U8127 ( .B(n6778), .A(n6775), .S(n8398), .Y(n6789) );
  MUX2X1 U8128 ( .B(ram[1612]), .A(ram[1548]), .S(n8499), .Y(n6783) );
  MUX2X1 U8129 ( .B(ram[1740]), .A(ram[1676]), .S(n8499), .Y(n6782) );
  MUX2X1 U8130 ( .B(ram[1868]), .A(ram[1804]), .S(n8499), .Y(n6786) );
  MUX2X1 U8131 ( .B(ram[1996]), .A(ram[1932]), .S(n8499), .Y(n6785) );
  MUX2X1 U8132 ( .B(n6784), .A(n6781), .S(n8398), .Y(n6788) );
  MUX2X1 U8133 ( .B(n6787), .A(n6772), .S(n8387), .Y(n8332) );
  MUX2X1 U8134 ( .B(ram[77]), .A(ram[13]), .S(n8500), .Y(n6792) );
  MUX2X1 U8135 ( .B(ram[205]), .A(ram[141]), .S(n8500), .Y(n6791) );
  MUX2X1 U8136 ( .B(ram[333]), .A(ram[269]), .S(n8500), .Y(n6795) );
  MUX2X1 U8137 ( .B(ram[461]), .A(ram[397]), .S(n8500), .Y(n6794) );
  MUX2X1 U8138 ( .B(n6793), .A(n6790), .S(n8399), .Y(n6804) );
  MUX2X1 U8139 ( .B(ram[589]), .A(ram[525]), .S(n8500), .Y(n6798) );
  MUX2X1 U8140 ( .B(ram[717]), .A(ram[653]), .S(n8500), .Y(n6797) );
  MUX2X1 U8141 ( .B(ram[845]), .A(ram[781]), .S(n8500), .Y(n6801) );
  MUX2X1 U8142 ( .B(ram[973]), .A(ram[909]), .S(n8500), .Y(n6800) );
  MUX2X1 U8143 ( .B(n6799), .A(n6796), .S(n8399), .Y(n6803) );
  MUX2X1 U8144 ( .B(ram[1101]), .A(ram[1037]), .S(n8500), .Y(n6807) );
  MUX2X1 U8145 ( .B(ram[1229]), .A(ram[1165]), .S(n8500), .Y(n6806) );
  MUX2X1 U8146 ( .B(ram[1357]), .A(ram[1293]), .S(n8500), .Y(n6810) );
  MUX2X1 U8147 ( .B(ram[1485]), .A(ram[1421]), .S(n8500), .Y(n6809) );
  MUX2X1 U8148 ( .B(n6808), .A(n6805), .S(n8399), .Y(n6819) );
  MUX2X1 U8149 ( .B(ram[1613]), .A(ram[1549]), .S(n8501), .Y(n6813) );
  MUX2X1 U8150 ( .B(ram[1741]), .A(ram[1677]), .S(n8501), .Y(n6812) );
  MUX2X1 U8151 ( .B(ram[1869]), .A(ram[1805]), .S(n8501), .Y(n6816) );
  MUX2X1 U8152 ( .B(ram[1997]), .A(ram[1933]), .S(n8501), .Y(n6815) );
  MUX2X1 U8153 ( .B(n6814), .A(n6811), .S(n8399), .Y(n6818) );
  MUX2X1 U8154 ( .B(n6817), .A(n6802), .S(n8387), .Y(n8333) );
  MUX2X1 U8155 ( .B(ram[78]), .A(ram[14]), .S(n8501), .Y(n6822) );
  MUX2X1 U8156 ( .B(ram[206]), .A(ram[142]), .S(n8501), .Y(n6821) );
  MUX2X1 U8157 ( .B(ram[334]), .A(ram[270]), .S(n8501), .Y(n6825) );
  MUX2X1 U8158 ( .B(ram[462]), .A(ram[398]), .S(n8501), .Y(n6824) );
  MUX2X1 U8159 ( .B(n6823), .A(n6820), .S(n8399), .Y(n6834) );
  MUX2X1 U8160 ( .B(ram[590]), .A(ram[526]), .S(n8501), .Y(n6828) );
  MUX2X1 U8161 ( .B(ram[718]), .A(ram[654]), .S(n8501), .Y(n6827) );
  MUX2X1 U8162 ( .B(ram[846]), .A(ram[782]), .S(n8501), .Y(n6831) );
  MUX2X1 U8163 ( .B(ram[974]), .A(ram[910]), .S(n8501), .Y(n6830) );
  MUX2X1 U8164 ( .B(n6829), .A(n6826), .S(n8399), .Y(n6833) );
  MUX2X1 U8165 ( .B(ram[1102]), .A(ram[1038]), .S(n8502), .Y(n6837) );
  MUX2X1 U8166 ( .B(ram[1230]), .A(ram[1166]), .S(n8502), .Y(n6836) );
  MUX2X1 U8167 ( .B(ram[1358]), .A(ram[1294]), .S(n8502), .Y(n6840) );
  MUX2X1 U8168 ( .B(ram[1486]), .A(ram[1422]), .S(n8502), .Y(n6839) );
  MUX2X1 U8169 ( .B(n6838), .A(n6835), .S(n8399), .Y(n6849) );
  MUX2X1 U8170 ( .B(ram[1614]), .A(ram[1550]), .S(n8502), .Y(n6843) );
  MUX2X1 U8171 ( .B(ram[1742]), .A(ram[1678]), .S(n8502), .Y(n6842) );
  MUX2X1 U8172 ( .B(ram[1870]), .A(ram[1806]), .S(n8502), .Y(n6846) );
  MUX2X1 U8173 ( .B(ram[1998]), .A(ram[1934]), .S(n8502), .Y(n6845) );
  MUX2X1 U8174 ( .B(n6844), .A(n6841), .S(n8399), .Y(n6848) );
  MUX2X1 U8175 ( .B(n6847), .A(n6832), .S(n8387), .Y(n8334) );
  MUX2X1 U8176 ( .B(ram[79]), .A(ram[15]), .S(n8502), .Y(n6852) );
  MUX2X1 U8177 ( .B(ram[207]), .A(ram[143]), .S(n8502), .Y(n6851) );
  MUX2X1 U8178 ( .B(ram[335]), .A(ram[271]), .S(n8502), .Y(n6855) );
  MUX2X1 U8179 ( .B(ram[463]), .A(ram[399]), .S(n8502), .Y(n6854) );
  MUX2X1 U8180 ( .B(n6853), .A(n6850), .S(n8399), .Y(n6864) );
  MUX2X1 U8181 ( .B(ram[591]), .A(ram[527]), .S(n8503), .Y(n6858) );
  MUX2X1 U8182 ( .B(ram[719]), .A(ram[655]), .S(n8503), .Y(n6857) );
  MUX2X1 U8183 ( .B(ram[847]), .A(ram[783]), .S(n8503), .Y(n6861) );
  MUX2X1 U8184 ( .B(ram[975]), .A(ram[911]), .S(n8503), .Y(n6860) );
  MUX2X1 U8185 ( .B(n6859), .A(n6856), .S(n8399), .Y(n6863) );
  MUX2X1 U8186 ( .B(ram[1103]), .A(ram[1039]), .S(n8503), .Y(n6867) );
  MUX2X1 U8187 ( .B(ram[1231]), .A(ram[1167]), .S(n8503), .Y(n6866) );
  MUX2X1 U8188 ( .B(ram[1359]), .A(ram[1295]), .S(n8503), .Y(n6870) );
  MUX2X1 U8189 ( .B(ram[1487]), .A(ram[1423]), .S(n8503), .Y(n6869) );
  MUX2X1 U8190 ( .B(n6868), .A(n6865), .S(n8399), .Y(n6879) );
  MUX2X1 U8191 ( .B(ram[1615]), .A(ram[1551]), .S(n8503), .Y(n6873) );
  MUX2X1 U8192 ( .B(ram[1743]), .A(ram[1679]), .S(n8503), .Y(n6872) );
  MUX2X1 U8193 ( .B(ram[1871]), .A(ram[1807]), .S(n8503), .Y(n6876) );
  MUX2X1 U8194 ( .B(ram[1999]), .A(ram[1935]), .S(n8503), .Y(n6875) );
  MUX2X1 U8195 ( .B(n6874), .A(n6871), .S(n8399), .Y(n6878) );
  MUX2X1 U8196 ( .B(n6877), .A(n6862), .S(n8387), .Y(n8335) );
  MUX2X1 U8197 ( .B(ram[80]), .A(ram[16]), .S(n8504), .Y(n6882) );
  MUX2X1 U8198 ( .B(ram[208]), .A(ram[144]), .S(n8504), .Y(n6881) );
  MUX2X1 U8199 ( .B(ram[336]), .A(ram[272]), .S(n8504), .Y(n6885) );
  MUX2X1 U8200 ( .B(ram[464]), .A(ram[400]), .S(n8504), .Y(n6884) );
  MUX2X1 U8201 ( .B(n6883), .A(n6880), .S(n8400), .Y(n6894) );
  MUX2X1 U8202 ( .B(ram[592]), .A(ram[528]), .S(n8504), .Y(n6888) );
  MUX2X1 U8203 ( .B(ram[720]), .A(ram[656]), .S(n8504), .Y(n6887) );
  MUX2X1 U8204 ( .B(ram[848]), .A(ram[784]), .S(n8504), .Y(n6891) );
  MUX2X1 U8205 ( .B(ram[976]), .A(ram[912]), .S(n8504), .Y(n6890) );
  MUX2X1 U8206 ( .B(n6889), .A(n6886), .S(n8400), .Y(n6893) );
  MUX2X1 U8207 ( .B(ram[1104]), .A(ram[1040]), .S(n8504), .Y(n6897) );
  MUX2X1 U8208 ( .B(ram[1232]), .A(ram[1168]), .S(n8504), .Y(n6896) );
  MUX2X1 U8209 ( .B(ram[1360]), .A(ram[1296]), .S(n8504), .Y(n6900) );
  MUX2X1 U8210 ( .B(ram[1488]), .A(ram[1424]), .S(n8504), .Y(n6899) );
  MUX2X1 U8211 ( .B(n6898), .A(n6895), .S(n8400), .Y(n6909) );
  MUX2X1 U8212 ( .B(ram[1616]), .A(ram[1552]), .S(n8505), .Y(n6903) );
  MUX2X1 U8213 ( .B(ram[1744]), .A(ram[1680]), .S(n8505), .Y(n6902) );
  MUX2X1 U8214 ( .B(ram[1872]), .A(ram[1808]), .S(n8505), .Y(n6906) );
  MUX2X1 U8215 ( .B(ram[2000]), .A(ram[1936]), .S(n8505), .Y(n6905) );
  MUX2X1 U8216 ( .B(n6904), .A(n6901), .S(n8400), .Y(n6908) );
  MUX2X1 U8217 ( .B(n6907), .A(n6892), .S(n8387), .Y(n8336) );
  MUX2X1 U8218 ( .B(ram[81]), .A(ram[17]), .S(n8505), .Y(n6912) );
  MUX2X1 U8219 ( .B(ram[209]), .A(ram[145]), .S(n8505), .Y(n6911) );
  MUX2X1 U8220 ( .B(ram[337]), .A(ram[273]), .S(n8505), .Y(n6915) );
  MUX2X1 U8221 ( .B(ram[465]), .A(ram[401]), .S(n8505), .Y(n6914) );
  MUX2X1 U8222 ( .B(n6913), .A(n6910), .S(n8400), .Y(n6924) );
  MUX2X1 U8223 ( .B(ram[593]), .A(ram[529]), .S(n8505), .Y(n6918) );
  MUX2X1 U8224 ( .B(ram[721]), .A(ram[657]), .S(n8505), .Y(n6917) );
  MUX2X1 U8225 ( .B(ram[849]), .A(ram[785]), .S(n8505), .Y(n6921) );
  MUX2X1 U8226 ( .B(ram[977]), .A(ram[913]), .S(n8505), .Y(n6920) );
  MUX2X1 U8227 ( .B(n6919), .A(n6916), .S(n8400), .Y(n6923) );
  MUX2X1 U8228 ( .B(ram[1105]), .A(ram[1041]), .S(n8506), .Y(n6927) );
  MUX2X1 U8229 ( .B(ram[1233]), .A(ram[1169]), .S(n8506), .Y(n6926) );
  MUX2X1 U8230 ( .B(ram[1361]), .A(ram[1297]), .S(n8506), .Y(n6930) );
  MUX2X1 U8231 ( .B(ram[1489]), .A(ram[1425]), .S(n8506), .Y(n6929) );
  MUX2X1 U8232 ( .B(n6928), .A(n6925), .S(n8400), .Y(n6939) );
  MUX2X1 U8233 ( .B(ram[1617]), .A(ram[1553]), .S(n8506), .Y(n6933) );
  MUX2X1 U8234 ( .B(ram[1745]), .A(ram[1681]), .S(n8506), .Y(n6932) );
  MUX2X1 U8235 ( .B(ram[1873]), .A(ram[1809]), .S(n8506), .Y(n6936) );
  MUX2X1 U8236 ( .B(ram[2001]), .A(ram[1937]), .S(n8506), .Y(n6935) );
  MUX2X1 U8237 ( .B(n6934), .A(n6931), .S(n8400), .Y(n6938) );
  MUX2X1 U8238 ( .B(n6937), .A(n6922), .S(n8387), .Y(n8337) );
  MUX2X1 U8239 ( .B(ram[82]), .A(ram[18]), .S(n8506), .Y(n6942) );
  MUX2X1 U8240 ( .B(ram[210]), .A(ram[146]), .S(n8506), .Y(n6941) );
  MUX2X1 U8241 ( .B(ram[338]), .A(ram[274]), .S(n8506), .Y(n6945) );
  MUX2X1 U8242 ( .B(ram[466]), .A(ram[402]), .S(n8506), .Y(n6944) );
  MUX2X1 U8243 ( .B(n6943), .A(n6940), .S(n8400), .Y(n6954) );
  MUX2X1 U8244 ( .B(ram[594]), .A(ram[530]), .S(n8507), .Y(n6948) );
  MUX2X1 U8245 ( .B(ram[722]), .A(ram[658]), .S(n8507), .Y(n6947) );
  MUX2X1 U8246 ( .B(ram[850]), .A(ram[786]), .S(n8507), .Y(n6951) );
  MUX2X1 U8247 ( .B(ram[978]), .A(ram[914]), .S(n8507), .Y(n6950) );
  MUX2X1 U8248 ( .B(n6949), .A(n6946), .S(n8400), .Y(n6953) );
  MUX2X1 U8249 ( .B(ram[1106]), .A(ram[1042]), .S(n8507), .Y(n6957) );
  MUX2X1 U8250 ( .B(ram[1234]), .A(ram[1170]), .S(n8507), .Y(n6956) );
  MUX2X1 U8251 ( .B(ram[1362]), .A(ram[1298]), .S(n8507), .Y(n6960) );
  MUX2X1 U8252 ( .B(ram[1490]), .A(ram[1426]), .S(n8507), .Y(n6959) );
  MUX2X1 U8253 ( .B(n6958), .A(n6955), .S(n8400), .Y(n6969) );
  MUX2X1 U8254 ( .B(ram[1618]), .A(ram[1554]), .S(n8507), .Y(n6963) );
  MUX2X1 U8255 ( .B(ram[1746]), .A(ram[1682]), .S(n8507), .Y(n6962) );
  MUX2X1 U8256 ( .B(ram[1874]), .A(ram[1810]), .S(n8507), .Y(n6966) );
  MUX2X1 U8257 ( .B(ram[2002]), .A(ram[1938]), .S(n8507), .Y(n6965) );
  MUX2X1 U8258 ( .B(n6964), .A(n6961), .S(n8400), .Y(n6968) );
  MUX2X1 U8259 ( .B(n6967), .A(n6952), .S(n8387), .Y(n8338) );
  MUX2X1 U8260 ( .B(ram[83]), .A(ram[19]), .S(n8508), .Y(n6972) );
  MUX2X1 U8261 ( .B(ram[211]), .A(ram[147]), .S(n8508), .Y(n6971) );
  MUX2X1 U8262 ( .B(ram[339]), .A(ram[275]), .S(n8508), .Y(n6975) );
  MUX2X1 U8263 ( .B(ram[467]), .A(ram[403]), .S(n8508), .Y(n6974) );
  MUX2X1 U8264 ( .B(n6973), .A(n6970), .S(n8401), .Y(n6984) );
  MUX2X1 U8265 ( .B(ram[595]), .A(ram[531]), .S(n8508), .Y(n6978) );
  MUX2X1 U8266 ( .B(ram[723]), .A(ram[659]), .S(n8508), .Y(n6977) );
  MUX2X1 U8267 ( .B(ram[851]), .A(ram[787]), .S(n8508), .Y(n6981) );
  MUX2X1 U8268 ( .B(ram[979]), .A(ram[915]), .S(n8508), .Y(n6980) );
  MUX2X1 U8269 ( .B(n6979), .A(n6976), .S(n8401), .Y(n6983) );
  MUX2X1 U8270 ( .B(ram[1107]), .A(ram[1043]), .S(n8508), .Y(n6987) );
  MUX2X1 U8271 ( .B(ram[1235]), .A(ram[1171]), .S(n8508), .Y(n6986) );
  MUX2X1 U8272 ( .B(ram[1363]), .A(ram[1299]), .S(n8508), .Y(n6990) );
  MUX2X1 U8273 ( .B(ram[1491]), .A(ram[1427]), .S(n8508), .Y(n6989) );
  MUX2X1 U8274 ( .B(n6988), .A(n6985), .S(n8401), .Y(n6999) );
  MUX2X1 U8275 ( .B(ram[1619]), .A(ram[1555]), .S(n8509), .Y(n6993) );
  MUX2X1 U8276 ( .B(ram[1747]), .A(ram[1683]), .S(n8509), .Y(n6992) );
  MUX2X1 U8277 ( .B(ram[1875]), .A(ram[1811]), .S(n8509), .Y(n6996) );
  MUX2X1 U8278 ( .B(ram[2003]), .A(ram[1939]), .S(n8509), .Y(n6995) );
  MUX2X1 U8279 ( .B(n6994), .A(n6991), .S(n8401), .Y(n6998) );
  MUX2X1 U8280 ( .B(n6997), .A(n6982), .S(n8387), .Y(n8339) );
  MUX2X1 U8281 ( .B(ram[84]), .A(ram[20]), .S(n8509), .Y(n7002) );
  MUX2X1 U8282 ( .B(ram[212]), .A(ram[148]), .S(n8509), .Y(n7001) );
  MUX2X1 U8283 ( .B(ram[340]), .A(ram[276]), .S(n8509), .Y(n7005) );
  MUX2X1 U8284 ( .B(ram[468]), .A(ram[404]), .S(n8509), .Y(n7004) );
  MUX2X1 U8285 ( .B(n7003), .A(n7000), .S(n8401), .Y(n7014) );
  MUX2X1 U8286 ( .B(ram[596]), .A(ram[532]), .S(n8509), .Y(n7008) );
  MUX2X1 U8287 ( .B(ram[724]), .A(ram[660]), .S(n8509), .Y(n7007) );
  MUX2X1 U8288 ( .B(ram[852]), .A(ram[788]), .S(n8509), .Y(n7011) );
  MUX2X1 U8289 ( .B(ram[980]), .A(ram[916]), .S(n8509), .Y(n7010) );
  MUX2X1 U8290 ( .B(n7009), .A(n7006), .S(n8401), .Y(n7013) );
  MUX2X1 U8291 ( .B(ram[1108]), .A(ram[1044]), .S(n8510), .Y(n7017) );
  MUX2X1 U8292 ( .B(ram[1236]), .A(ram[1172]), .S(n8510), .Y(n7016) );
  MUX2X1 U8293 ( .B(ram[1364]), .A(ram[1300]), .S(n8510), .Y(n7020) );
  MUX2X1 U8294 ( .B(ram[1492]), .A(ram[1428]), .S(n8510), .Y(n7019) );
  MUX2X1 U8295 ( .B(n7018), .A(n7015), .S(n8401), .Y(n7029) );
  MUX2X1 U8296 ( .B(ram[1620]), .A(ram[1556]), .S(n8510), .Y(n7023) );
  MUX2X1 U8297 ( .B(ram[1748]), .A(ram[1684]), .S(n8510), .Y(n7022) );
  MUX2X1 U8298 ( .B(ram[1876]), .A(ram[1812]), .S(n8510), .Y(n7026) );
  MUX2X1 U8299 ( .B(ram[2004]), .A(ram[1940]), .S(n8510), .Y(n7025) );
  MUX2X1 U8300 ( .B(n7024), .A(n7021), .S(n8401), .Y(n7028) );
  MUX2X1 U8301 ( .B(n7027), .A(n7012), .S(n8387), .Y(n8340) );
  MUX2X1 U8302 ( .B(ram[85]), .A(ram[21]), .S(n8510), .Y(n7032) );
  MUX2X1 U8303 ( .B(ram[213]), .A(ram[149]), .S(n8510), .Y(n7031) );
  MUX2X1 U8304 ( .B(ram[341]), .A(ram[277]), .S(n8510), .Y(n7035) );
  MUX2X1 U8305 ( .B(ram[469]), .A(ram[405]), .S(n8510), .Y(n7034) );
  MUX2X1 U8306 ( .B(n7033), .A(n7030), .S(n8401), .Y(n7044) );
  MUX2X1 U8307 ( .B(ram[597]), .A(ram[533]), .S(n8511), .Y(n7038) );
  MUX2X1 U8308 ( .B(ram[725]), .A(ram[661]), .S(n8511), .Y(n7037) );
  MUX2X1 U8309 ( .B(ram[853]), .A(ram[789]), .S(n8511), .Y(n7041) );
  MUX2X1 U8310 ( .B(ram[981]), .A(ram[917]), .S(n8511), .Y(n7040) );
  MUX2X1 U8311 ( .B(n7039), .A(n7036), .S(n8401), .Y(n7043) );
  MUX2X1 U8312 ( .B(ram[1109]), .A(ram[1045]), .S(n8511), .Y(n7047) );
  MUX2X1 U8313 ( .B(ram[1237]), .A(ram[1173]), .S(n8511), .Y(n7046) );
  MUX2X1 U8314 ( .B(ram[1365]), .A(ram[1301]), .S(n8511), .Y(n7050) );
  MUX2X1 U8315 ( .B(ram[1493]), .A(ram[1429]), .S(n8511), .Y(n7049) );
  MUX2X1 U8316 ( .B(n7048), .A(n7045), .S(n8401), .Y(n7059) );
  MUX2X1 U8317 ( .B(ram[1621]), .A(ram[1557]), .S(n8511), .Y(n7053) );
  MUX2X1 U8318 ( .B(ram[1749]), .A(ram[1685]), .S(n8511), .Y(n7052) );
  MUX2X1 U8319 ( .B(ram[1877]), .A(ram[1813]), .S(n8511), .Y(n7056) );
  MUX2X1 U8320 ( .B(ram[2005]), .A(ram[1941]), .S(n8511), .Y(n7055) );
  MUX2X1 U8321 ( .B(n7054), .A(n7051), .S(n8401), .Y(n7058) );
  MUX2X1 U8322 ( .B(n7057), .A(n7042), .S(n8387), .Y(n8341) );
  MUX2X1 U8323 ( .B(ram[86]), .A(ram[22]), .S(n8512), .Y(n7062) );
  MUX2X1 U8324 ( .B(ram[214]), .A(ram[150]), .S(n8512), .Y(n7061) );
  MUX2X1 U8325 ( .B(ram[342]), .A(ram[278]), .S(n8512), .Y(n7065) );
  MUX2X1 U8326 ( .B(ram[470]), .A(ram[406]), .S(n8512), .Y(n7064) );
  MUX2X1 U8327 ( .B(n7063), .A(n7060), .S(n8405), .Y(n7074) );
  MUX2X1 U8328 ( .B(ram[598]), .A(ram[534]), .S(n8512), .Y(n7068) );
  MUX2X1 U8329 ( .B(ram[726]), .A(ram[662]), .S(n8512), .Y(n7067) );
  MUX2X1 U8330 ( .B(ram[854]), .A(ram[790]), .S(n8512), .Y(n7071) );
  MUX2X1 U8331 ( .B(ram[982]), .A(ram[918]), .S(n8512), .Y(n7070) );
  MUX2X1 U8332 ( .B(n7069), .A(n7066), .S(n8406), .Y(n7073) );
  MUX2X1 U8333 ( .B(ram[1110]), .A(ram[1046]), .S(n8512), .Y(n7077) );
  MUX2X1 U8334 ( .B(ram[1238]), .A(ram[1174]), .S(n8512), .Y(n7076) );
  MUX2X1 U8335 ( .B(ram[1366]), .A(ram[1302]), .S(n8512), .Y(n7080) );
  MUX2X1 U8336 ( .B(ram[1494]), .A(ram[1430]), .S(n8512), .Y(n7079) );
  MUX2X1 U8337 ( .B(n7078), .A(n7075), .S(n8407), .Y(n7089) );
  MUX2X1 U8338 ( .B(ram[1622]), .A(ram[1558]), .S(n8513), .Y(n7083) );
  MUX2X1 U8339 ( .B(ram[1750]), .A(ram[1686]), .S(n8513), .Y(n7082) );
  MUX2X1 U8340 ( .B(ram[1878]), .A(ram[1814]), .S(n8513), .Y(n7086) );
  MUX2X1 U8341 ( .B(ram[2006]), .A(ram[1942]), .S(n8513), .Y(n7085) );
  MUX2X1 U8342 ( .B(n7084), .A(n7081), .S(n8410), .Y(n7088) );
  MUX2X1 U8343 ( .B(n7087), .A(n7072), .S(n8387), .Y(n8342) );
  MUX2X1 U8344 ( .B(ram[87]), .A(ram[23]), .S(n8513), .Y(n7092) );
  MUX2X1 U8345 ( .B(ram[215]), .A(ram[151]), .S(n8513), .Y(n7091) );
  MUX2X1 U8346 ( .B(ram[343]), .A(ram[279]), .S(n8513), .Y(n7095) );
  MUX2X1 U8347 ( .B(ram[471]), .A(ram[407]), .S(n8513), .Y(n7094) );
  MUX2X1 U8348 ( .B(n7093), .A(n7090), .S(n8409), .Y(n7104) );
  MUX2X1 U8349 ( .B(ram[599]), .A(ram[535]), .S(n8513), .Y(n7098) );
  MUX2X1 U8350 ( .B(ram[727]), .A(ram[663]), .S(n8513), .Y(n7097) );
  MUX2X1 U8351 ( .B(ram[855]), .A(ram[791]), .S(n8513), .Y(n7101) );
  MUX2X1 U8352 ( .B(ram[983]), .A(ram[919]), .S(n8513), .Y(n7100) );
  MUX2X1 U8353 ( .B(n7099), .A(n7096), .S(n8398), .Y(n7103) );
  MUX2X1 U8354 ( .B(ram[1111]), .A(ram[1047]), .S(n8514), .Y(n7107) );
  MUX2X1 U8355 ( .B(ram[1239]), .A(ram[1175]), .S(n8514), .Y(n7106) );
  MUX2X1 U8356 ( .B(ram[1367]), .A(ram[1303]), .S(n8514), .Y(n7110) );
  MUX2X1 U8357 ( .B(ram[1495]), .A(ram[1431]), .S(n8514), .Y(n7109) );
  MUX2X1 U8358 ( .B(n7108), .A(n7105), .S(n8408), .Y(n7119) );
  MUX2X1 U8359 ( .B(ram[1623]), .A(ram[1559]), .S(n8514), .Y(n7113) );
  MUX2X1 U8360 ( .B(ram[1751]), .A(ram[1687]), .S(n8514), .Y(n7112) );
  MUX2X1 U8361 ( .B(ram[1879]), .A(ram[1815]), .S(n8514), .Y(n7116) );
  MUX2X1 U8362 ( .B(ram[2007]), .A(ram[1943]), .S(n8514), .Y(n7115) );
  MUX2X1 U8363 ( .B(n7114), .A(n7111), .S(n8397), .Y(n7118) );
  MUX2X1 U8364 ( .B(n7117), .A(n7102), .S(n8387), .Y(n8343) );
  MUX2X1 U8365 ( .B(ram[88]), .A(ram[24]), .S(n8514), .Y(n7122) );
  MUX2X1 U8366 ( .B(ram[216]), .A(ram[152]), .S(n8514), .Y(n7121) );
  MUX2X1 U8367 ( .B(ram[344]), .A(ram[280]), .S(n8514), .Y(n7125) );
  MUX2X1 U8368 ( .B(ram[472]), .A(ram[408]), .S(n8514), .Y(n7124) );
  MUX2X1 U8369 ( .B(n7123), .A(n7120), .S(n8409), .Y(n7134) );
  MUX2X1 U8370 ( .B(ram[600]), .A(ram[536]), .S(n8515), .Y(n7128) );
  MUX2X1 U8371 ( .B(ram[728]), .A(ram[664]), .S(n8515), .Y(n7127) );
  MUX2X1 U8372 ( .B(ram[856]), .A(ram[792]), .S(n8515), .Y(n7131) );
  MUX2X1 U8373 ( .B(ram[984]), .A(ram[920]), .S(n8515), .Y(n7130) );
  MUX2X1 U8374 ( .B(n7129), .A(n7126), .S(n8398), .Y(n7133) );
  MUX2X1 U8375 ( .B(ram[1112]), .A(ram[1048]), .S(n8515), .Y(n7137) );
  MUX2X1 U8376 ( .B(ram[1240]), .A(ram[1176]), .S(n8515), .Y(n7136) );
  MUX2X1 U8377 ( .B(ram[1368]), .A(ram[1304]), .S(n8515), .Y(n7140) );
  MUX2X1 U8378 ( .B(ram[1496]), .A(ram[1432]), .S(n8515), .Y(n7139) );
  MUX2X1 U8379 ( .B(n7138), .A(n7135), .S(n8407), .Y(n7149) );
  MUX2X1 U8380 ( .B(ram[1624]), .A(ram[1560]), .S(n8515), .Y(n7143) );
  MUX2X1 U8381 ( .B(ram[1752]), .A(ram[1688]), .S(n8515), .Y(n7142) );
  MUX2X1 U8382 ( .B(ram[1880]), .A(ram[1816]), .S(n8515), .Y(n7146) );
  MUX2X1 U8383 ( .B(ram[2008]), .A(ram[1944]), .S(n8515), .Y(n7145) );
  MUX2X1 U8384 ( .B(n7144), .A(n7141), .S(n8405), .Y(n7148) );
  MUX2X1 U8385 ( .B(n7147), .A(n7132), .S(n8385), .Y(n8344) );
  MUX2X1 U8386 ( .B(ram[89]), .A(ram[25]), .S(n8516), .Y(n7152) );
  MUX2X1 U8387 ( .B(ram[217]), .A(ram[153]), .S(n8516), .Y(n7151) );
  MUX2X1 U8388 ( .B(ram[345]), .A(ram[281]), .S(n8516), .Y(n7155) );
  MUX2X1 U8389 ( .B(ram[473]), .A(ram[409]), .S(n8516), .Y(n7154) );
  MUX2X1 U8390 ( .B(n7153), .A(n7150), .S(n8405), .Y(n7164) );
  MUX2X1 U8391 ( .B(ram[601]), .A(ram[537]), .S(n8516), .Y(n7158) );
  MUX2X1 U8392 ( .B(ram[729]), .A(ram[665]), .S(n8516), .Y(n7157) );
  MUX2X1 U8393 ( .B(ram[857]), .A(ram[793]), .S(n8516), .Y(n7161) );
  MUX2X1 U8394 ( .B(ram[985]), .A(ram[921]), .S(n8516), .Y(n7160) );
  MUX2X1 U8395 ( .B(n7159), .A(n7156), .S(n8408), .Y(n7163) );
  MUX2X1 U8396 ( .B(ram[1113]), .A(ram[1049]), .S(n8516), .Y(n7167) );
  MUX2X1 U8397 ( .B(ram[1241]), .A(ram[1177]), .S(n8516), .Y(n7166) );
  MUX2X1 U8398 ( .B(ram[1369]), .A(ram[1305]), .S(n8516), .Y(n7170) );
  MUX2X1 U8399 ( .B(ram[1497]), .A(ram[1433]), .S(n8516), .Y(n7169) );
  MUX2X1 U8400 ( .B(n7168), .A(n7165), .S(n8410), .Y(n7179) );
  MUX2X1 U8401 ( .B(ram[1625]), .A(ram[1561]), .S(n8517), .Y(n7173) );
  MUX2X1 U8402 ( .B(ram[1753]), .A(ram[1689]), .S(n8517), .Y(n7172) );
  MUX2X1 U8403 ( .B(ram[1881]), .A(ram[1817]), .S(n8517), .Y(n7176) );
  MUX2X1 U8404 ( .B(ram[2009]), .A(ram[1945]), .S(n8517), .Y(n7175) );
  MUX2X1 U8405 ( .B(n7174), .A(n7171), .S(n8409), .Y(n7178) );
  MUX2X1 U8406 ( .B(n7177), .A(n7162), .S(n8387), .Y(n8345) );
  MUX2X1 U8407 ( .B(ram[90]), .A(ram[26]), .S(n8517), .Y(n7182) );
  MUX2X1 U8408 ( .B(ram[218]), .A(ram[154]), .S(n8517), .Y(n7181) );
  MUX2X1 U8409 ( .B(ram[346]), .A(ram[282]), .S(n8517), .Y(n7185) );
  MUX2X1 U8410 ( .B(ram[474]), .A(ram[410]), .S(n8517), .Y(n7184) );
  MUX2X1 U8411 ( .B(n7183), .A(n7180), .S(n8398), .Y(n7194) );
  MUX2X1 U8412 ( .B(ram[602]), .A(ram[538]), .S(n8517), .Y(n7188) );
  MUX2X1 U8413 ( .B(ram[730]), .A(ram[666]), .S(n8517), .Y(n7187) );
  MUX2X1 U8414 ( .B(ram[858]), .A(ram[794]), .S(n8517), .Y(n7191) );
  MUX2X1 U8415 ( .B(ram[986]), .A(ram[922]), .S(n8517), .Y(n7190) );
  MUX2X1 U8416 ( .B(n7189), .A(n7186), .S(n8408), .Y(n7193) );
  MUX2X1 U8417 ( .B(ram[1114]), .A(ram[1050]), .S(n8518), .Y(n7197) );
  MUX2X1 U8418 ( .B(ram[1242]), .A(ram[1178]), .S(n8518), .Y(n7196) );
  MUX2X1 U8419 ( .B(ram[1370]), .A(ram[1306]), .S(n8518), .Y(n7200) );
  MUX2X1 U8420 ( .B(ram[1498]), .A(ram[1434]), .S(n8518), .Y(n7199) );
  MUX2X1 U8421 ( .B(n7198), .A(n7195), .S(n8407), .Y(n7209) );
  MUX2X1 U8422 ( .B(ram[1626]), .A(ram[1562]), .S(n8518), .Y(n7203) );
  MUX2X1 U8423 ( .B(ram[1754]), .A(ram[1690]), .S(n8518), .Y(n7202) );
  MUX2X1 U8424 ( .B(ram[1882]), .A(ram[1818]), .S(n8518), .Y(n7206) );
  MUX2X1 U8425 ( .B(ram[2010]), .A(ram[1946]), .S(n8518), .Y(n7205) );
  MUX2X1 U8426 ( .B(n7204), .A(n7201), .S(n8409), .Y(n7208) );
  MUX2X1 U8427 ( .B(n7207), .A(n7192), .S(n8387), .Y(n8346) );
  MUX2X1 U8428 ( .B(ram[91]), .A(ram[27]), .S(n8518), .Y(n7212) );
  MUX2X1 U8429 ( .B(ram[219]), .A(ram[155]), .S(n8518), .Y(n7211) );
  MUX2X1 U8430 ( .B(ram[347]), .A(ram[283]), .S(n8518), .Y(n7215) );
  MUX2X1 U8431 ( .B(ram[475]), .A(ram[411]), .S(n8518), .Y(n7214) );
  MUX2X1 U8432 ( .B(n7213), .A(n7210), .S(n8405), .Y(n7224) );
  MUX2X1 U8433 ( .B(ram[603]), .A(ram[539]), .S(n8519), .Y(n7218) );
  MUX2X1 U8434 ( .B(ram[731]), .A(ram[667]), .S(n8519), .Y(n7217) );
  MUX2X1 U8435 ( .B(ram[859]), .A(ram[795]), .S(n8519), .Y(n7221) );
  MUX2X1 U8436 ( .B(ram[987]), .A(ram[923]), .S(n8519), .Y(n7220) );
  MUX2X1 U8437 ( .B(n7219), .A(n7216), .S(n8410), .Y(n7223) );
  MUX2X1 U8438 ( .B(ram[1115]), .A(ram[1051]), .S(n8519), .Y(n7227) );
  MUX2X1 U8439 ( .B(ram[1243]), .A(ram[1179]), .S(n8519), .Y(n7226) );
  MUX2X1 U8440 ( .B(ram[1371]), .A(ram[1307]), .S(n8519), .Y(n7230) );
  MUX2X1 U8441 ( .B(ram[1499]), .A(ram[1435]), .S(n8519), .Y(n7229) );
  MUX2X1 U8442 ( .B(n7228), .A(n7225), .S(n8398), .Y(n7239) );
  MUX2X1 U8443 ( .B(ram[1627]), .A(ram[1563]), .S(n8519), .Y(n7233) );
  MUX2X1 U8444 ( .B(ram[1755]), .A(ram[1691]), .S(n8519), .Y(n7232) );
  MUX2X1 U8445 ( .B(ram[1883]), .A(ram[1819]), .S(n8519), .Y(n7236) );
  MUX2X1 U8446 ( .B(ram[2011]), .A(ram[1947]), .S(n8519), .Y(n7235) );
  MUX2X1 U8447 ( .B(n7234), .A(n7231), .S(n8408), .Y(n7238) );
  MUX2X1 U8448 ( .B(n7237), .A(n7222), .S(n8386), .Y(n8347) );
  MUX2X1 U8449 ( .B(ram[92]), .A(ram[28]), .S(n8520), .Y(n7242) );
  MUX2X1 U8450 ( .B(ram[220]), .A(ram[156]), .S(n8520), .Y(n7241) );
  MUX2X1 U8451 ( .B(ram[348]), .A(ram[284]), .S(n8520), .Y(n7245) );
  MUX2X1 U8452 ( .B(ram[476]), .A(ram[412]), .S(n8520), .Y(n7244) );
  MUX2X1 U8453 ( .B(n7243), .A(n7240), .S(n8402), .Y(n7254) );
  MUX2X1 U8454 ( .B(ram[604]), .A(ram[540]), .S(n8520), .Y(n7248) );
  MUX2X1 U8455 ( .B(ram[732]), .A(ram[668]), .S(n8520), .Y(n7247) );
  MUX2X1 U8456 ( .B(ram[860]), .A(ram[796]), .S(n8520), .Y(n7251) );
  MUX2X1 U8457 ( .B(ram[988]), .A(ram[924]), .S(n8520), .Y(n7250) );
  MUX2X1 U8458 ( .B(n7249), .A(n7246), .S(n8402), .Y(n7253) );
  MUX2X1 U8459 ( .B(ram[1116]), .A(ram[1052]), .S(n8520), .Y(n7257) );
  MUX2X1 U8460 ( .B(ram[1244]), .A(ram[1180]), .S(n8520), .Y(n7256) );
  MUX2X1 U8461 ( .B(ram[1372]), .A(ram[1308]), .S(n8520), .Y(n7260) );
  MUX2X1 U8462 ( .B(ram[1500]), .A(ram[1436]), .S(n8520), .Y(n7259) );
  MUX2X1 U8463 ( .B(n7258), .A(n7255), .S(n8402), .Y(n7269) );
  MUX2X1 U8464 ( .B(ram[1628]), .A(ram[1564]), .S(n8521), .Y(n7263) );
  MUX2X1 U8465 ( .B(ram[1756]), .A(ram[1692]), .S(n8521), .Y(n7262) );
  MUX2X1 U8466 ( .B(ram[1884]), .A(ram[1820]), .S(n8521), .Y(n7266) );
  MUX2X1 U8467 ( .B(ram[2012]), .A(ram[1948]), .S(n8521), .Y(n7265) );
  MUX2X1 U8468 ( .B(n7264), .A(n7261), .S(n8402), .Y(n7268) );
  MUX2X1 U8469 ( .B(n7267), .A(n7252), .S(n8386), .Y(n8348) );
  MUX2X1 U8470 ( .B(ram[93]), .A(ram[29]), .S(n8521), .Y(n7272) );
  MUX2X1 U8471 ( .B(ram[221]), .A(ram[157]), .S(n8521), .Y(n7271) );
  MUX2X1 U8472 ( .B(ram[349]), .A(ram[285]), .S(n8521), .Y(n7275) );
  MUX2X1 U8473 ( .B(ram[477]), .A(ram[413]), .S(n8521), .Y(n7274) );
  MUX2X1 U8474 ( .B(n7273), .A(n7270), .S(n8402), .Y(n7284) );
  MUX2X1 U8475 ( .B(ram[605]), .A(ram[541]), .S(n8521), .Y(n7278) );
  MUX2X1 U8476 ( .B(ram[733]), .A(ram[669]), .S(n8521), .Y(n7277) );
  MUX2X1 U8477 ( .B(ram[861]), .A(ram[797]), .S(n8521), .Y(n7281) );
  MUX2X1 U8478 ( .B(ram[989]), .A(ram[925]), .S(n8521), .Y(n7280) );
  MUX2X1 U8479 ( .B(n7279), .A(n7276), .S(n8402), .Y(n7283) );
  MUX2X1 U8480 ( .B(ram[1117]), .A(ram[1053]), .S(n8522), .Y(n7287) );
  MUX2X1 U8481 ( .B(ram[1245]), .A(ram[1181]), .S(n8522), .Y(n7286) );
  MUX2X1 U8482 ( .B(ram[1373]), .A(ram[1309]), .S(n8522), .Y(n7290) );
  MUX2X1 U8483 ( .B(ram[1501]), .A(ram[1437]), .S(n8522), .Y(n7289) );
  MUX2X1 U8484 ( .B(n7288), .A(n7285), .S(n8402), .Y(n7299) );
  MUX2X1 U8485 ( .B(ram[1629]), .A(ram[1565]), .S(n8522), .Y(n7293) );
  MUX2X1 U8486 ( .B(ram[1757]), .A(ram[1693]), .S(n8522), .Y(n7292) );
  MUX2X1 U8487 ( .B(ram[1885]), .A(ram[1821]), .S(n8522), .Y(n7296) );
  MUX2X1 U8488 ( .B(ram[2013]), .A(ram[1949]), .S(n8522), .Y(n7295) );
  MUX2X1 U8489 ( .B(n7294), .A(n7291), .S(n8402), .Y(n7298) );
  MUX2X1 U8490 ( .B(n7297), .A(n7282), .S(n8385), .Y(n8349) );
  MUX2X1 U8491 ( .B(ram[94]), .A(ram[30]), .S(n8522), .Y(n7302) );
  MUX2X1 U8492 ( .B(ram[222]), .A(ram[158]), .S(n8522), .Y(n7301) );
  MUX2X1 U8493 ( .B(ram[350]), .A(ram[286]), .S(n8522), .Y(n7305) );
  MUX2X1 U8494 ( .B(ram[478]), .A(ram[414]), .S(n8522), .Y(n7304) );
  MUX2X1 U8495 ( .B(n7303), .A(n7300), .S(n8402), .Y(n7314) );
  MUX2X1 U8496 ( .B(ram[606]), .A(ram[542]), .S(n8523), .Y(n7308) );
  MUX2X1 U8497 ( .B(ram[734]), .A(ram[670]), .S(n8523), .Y(n7307) );
  MUX2X1 U8498 ( .B(ram[862]), .A(ram[798]), .S(n8523), .Y(n7311) );
  MUX2X1 U8499 ( .B(ram[990]), .A(ram[926]), .S(n8523), .Y(n7310) );
  MUX2X1 U8500 ( .B(n7309), .A(n7306), .S(n8402), .Y(n7313) );
  MUX2X1 U8501 ( .B(ram[1118]), .A(ram[1054]), .S(n8523), .Y(n7317) );
  MUX2X1 U8502 ( .B(ram[1246]), .A(ram[1182]), .S(n8523), .Y(n7316) );
  MUX2X1 U8503 ( .B(ram[1374]), .A(ram[1310]), .S(n8523), .Y(n7320) );
  MUX2X1 U8504 ( .B(ram[1502]), .A(ram[1438]), .S(n8523), .Y(n7319) );
  MUX2X1 U8505 ( .B(n7318), .A(n7315), .S(n8402), .Y(n7329) );
  MUX2X1 U8506 ( .B(ram[1630]), .A(ram[1566]), .S(n8523), .Y(n7323) );
  MUX2X1 U8507 ( .B(ram[1758]), .A(ram[1694]), .S(n8523), .Y(n7322) );
  MUX2X1 U8508 ( .B(ram[1886]), .A(ram[1822]), .S(n8523), .Y(n7326) );
  MUX2X1 U8509 ( .B(ram[2014]), .A(ram[1950]), .S(n8523), .Y(n7325) );
  MUX2X1 U8510 ( .B(n7324), .A(n7321), .S(n8402), .Y(n7328) );
  MUX2X1 U8511 ( .B(n7327), .A(n7312), .S(n8386), .Y(n8350) );
  MUX2X1 U8512 ( .B(ram[95]), .A(ram[31]), .S(n8524), .Y(n7332) );
  MUX2X1 U8513 ( .B(ram[223]), .A(ram[159]), .S(n8524), .Y(n7331) );
  MUX2X1 U8514 ( .B(ram[351]), .A(ram[287]), .S(n8524), .Y(n7335) );
  MUX2X1 U8515 ( .B(ram[479]), .A(ram[415]), .S(n8524), .Y(n7334) );
  MUX2X1 U8516 ( .B(n7333), .A(n7330), .S(n8403), .Y(n7344) );
  MUX2X1 U8517 ( .B(ram[607]), .A(ram[543]), .S(n8524), .Y(n7338) );
  MUX2X1 U8518 ( .B(ram[735]), .A(ram[671]), .S(n8524), .Y(n7337) );
  MUX2X1 U8519 ( .B(ram[863]), .A(ram[799]), .S(n8524), .Y(n7341) );
  MUX2X1 U8520 ( .B(ram[991]), .A(ram[927]), .S(n8524), .Y(n7340) );
  MUX2X1 U8521 ( .B(n7339), .A(n7336), .S(n8403), .Y(n7343) );
  MUX2X1 U8522 ( .B(ram[1119]), .A(ram[1055]), .S(n8524), .Y(n7347) );
  MUX2X1 U8523 ( .B(ram[1247]), .A(ram[1183]), .S(n8524), .Y(n7346) );
  MUX2X1 U8524 ( .B(ram[1375]), .A(ram[1311]), .S(n8524), .Y(n7350) );
  MUX2X1 U8525 ( .B(ram[1503]), .A(ram[1439]), .S(n8524), .Y(n7349) );
  MUX2X1 U8526 ( .B(n7348), .A(n7345), .S(n8403), .Y(n7359) );
  MUX2X1 U8527 ( .B(ram[1631]), .A(ram[1567]), .S(n8525), .Y(n7353) );
  MUX2X1 U8528 ( .B(ram[1759]), .A(ram[1695]), .S(n8525), .Y(n7352) );
  MUX2X1 U8529 ( .B(ram[1887]), .A(ram[1823]), .S(n8525), .Y(n7356) );
  MUX2X1 U8530 ( .B(ram[2015]), .A(ram[1951]), .S(n8525), .Y(n7355) );
  MUX2X1 U8531 ( .B(n7354), .A(n7351), .S(n8403), .Y(n7358) );
  MUX2X1 U8532 ( .B(n7357), .A(n7342), .S(n8386), .Y(n8351) );
  MUX2X1 U8533 ( .B(ram[96]), .A(ram[32]), .S(n8525), .Y(n7362) );
  MUX2X1 U8534 ( .B(ram[224]), .A(ram[160]), .S(n8525), .Y(n7361) );
  MUX2X1 U8535 ( .B(ram[352]), .A(ram[288]), .S(n8525), .Y(n7365) );
  MUX2X1 U8536 ( .B(ram[480]), .A(ram[416]), .S(n8525), .Y(n7364) );
  MUX2X1 U8537 ( .B(n7363), .A(n7360), .S(n8403), .Y(n7374) );
  MUX2X1 U8538 ( .B(ram[608]), .A(ram[544]), .S(n8525), .Y(n7368) );
  MUX2X1 U8539 ( .B(ram[736]), .A(ram[672]), .S(n8525), .Y(n7367) );
  MUX2X1 U8540 ( .B(ram[864]), .A(ram[800]), .S(n8525), .Y(n7371) );
  MUX2X1 U8541 ( .B(ram[992]), .A(ram[928]), .S(n8525), .Y(n7370) );
  MUX2X1 U8542 ( .B(n7369), .A(n7366), .S(n8403), .Y(n7373) );
  MUX2X1 U8543 ( .B(ram[1120]), .A(ram[1056]), .S(n8526), .Y(n7377) );
  MUX2X1 U8544 ( .B(ram[1248]), .A(ram[1184]), .S(n8526), .Y(n7376) );
  MUX2X1 U8545 ( .B(ram[1376]), .A(ram[1312]), .S(n8526), .Y(n7380) );
  MUX2X1 U8546 ( .B(ram[1504]), .A(ram[1440]), .S(n8526), .Y(n7379) );
  MUX2X1 U8547 ( .B(n7378), .A(n7375), .S(n8403), .Y(n7389) );
  MUX2X1 U8548 ( .B(ram[1632]), .A(ram[1568]), .S(n8526), .Y(n7383) );
  MUX2X1 U8549 ( .B(ram[1760]), .A(ram[1696]), .S(n8526), .Y(n7382) );
  MUX2X1 U8550 ( .B(ram[1888]), .A(ram[1824]), .S(n8526), .Y(n7386) );
  MUX2X1 U8551 ( .B(ram[2016]), .A(ram[1952]), .S(n8526), .Y(n7385) );
  MUX2X1 U8552 ( .B(n7384), .A(n7381), .S(n8403), .Y(n7388) );
  MUX2X1 U8553 ( .B(n7387), .A(n7372), .S(n8385), .Y(n8352) );
  MUX2X1 U8554 ( .B(ram[97]), .A(ram[33]), .S(n8526), .Y(n7392) );
  MUX2X1 U8555 ( .B(ram[225]), .A(ram[161]), .S(n8526), .Y(n7391) );
  MUX2X1 U8556 ( .B(ram[353]), .A(ram[289]), .S(n8526), .Y(n7395) );
  MUX2X1 U8557 ( .B(ram[481]), .A(ram[417]), .S(n8526), .Y(n7394) );
  MUX2X1 U8558 ( .B(n7393), .A(n7390), .S(n8403), .Y(n7404) );
  MUX2X1 U8559 ( .B(ram[609]), .A(ram[545]), .S(n8527), .Y(n7398) );
  MUX2X1 U8560 ( .B(ram[737]), .A(ram[673]), .S(n8527), .Y(n7397) );
  MUX2X1 U8561 ( .B(ram[865]), .A(ram[801]), .S(n8527), .Y(n7401) );
  MUX2X1 U8562 ( .B(ram[993]), .A(ram[929]), .S(n8527), .Y(n7400) );
  MUX2X1 U8563 ( .B(n7399), .A(n7396), .S(n8403), .Y(n7403) );
  MUX2X1 U8564 ( .B(ram[1121]), .A(ram[1057]), .S(n8527), .Y(n7407) );
  MUX2X1 U8565 ( .B(ram[1249]), .A(ram[1185]), .S(n8527), .Y(n7406) );
  MUX2X1 U8566 ( .B(ram[1377]), .A(ram[1313]), .S(n8527), .Y(n7410) );
  MUX2X1 U8567 ( .B(ram[1505]), .A(ram[1441]), .S(n8527), .Y(n7409) );
  MUX2X1 U8568 ( .B(n7408), .A(n7405), .S(n8403), .Y(n7419) );
  MUX2X1 U8569 ( .B(ram[1633]), .A(ram[1569]), .S(n8527), .Y(n7413) );
  MUX2X1 U8570 ( .B(ram[1761]), .A(ram[1697]), .S(n8527), .Y(n7412) );
  MUX2X1 U8571 ( .B(ram[1889]), .A(ram[1825]), .S(n8527), .Y(n7416) );
  MUX2X1 U8572 ( .B(ram[2017]), .A(ram[1953]), .S(n8527), .Y(n7415) );
  MUX2X1 U8573 ( .B(n7414), .A(n7411), .S(n8403), .Y(n7418) );
  MUX2X1 U8574 ( .B(n7417), .A(n7402), .S(n8387), .Y(n8353) );
  MUX2X1 U8575 ( .B(ram[98]), .A(ram[34]), .S(n8528), .Y(n7422) );
  MUX2X1 U8576 ( .B(ram[226]), .A(ram[162]), .S(n8528), .Y(n7421) );
  MUX2X1 U8577 ( .B(ram[354]), .A(ram[290]), .S(n8528), .Y(n7425) );
  MUX2X1 U8578 ( .B(ram[482]), .A(ram[418]), .S(n8528), .Y(n7424) );
  MUX2X1 U8579 ( .B(n7423), .A(n7420), .S(n8404), .Y(n7434) );
  MUX2X1 U8580 ( .B(ram[610]), .A(ram[546]), .S(n8528), .Y(n7428) );
  MUX2X1 U8581 ( .B(ram[738]), .A(ram[674]), .S(n8528), .Y(n7427) );
  MUX2X1 U8582 ( .B(ram[866]), .A(ram[802]), .S(n8528), .Y(n7431) );
  MUX2X1 U8583 ( .B(ram[994]), .A(ram[930]), .S(n8528), .Y(n7430) );
  MUX2X1 U8584 ( .B(n7429), .A(n7426), .S(n8404), .Y(n7433) );
  MUX2X1 U8585 ( .B(ram[1122]), .A(ram[1058]), .S(n8528), .Y(n7437) );
  MUX2X1 U8586 ( .B(ram[1250]), .A(ram[1186]), .S(n8528), .Y(n7436) );
  MUX2X1 U8587 ( .B(ram[1378]), .A(ram[1314]), .S(n8528), .Y(n7440) );
  MUX2X1 U8588 ( .B(ram[1506]), .A(ram[1442]), .S(n8528), .Y(n7439) );
  MUX2X1 U8589 ( .B(n7438), .A(n7435), .S(n8404), .Y(n7449) );
  MUX2X1 U8590 ( .B(ram[1634]), .A(ram[1570]), .S(n8529), .Y(n7443) );
  MUX2X1 U8591 ( .B(ram[1762]), .A(ram[1698]), .S(n8529), .Y(n7442) );
  MUX2X1 U8592 ( .B(ram[1890]), .A(ram[1826]), .S(n8529), .Y(n7446) );
  MUX2X1 U8593 ( .B(ram[2018]), .A(ram[1954]), .S(n8529), .Y(n7445) );
  MUX2X1 U8594 ( .B(n7444), .A(n7441), .S(n8404), .Y(n7448) );
  MUX2X1 U8595 ( .B(n7447), .A(n7432), .S(n8385), .Y(n8354) );
  MUX2X1 U8596 ( .B(ram[99]), .A(ram[35]), .S(n8529), .Y(n7452) );
  MUX2X1 U8597 ( .B(ram[227]), .A(ram[163]), .S(n8529), .Y(n7451) );
  MUX2X1 U8598 ( .B(ram[355]), .A(ram[291]), .S(n8529), .Y(n7455) );
  MUX2X1 U8599 ( .B(ram[483]), .A(ram[419]), .S(n8529), .Y(n7454) );
  MUX2X1 U8600 ( .B(n7453), .A(n7450), .S(n8404), .Y(n7464) );
  MUX2X1 U8601 ( .B(ram[611]), .A(ram[547]), .S(n8529), .Y(n7458) );
  MUX2X1 U8602 ( .B(ram[739]), .A(ram[675]), .S(n8529), .Y(n7457) );
  MUX2X1 U8603 ( .B(ram[867]), .A(ram[803]), .S(n8529), .Y(n7461) );
  MUX2X1 U8604 ( .B(ram[995]), .A(ram[931]), .S(n8529), .Y(n7460) );
  MUX2X1 U8605 ( .B(n7459), .A(n7456), .S(n8404), .Y(n7463) );
  MUX2X1 U8606 ( .B(ram[1123]), .A(ram[1059]), .S(n8530), .Y(n7467) );
  MUX2X1 U8607 ( .B(ram[1251]), .A(ram[1187]), .S(n8530), .Y(n7466) );
  MUX2X1 U8608 ( .B(ram[1379]), .A(ram[1315]), .S(n8530), .Y(n7470) );
  MUX2X1 U8609 ( .B(ram[1507]), .A(ram[1443]), .S(n8530), .Y(n7469) );
  MUX2X1 U8610 ( .B(n7468), .A(n7465), .S(n8404), .Y(n7479) );
  MUX2X1 U8611 ( .B(ram[1635]), .A(ram[1571]), .S(n8530), .Y(n7473) );
  MUX2X1 U8612 ( .B(ram[1763]), .A(ram[1699]), .S(n8530), .Y(n7472) );
  MUX2X1 U8613 ( .B(ram[1891]), .A(ram[1827]), .S(n8530), .Y(n7476) );
  MUX2X1 U8614 ( .B(ram[2019]), .A(ram[1955]), .S(n8530), .Y(n7475) );
  MUX2X1 U8615 ( .B(n7474), .A(n7471), .S(n8404), .Y(n7478) );
  MUX2X1 U8616 ( .B(n7477), .A(n7462), .S(n8387), .Y(n8355) );
  MUX2X1 U8617 ( .B(ram[100]), .A(ram[36]), .S(n8530), .Y(n7482) );
  MUX2X1 U8618 ( .B(ram[228]), .A(ram[164]), .S(n8530), .Y(n7481) );
  MUX2X1 U8619 ( .B(ram[356]), .A(ram[292]), .S(n8530), .Y(n7485) );
  MUX2X1 U8620 ( .B(ram[484]), .A(ram[420]), .S(n8530), .Y(n7484) );
  MUX2X1 U8621 ( .B(n7483), .A(n7480), .S(n8404), .Y(n7494) );
  MUX2X1 U8622 ( .B(ram[612]), .A(ram[548]), .S(n8531), .Y(n7488) );
  MUX2X1 U8623 ( .B(ram[740]), .A(ram[676]), .S(n8531), .Y(n7487) );
  MUX2X1 U8624 ( .B(ram[868]), .A(ram[804]), .S(n8531), .Y(n7491) );
  MUX2X1 U8625 ( .B(ram[996]), .A(ram[932]), .S(n8531), .Y(n7490) );
  MUX2X1 U8626 ( .B(n7489), .A(n7486), .S(n8404), .Y(n7493) );
  MUX2X1 U8627 ( .B(ram[1124]), .A(ram[1060]), .S(n8531), .Y(n7497) );
  MUX2X1 U8628 ( .B(ram[1252]), .A(ram[1188]), .S(n8531), .Y(n7496) );
  MUX2X1 U8629 ( .B(ram[1380]), .A(ram[1316]), .S(n8531), .Y(n7500) );
  MUX2X1 U8630 ( .B(ram[1508]), .A(ram[1444]), .S(n8531), .Y(n7499) );
  MUX2X1 U8631 ( .B(n7498), .A(n7495), .S(n8404), .Y(n7509) );
  MUX2X1 U8632 ( .B(ram[1636]), .A(ram[1572]), .S(n8531), .Y(n7503) );
  MUX2X1 U8633 ( .B(ram[1764]), .A(ram[1700]), .S(n8531), .Y(n7502) );
  MUX2X1 U8634 ( .B(ram[1892]), .A(ram[1828]), .S(n8531), .Y(n7506) );
  MUX2X1 U8635 ( .B(ram[2020]), .A(ram[1956]), .S(n8531), .Y(n7505) );
  MUX2X1 U8636 ( .B(n7504), .A(n7501), .S(n8404), .Y(n7508) );
  MUX2X1 U8637 ( .B(n7507), .A(n7492), .S(n8386), .Y(n8356) );
  MUX2X1 U8638 ( .B(ram[101]), .A(ram[37]), .S(n8532), .Y(n7512) );
  MUX2X1 U8639 ( .B(ram[229]), .A(ram[165]), .S(n8532), .Y(n7511) );
  MUX2X1 U8640 ( .B(ram[357]), .A(ram[293]), .S(n8532), .Y(n7515) );
  MUX2X1 U8641 ( .B(ram[485]), .A(ram[421]), .S(n8532), .Y(n7514) );
  MUX2X1 U8642 ( .B(n7513), .A(n7510), .S(n8405), .Y(n7524) );
  MUX2X1 U8643 ( .B(ram[613]), .A(ram[549]), .S(n8532), .Y(n7518) );
  MUX2X1 U8644 ( .B(ram[741]), .A(ram[677]), .S(n8532), .Y(n7517) );
  MUX2X1 U8645 ( .B(ram[869]), .A(ram[805]), .S(n8532), .Y(n7521) );
  MUX2X1 U8646 ( .B(ram[997]), .A(ram[933]), .S(n8532), .Y(n7520) );
  MUX2X1 U8647 ( .B(n7519), .A(n7516), .S(n8405), .Y(n7523) );
  MUX2X1 U8648 ( .B(ram[1125]), .A(ram[1061]), .S(n8532), .Y(n7527) );
  MUX2X1 U8649 ( .B(ram[1253]), .A(ram[1189]), .S(n8532), .Y(n7526) );
  MUX2X1 U8650 ( .B(ram[1381]), .A(ram[1317]), .S(n8532), .Y(n7530) );
  MUX2X1 U8651 ( .B(ram[1509]), .A(ram[1445]), .S(n8532), .Y(n7529) );
  MUX2X1 U8652 ( .B(n7528), .A(n7525), .S(n8405), .Y(n7539) );
  MUX2X1 U8653 ( .B(ram[1637]), .A(ram[1573]), .S(n8533), .Y(n7533) );
  MUX2X1 U8654 ( .B(ram[1765]), .A(ram[1701]), .S(n8533), .Y(n7532) );
  MUX2X1 U8655 ( .B(ram[1893]), .A(ram[1829]), .S(n8533), .Y(n7536) );
  MUX2X1 U8656 ( .B(ram[2021]), .A(ram[1957]), .S(n8533), .Y(n7535) );
  MUX2X1 U8657 ( .B(n7534), .A(n7531), .S(n8405), .Y(n7538) );
  MUX2X1 U8658 ( .B(n7537), .A(n7522), .S(n8386), .Y(n8357) );
  MUX2X1 U8659 ( .B(ram[102]), .A(ram[38]), .S(n8533), .Y(n7542) );
  MUX2X1 U8660 ( .B(ram[230]), .A(ram[166]), .S(n8533), .Y(n7541) );
  MUX2X1 U8661 ( .B(ram[358]), .A(ram[294]), .S(n8533), .Y(n7545) );
  MUX2X1 U8662 ( .B(ram[486]), .A(ram[422]), .S(n8533), .Y(n7544) );
  MUX2X1 U8663 ( .B(n7543), .A(n7540), .S(n8405), .Y(n7554) );
  MUX2X1 U8664 ( .B(ram[614]), .A(ram[550]), .S(n8533), .Y(n7548) );
  MUX2X1 U8665 ( .B(ram[742]), .A(ram[678]), .S(n8533), .Y(n7547) );
  MUX2X1 U8666 ( .B(ram[870]), .A(ram[806]), .S(n8533), .Y(n7551) );
  MUX2X1 U8667 ( .B(ram[998]), .A(ram[934]), .S(n8533), .Y(n7550) );
  MUX2X1 U8668 ( .B(n7549), .A(n7546), .S(n8405), .Y(n7553) );
  MUX2X1 U8669 ( .B(ram[1126]), .A(ram[1062]), .S(n8534), .Y(n7557) );
  MUX2X1 U8670 ( .B(ram[1254]), .A(ram[1190]), .S(n8534), .Y(n7556) );
  MUX2X1 U8671 ( .B(ram[1382]), .A(ram[1318]), .S(n8534), .Y(n7560) );
  MUX2X1 U8672 ( .B(ram[1510]), .A(ram[1446]), .S(n8534), .Y(n7559) );
  MUX2X1 U8673 ( .B(n7558), .A(n7555), .S(n8405), .Y(n7569) );
  MUX2X1 U8674 ( .B(ram[1638]), .A(ram[1574]), .S(n8534), .Y(n7563) );
  MUX2X1 U8675 ( .B(ram[1766]), .A(ram[1702]), .S(n8534), .Y(n7562) );
  MUX2X1 U8676 ( .B(ram[1894]), .A(ram[1830]), .S(n8534), .Y(n7566) );
  MUX2X1 U8677 ( .B(ram[2022]), .A(ram[1958]), .S(n8534), .Y(n7565) );
  MUX2X1 U8678 ( .B(n7564), .A(n7561), .S(n8405), .Y(n7568) );
  MUX2X1 U8679 ( .B(n7567), .A(n7552), .S(n8386), .Y(n8358) );
  MUX2X1 U8680 ( .B(ram[103]), .A(ram[39]), .S(n8534), .Y(n7572) );
  MUX2X1 U8681 ( .B(ram[231]), .A(ram[167]), .S(n8534), .Y(n7571) );
  MUX2X1 U8682 ( .B(ram[359]), .A(ram[295]), .S(n8534), .Y(n7575) );
  MUX2X1 U8683 ( .B(ram[487]), .A(ram[423]), .S(n8534), .Y(n7574) );
  MUX2X1 U8684 ( .B(n7573), .A(n7570), .S(n8405), .Y(n7584) );
  MUX2X1 U8685 ( .B(ram[615]), .A(ram[551]), .S(n8535), .Y(n7578) );
  MUX2X1 U8686 ( .B(ram[743]), .A(ram[679]), .S(n8535), .Y(n7577) );
  MUX2X1 U8687 ( .B(ram[871]), .A(ram[807]), .S(n8535), .Y(n7581) );
  MUX2X1 U8688 ( .B(ram[999]), .A(ram[935]), .S(n8535), .Y(n7580) );
  MUX2X1 U8689 ( .B(n7579), .A(n7576), .S(n8405), .Y(n7583) );
  MUX2X1 U8690 ( .B(ram[1127]), .A(ram[1063]), .S(n8535), .Y(n7587) );
  MUX2X1 U8691 ( .B(ram[1255]), .A(ram[1191]), .S(n8535), .Y(n7586) );
  MUX2X1 U8692 ( .B(ram[1383]), .A(ram[1319]), .S(n8535), .Y(n7590) );
  MUX2X1 U8693 ( .B(ram[1511]), .A(ram[1447]), .S(n8535), .Y(n7589) );
  MUX2X1 U8694 ( .B(n7588), .A(n7585), .S(n8405), .Y(n7599) );
  MUX2X1 U8695 ( .B(ram[1639]), .A(ram[1575]), .S(n8535), .Y(n7593) );
  MUX2X1 U8696 ( .B(ram[1767]), .A(ram[1703]), .S(n8535), .Y(n7592) );
  MUX2X1 U8697 ( .B(ram[1895]), .A(ram[1831]), .S(n8535), .Y(n7596) );
  MUX2X1 U8698 ( .B(ram[2023]), .A(ram[1959]), .S(n8535), .Y(n7595) );
  MUX2X1 U8699 ( .B(n7594), .A(n7591), .S(n8405), .Y(n7598) );
  MUX2X1 U8700 ( .B(n7597), .A(n7582), .S(n8386), .Y(n8359) );
  MUX2X1 U8701 ( .B(ram[104]), .A(ram[40]), .S(n8536), .Y(n7602) );
  MUX2X1 U8702 ( .B(ram[232]), .A(ram[168]), .S(n8536), .Y(n7601) );
  MUX2X1 U8703 ( .B(ram[360]), .A(ram[296]), .S(n8536), .Y(n7605) );
  MUX2X1 U8704 ( .B(ram[488]), .A(ram[424]), .S(n8536), .Y(n7604) );
  MUX2X1 U8705 ( .B(n7603), .A(n7600), .S(n8401), .Y(n7614) );
  MUX2X1 U8706 ( .B(ram[616]), .A(ram[552]), .S(n8536), .Y(n7608) );
  MUX2X1 U8707 ( .B(ram[744]), .A(ram[680]), .S(n8536), .Y(n7607) );
  MUX2X1 U8708 ( .B(ram[872]), .A(ram[808]), .S(n8536), .Y(n7611) );
  MUX2X1 U8709 ( .B(ram[1000]), .A(ram[936]), .S(n8536), .Y(n7610) );
  MUX2X1 U8710 ( .B(n7609), .A(n7606), .S(n8403), .Y(n7613) );
  MUX2X1 U8711 ( .B(ram[1128]), .A(ram[1064]), .S(n8536), .Y(n7617) );
  MUX2X1 U8712 ( .B(ram[1256]), .A(ram[1192]), .S(n8536), .Y(n7616) );
  MUX2X1 U8713 ( .B(ram[1384]), .A(ram[1320]), .S(n8536), .Y(n7620) );
  MUX2X1 U8714 ( .B(ram[1512]), .A(ram[1448]), .S(n8536), .Y(n7619) );
  MUX2X1 U8715 ( .B(n7618), .A(n7615), .S(n8410), .Y(n7629) );
  MUX2X1 U8716 ( .B(ram[1640]), .A(ram[1576]), .S(n8537), .Y(n7623) );
  MUX2X1 U8717 ( .B(ram[1768]), .A(ram[1704]), .S(n8537), .Y(n7622) );
  MUX2X1 U8718 ( .B(ram[1896]), .A(ram[1832]), .S(n8537), .Y(n7626) );
  MUX2X1 U8719 ( .B(ram[2024]), .A(ram[1960]), .S(n8537), .Y(n7625) );
  MUX2X1 U8720 ( .B(n7624), .A(n7621), .S(n8407), .Y(n7628) );
  MUX2X1 U8721 ( .B(n7627), .A(n7612), .S(n8386), .Y(n8360) );
  MUX2X1 U8722 ( .B(ram[105]), .A(ram[41]), .S(n8537), .Y(n7632) );
  MUX2X1 U8723 ( .B(ram[233]), .A(ram[169]), .S(n8537), .Y(n7631) );
  MUX2X1 U8724 ( .B(ram[361]), .A(ram[297]), .S(n8537), .Y(n7635) );
  MUX2X1 U8725 ( .B(ram[489]), .A(ram[425]), .S(n8537), .Y(n7634) );
  MUX2X1 U8726 ( .B(n7633), .A(n7630), .S(n8402), .Y(n7644) );
  MUX2X1 U8727 ( .B(ram[617]), .A(ram[553]), .S(n8537), .Y(n7638) );
  MUX2X1 U8728 ( .B(ram[745]), .A(ram[681]), .S(n8537), .Y(n7637) );
  MUX2X1 U8729 ( .B(ram[873]), .A(ram[809]), .S(n8537), .Y(n7641) );
  MUX2X1 U8730 ( .B(ram[1001]), .A(ram[937]), .S(n8537), .Y(n7640) );
  MUX2X1 U8731 ( .B(n7639), .A(n7636), .S(n8405), .Y(n7643) );
  MUX2X1 U8732 ( .B(ram[1129]), .A(ram[1065]), .S(n8538), .Y(n7647) );
  MUX2X1 U8733 ( .B(ram[1257]), .A(ram[1193]), .S(n8538), .Y(n7646) );
  MUX2X1 U8734 ( .B(ram[1385]), .A(ram[1321]), .S(n8538), .Y(n7650) );
  MUX2X1 U8735 ( .B(ram[1513]), .A(ram[1449]), .S(n8538), .Y(n7649) );
  MUX2X1 U8736 ( .B(n7648), .A(n7645), .S(n8408), .Y(n7659) );
  MUX2X1 U8737 ( .B(ram[1641]), .A(ram[1577]), .S(n8538), .Y(n7653) );
  MUX2X1 U8738 ( .B(ram[1769]), .A(ram[1705]), .S(n8538), .Y(n7652) );
  MUX2X1 U8739 ( .B(ram[1897]), .A(ram[1833]), .S(n8538), .Y(n7656) );
  MUX2X1 U8740 ( .B(ram[2025]), .A(ram[1961]), .S(n8538), .Y(n7655) );
  MUX2X1 U8741 ( .B(n7654), .A(n7651), .S(n8397), .Y(n7658) );
  MUX2X1 U8742 ( .B(n7657), .A(n7642), .S(n8386), .Y(n8361) );
  MUX2X1 U8743 ( .B(ram[106]), .A(ram[42]), .S(n8538), .Y(n7662) );
  MUX2X1 U8744 ( .B(ram[234]), .A(ram[170]), .S(n8538), .Y(n7661) );
  MUX2X1 U8745 ( .B(ram[362]), .A(ram[298]), .S(n8538), .Y(n7665) );
  MUX2X1 U8746 ( .B(ram[490]), .A(ram[426]), .S(n8538), .Y(n7664) );
  MUX2X1 U8747 ( .B(n7663), .A(n7660), .S(n8399), .Y(n7674) );
  MUX2X1 U8748 ( .B(ram[618]), .A(ram[554]), .S(n8539), .Y(n7668) );
  MUX2X1 U8749 ( .B(ram[746]), .A(ram[682]), .S(n8539), .Y(n7667) );
  MUX2X1 U8750 ( .B(ram[874]), .A(ram[810]), .S(n8539), .Y(n7671) );
  MUX2X1 U8751 ( .B(ram[1002]), .A(ram[938]), .S(n8539), .Y(n7670) );
  MUX2X1 U8752 ( .B(n7669), .A(n7666), .S(n8404), .Y(n7673) );
  MUX2X1 U8753 ( .B(ram[1130]), .A(ram[1066]), .S(n8539), .Y(n7677) );
  MUX2X1 U8754 ( .B(ram[1258]), .A(ram[1194]), .S(n8539), .Y(n7676) );
  MUX2X1 U8755 ( .B(ram[1386]), .A(ram[1322]), .S(n8539), .Y(n7680) );
  MUX2X1 U8756 ( .B(ram[1514]), .A(ram[1450]), .S(n8539), .Y(n7679) );
  MUX2X1 U8757 ( .B(n7678), .A(n7675), .S(n8396), .Y(n7689) );
  MUX2X1 U8758 ( .B(ram[1642]), .A(ram[1578]), .S(n8539), .Y(n7683) );
  MUX2X1 U8759 ( .B(ram[1770]), .A(ram[1706]), .S(n8539), .Y(n7682) );
  MUX2X1 U8760 ( .B(ram[1898]), .A(ram[1834]), .S(n8539), .Y(n7686) );
  MUX2X1 U8761 ( .B(ram[2026]), .A(ram[1962]), .S(n8539), .Y(n7685) );
  MUX2X1 U8762 ( .B(n7684), .A(n7681), .S(n8406), .Y(n7688) );
  MUX2X1 U8763 ( .B(n7687), .A(n7672), .S(n8386), .Y(n8362) );
  MUX2X1 U8764 ( .B(ram[107]), .A(ram[43]), .S(n8540), .Y(n7692) );
  MUX2X1 U8765 ( .B(ram[235]), .A(ram[171]), .S(n8540), .Y(n7691) );
  MUX2X1 U8766 ( .B(ram[363]), .A(ram[299]), .S(n8540), .Y(n7695) );
  MUX2X1 U8767 ( .B(ram[491]), .A(ram[427]), .S(n8540), .Y(n7694) );
  MUX2X1 U8768 ( .B(n7693), .A(n7690), .S(n8406), .Y(n7704) );
  MUX2X1 U8769 ( .B(ram[619]), .A(ram[555]), .S(n8540), .Y(n7698) );
  MUX2X1 U8770 ( .B(ram[747]), .A(ram[683]), .S(n8540), .Y(n7697) );
  MUX2X1 U8771 ( .B(ram[875]), .A(ram[811]), .S(n8540), .Y(n7701) );
  MUX2X1 U8772 ( .B(ram[1003]), .A(ram[939]), .S(n8540), .Y(n7700) );
  MUX2X1 U8773 ( .B(n7699), .A(n7696), .S(n8406), .Y(n7703) );
  MUX2X1 U8774 ( .B(ram[1131]), .A(ram[1067]), .S(n8540), .Y(n7707) );
  MUX2X1 U8775 ( .B(ram[1259]), .A(ram[1195]), .S(n8540), .Y(n7706) );
  MUX2X1 U8776 ( .B(ram[1387]), .A(ram[1323]), .S(n8540), .Y(n7710) );
  MUX2X1 U8777 ( .B(ram[1515]), .A(ram[1451]), .S(n8540), .Y(n7709) );
  MUX2X1 U8778 ( .B(n7708), .A(n7705), .S(n8406), .Y(n7719) );
  MUX2X1 U8779 ( .B(ram[1643]), .A(ram[1579]), .S(n8541), .Y(n7713) );
  MUX2X1 U8780 ( .B(ram[1771]), .A(ram[1707]), .S(n8541), .Y(n7712) );
  MUX2X1 U8781 ( .B(ram[1899]), .A(ram[1835]), .S(n8541), .Y(n7716) );
  MUX2X1 U8782 ( .B(ram[2027]), .A(ram[1963]), .S(n8541), .Y(n7715) );
  MUX2X1 U8783 ( .B(n7714), .A(n7711), .S(n8406), .Y(n7718) );
  MUX2X1 U8784 ( .B(n7717), .A(n7702), .S(n8386), .Y(n8363) );
  MUX2X1 U8785 ( .B(ram[108]), .A(ram[44]), .S(n8541), .Y(n7722) );
  MUX2X1 U8786 ( .B(ram[236]), .A(ram[172]), .S(n8541), .Y(n7721) );
  MUX2X1 U8787 ( .B(ram[364]), .A(ram[300]), .S(n8541), .Y(n7725) );
  MUX2X1 U8788 ( .B(ram[492]), .A(ram[428]), .S(n8541), .Y(n7724) );
  MUX2X1 U8789 ( .B(n7723), .A(n7720), .S(n8406), .Y(n7734) );
  MUX2X1 U8790 ( .B(ram[620]), .A(ram[556]), .S(n8541), .Y(n7728) );
  MUX2X1 U8791 ( .B(ram[748]), .A(ram[684]), .S(n8541), .Y(n7727) );
  MUX2X1 U8792 ( .B(ram[876]), .A(ram[812]), .S(n8541), .Y(n7731) );
  MUX2X1 U8793 ( .B(ram[1004]), .A(ram[940]), .S(n8541), .Y(n7730) );
  MUX2X1 U8794 ( .B(n7729), .A(n7726), .S(n8406), .Y(n7733) );
  MUX2X1 U8795 ( .B(ram[1132]), .A(ram[1068]), .S(n8542), .Y(n7737) );
  MUX2X1 U8796 ( .B(ram[1260]), .A(ram[1196]), .S(n8542), .Y(n7736) );
  MUX2X1 U8797 ( .B(ram[1388]), .A(ram[1324]), .S(n8542), .Y(n7740) );
  MUX2X1 U8798 ( .B(ram[1516]), .A(ram[1452]), .S(n8542), .Y(n7739) );
  MUX2X1 U8799 ( .B(n7738), .A(n7735), .S(n8406), .Y(n7749) );
  MUX2X1 U8800 ( .B(ram[1644]), .A(ram[1580]), .S(n8542), .Y(n7743) );
  MUX2X1 U8801 ( .B(ram[1772]), .A(ram[1708]), .S(n8542), .Y(n7742) );
  MUX2X1 U8802 ( .B(ram[1900]), .A(ram[1836]), .S(n8542), .Y(n7746) );
  MUX2X1 U8803 ( .B(ram[2028]), .A(ram[1964]), .S(n8542), .Y(n7745) );
  MUX2X1 U8804 ( .B(n7744), .A(n7741), .S(n8406), .Y(n7748) );
  MUX2X1 U8805 ( .B(n7747), .A(n7732), .S(n8386), .Y(n8364) );
  MUX2X1 U8806 ( .B(ram[109]), .A(ram[45]), .S(n8542), .Y(n7752) );
  MUX2X1 U8807 ( .B(ram[237]), .A(ram[173]), .S(n8542), .Y(n7751) );
  MUX2X1 U8808 ( .B(ram[365]), .A(ram[301]), .S(n8542), .Y(n7755) );
  MUX2X1 U8809 ( .B(ram[493]), .A(ram[429]), .S(n8542), .Y(n7754) );
  MUX2X1 U8810 ( .B(n7753), .A(n7750), .S(n8406), .Y(n7764) );
  MUX2X1 U8811 ( .B(ram[621]), .A(ram[557]), .S(n8543), .Y(n7758) );
  MUX2X1 U8812 ( .B(ram[749]), .A(ram[685]), .S(n8543), .Y(n7757) );
  MUX2X1 U8813 ( .B(ram[877]), .A(ram[813]), .S(n8543), .Y(n7761) );
  MUX2X1 U8814 ( .B(ram[1005]), .A(ram[941]), .S(n8543), .Y(n7760) );
  MUX2X1 U8815 ( .B(n7759), .A(n7756), .S(n8406), .Y(n7763) );
  MUX2X1 U8816 ( .B(ram[1133]), .A(ram[1069]), .S(n8543), .Y(n7767) );
  MUX2X1 U8817 ( .B(ram[1261]), .A(ram[1197]), .S(n8543), .Y(n7766) );
  MUX2X1 U8818 ( .B(ram[1389]), .A(ram[1325]), .S(n8543), .Y(n7770) );
  MUX2X1 U8819 ( .B(ram[1517]), .A(ram[1453]), .S(n8543), .Y(n7769) );
  MUX2X1 U8820 ( .B(n7768), .A(n7765), .S(n8406), .Y(n7779) );
  MUX2X1 U8821 ( .B(ram[1645]), .A(ram[1581]), .S(n8543), .Y(n7773) );
  MUX2X1 U8822 ( .B(ram[1773]), .A(ram[1709]), .S(n8543), .Y(n7772) );
  MUX2X1 U8823 ( .B(ram[1901]), .A(ram[1837]), .S(n8543), .Y(n7776) );
  MUX2X1 U8824 ( .B(ram[2029]), .A(ram[1965]), .S(n8543), .Y(n7775) );
  MUX2X1 U8825 ( .B(n7774), .A(n7771), .S(n8406), .Y(n7778) );
  MUX2X1 U8826 ( .B(n7777), .A(n7762), .S(n8386), .Y(n8365) );
  MUX2X1 U8827 ( .B(ram[110]), .A(ram[46]), .S(n8544), .Y(n7782) );
  MUX2X1 U8828 ( .B(ram[238]), .A(ram[174]), .S(n8544), .Y(n7781) );
  MUX2X1 U8829 ( .B(ram[366]), .A(ram[302]), .S(n8544), .Y(n7785) );
  MUX2X1 U8830 ( .B(ram[494]), .A(ram[430]), .S(n8544), .Y(n7784) );
  MUX2X1 U8831 ( .B(n7783), .A(n7780), .S(n8407), .Y(n7794) );
  MUX2X1 U8832 ( .B(ram[622]), .A(ram[558]), .S(n8544), .Y(n7788) );
  MUX2X1 U8833 ( .B(ram[750]), .A(ram[686]), .S(n8544), .Y(n7787) );
  MUX2X1 U8834 ( .B(ram[878]), .A(ram[814]), .S(n8544), .Y(n7791) );
  MUX2X1 U8835 ( .B(ram[1006]), .A(ram[942]), .S(n8544), .Y(n7790) );
  MUX2X1 U8836 ( .B(n7789), .A(n7786), .S(n8407), .Y(n7793) );
  MUX2X1 U8837 ( .B(ram[1134]), .A(ram[1070]), .S(n8544), .Y(n7797) );
  MUX2X1 U8838 ( .B(ram[1262]), .A(ram[1198]), .S(n8544), .Y(n7796) );
  MUX2X1 U8839 ( .B(ram[1390]), .A(ram[1326]), .S(n8544), .Y(n7800) );
  MUX2X1 U8840 ( .B(ram[1518]), .A(ram[1454]), .S(n8544), .Y(n7799) );
  MUX2X1 U8841 ( .B(n7798), .A(n7795), .S(n8407), .Y(n7809) );
  MUX2X1 U8842 ( .B(ram[1646]), .A(ram[1582]), .S(n8545), .Y(n7803) );
  MUX2X1 U8843 ( .B(ram[1774]), .A(ram[1710]), .S(n8545), .Y(n7802) );
  MUX2X1 U8844 ( .B(ram[1902]), .A(ram[1838]), .S(n8545), .Y(n7806) );
  MUX2X1 U8845 ( .B(ram[2030]), .A(ram[1966]), .S(n8545), .Y(n7805) );
  MUX2X1 U8846 ( .B(n7804), .A(n7801), .S(n8407), .Y(n7808) );
  MUX2X1 U8847 ( .B(n7807), .A(n7792), .S(n8386), .Y(n8366) );
  MUX2X1 U8848 ( .B(ram[111]), .A(ram[47]), .S(n8545), .Y(n7812) );
  MUX2X1 U8849 ( .B(ram[239]), .A(ram[175]), .S(n8545), .Y(n7811) );
  MUX2X1 U8850 ( .B(ram[367]), .A(ram[303]), .S(n8545), .Y(n7815) );
  MUX2X1 U8851 ( .B(ram[495]), .A(ram[431]), .S(n8545), .Y(n7814) );
  MUX2X1 U8852 ( .B(n7813), .A(n7810), .S(n8407), .Y(n7824) );
  MUX2X1 U8853 ( .B(ram[623]), .A(ram[559]), .S(n8545), .Y(n7818) );
  MUX2X1 U8854 ( .B(ram[751]), .A(ram[687]), .S(n8545), .Y(n7817) );
  MUX2X1 U8855 ( .B(ram[879]), .A(ram[815]), .S(n8545), .Y(n7821) );
  MUX2X1 U8856 ( .B(ram[1007]), .A(ram[943]), .S(n8545), .Y(n7820) );
  MUX2X1 U8857 ( .B(n7819), .A(n7816), .S(n8407), .Y(n7823) );
  MUX2X1 U8858 ( .B(ram[1135]), .A(ram[1071]), .S(n8546), .Y(n7827) );
  MUX2X1 U8859 ( .B(ram[1263]), .A(ram[1199]), .S(n8546), .Y(n7826) );
  MUX2X1 U8860 ( .B(ram[1391]), .A(ram[1327]), .S(n8546), .Y(n7830) );
  MUX2X1 U8861 ( .B(ram[1519]), .A(ram[1455]), .S(n8546), .Y(n7829) );
  MUX2X1 U8862 ( .B(n7828), .A(n7825), .S(n8407), .Y(n7839) );
  MUX2X1 U8863 ( .B(ram[1647]), .A(ram[1583]), .S(n8546), .Y(n7833) );
  MUX2X1 U8864 ( .B(ram[1775]), .A(ram[1711]), .S(n8546), .Y(n7832) );
  MUX2X1 U8865 ( .B(ram[1903]), .A(ram[1839]), .S(n8546), .Y(n7836) );
  MUX2X1 U8866 ( .B(ram[2031]), .A(ram[1967]), .S(n8546), .Y(n7835) );
  MUX2X1 U8867 ( .B(n7834), .A(n7831), .S(n8407), .Y(n7838) );
  MUX2X1 U8868 ( .B(n7837), .A(n7822), .S(n8386), .Y(n8367) );
  MUX2X1 U8869 ( .B(ram[112]), .A(ram[48]), .S(n8546), .Y(n7842) );
  MUX2X1 U8870 ( .B(ram[240]), .A(ram[176]), .S(n8546), .Y(n7841) );
  MUX2X1 U8871 ( .B(ram[368]), .A(ram[304]), .S(n8546), .Y(n7845) );
  MUX2X1 U8872 ( .B(ram[496]), .A(ram[432]), .S(n8546), .Y(n7844) );
  MUX2X1 U8873 ( .B(n7843), .A(n7840), .S(n8407), .Y(n7854) );
  MUX2X1 U8874 ( .B(ram[624]), .A(ram[560]), .S(n8547), .Y(n7848) );
  MUX2X1 U8875 ( .B(ram[752]), .A(ram[688]), .S(n8547), .Y(n7847) );
  MUX2X1 U8876 ( .B(ram[880]), .A(ram[816]), .S(n8547), .Y(n7851) );
  MUX2X1 U8877 ( .B(ram[1008]), .A(ram[944]), .S(n8547), .Y(n7850) );
  MUX2X1 U8878 ( .B(n7849), .A(n7846), .S(n8407), .Y(n7853) );
  MUX2X1 U8879 ( .B(ram[1136]), .A(ram[1072]), .S(n8547), .Y(n7857) );
  MUX2X1 U8880 ( .B(ram[1264]), .A(ram[1200]), .S(n8547), .Y(n7856) );
  MUX2X1 U8881 ( .B(ram[1392]), .A(ram[1328]), .S(n8547), .Y(n7860) );
  MUX2X1 U8882 ( .B(ram[1520]), .A(ram[1456]), .S(n8547), .Y(n7859) );
  MUX2X1 U8883 ( .B(n7858), .A(n7855), .S(n8407), .Y(n7869) );
  MUX2X1 U8884 ( .B(ram[1648]), .A(ram[1584]), .S(n8547), .Y(n7863) );
  MUX2X1 U8885 ( .B(ram[1776]), .A(ram[1712]), .S(n8547), .Y(n7862) );
  MUX2X1 U8886 ( .B(ram[1904]), .A(ram[1840]), .S(n8547), .Y(n7866) );
  MUX2X1 U8887 ( .B(ram[2032]), .A(ram[1968]), .S(n8547), .Y(n7865) );
  MUX2X1 U8888 ( .B(n7864), .A(n7861), .S(n8407), .Y(n7868) );
  MUX2X1 U8889 ( .B(n7867), .A(n7852), .S(n8385), .Y(n8368) );
  MUX2X1 U8890 ( .B(ram[113]), .A(ram[49]), .S(n8548), .Y(n7872) );
  MUX2X1 U8891 ( .B(ram[241]), .A(ram[177]), .S(n8548), .Y(n7871) );
  MUX2X1 U8892 ( .B(ram[369]), .A(ram[305]), .S(n8548), .Y(n7875) );
  MUX2X1 U8893 ( .B(ram[497]), .A(ram[433]), .S(n8548), .Y(n7874) );
  MUX2X1 U8894 ( .B(n7873), .A(n7870), .S(n8404), .Y(n7884) );
  MUX2X1 U8895 ( .B(ram[625]), .A(ram[561]), .S(n8548), .Y(n7878) );
  MUX2X1 U8896 ( .B(ram[753]), .A(ram[689]), .S(n8548), .Y(n7877) );
  MUX2X1 U8897 ( .B(ram[881]), .A(ram[817]), .S(n8548), .Y(n7881) );
  MUX2X1 U8898 ( .B(ram[1009]), .A(ram[945]), .S(n8548), .Y(n7880) );
  MUX2X1 U8899 ( .B(n7879), .A(n7876), .S(n8410), .Y(n7883) );
  MUX2X1 U8900 ( .B(ram[1137]), .A(ram[1073]), .S(n8548), .Y(n7887) );
  MUX2X1 U8901 ( .B(ram[1265]), .A(ram[1201]), .S(n8548), .Y(n7886) );
  MUX2X1 U8902 ( .B(ram[1393]), .A(ram[1329]), .S(n8548), .Y(n7890) );
  MUX2X1 U8903 ( .B(ram[1521]), .A(ram[1457]), .S(n8548), .Y(n7889) );
  MUX2X1 U8904 ( .B(n7888), .A(n7885), .S(n8404), .Y(n7899) );
  MUX2X1 U8905 ( .B(ram[1649]), .A(ram[1585]), .S(n8549), .Y(n7893) );
  MUX2X1 U8906 ( .B(ram[1777]), .A(ram[1713]), .S(n8549), .Y(n7892) );
  MUX2X1 U8907 ( .B(ram[1905]), .A(ram[1841]), .S(n8549), .Y(n7896) );
  MUX2X1 U8908 ( .B(ram[2033]), .A(ram[1969]), .S(n8549), .Y(n7895) );
  MUX2X1 U8909 ( .B(n7894), .A(n7891), .S(n8399), .Y(n7898) );
  MUX2X1 U8910 ( .B(n7897), .A(n7882), .S(n8385), .Y(n8369) );
  MUX2X1 U8911 ( .B(ram[114]), .A(ram[50]), .S(n8549), .Y(n7902) );
  MUX2X1 U8912 ( .B(ram[242]), .A(ram[178]), .S(n8549), .Y(n7901) );
  MUX2X1 U8913 ( .B(ram[370]), .A(ram[306]), .S(n8549), .Y(n7905) );
  MUX2X1 U8914 ( .B(ram[498]), .A(ram[434]), .S(n8549), .Y(n7904) );
  MUX2X1 U8915 ( .B(n7903), .A(n7900), .S(n8402), .Y(n7914) );
  MUX2X1 U8916 ( .B(ram[626]), .A(ram[562]), .S(n8549), .Y(n7908) );
  MUX2X1 U8917 ( .B(ram[754]), .A(ram[690]), .S(n8549), .Y(n7907) );
  MUX2X1 U8918 ( .B(ram[882]), .A(ram[818]), .S(n8549), .Y(n7911) );
  MUX2X1 U8919 ( .B(ram[1010]), .A(ram[946]), .S(n8549), .Y(n7910) );
  MUX2X1 U8920 ( .B(n7909), .A(n7906), .S(n8403), .Y(n7913) );
  MUX2X1 U8921 ( .B(ram[1138]), .A(ram[1074]), .S(n8550), .Y(n7917) );
  MUX2X1 U8922 ( .B(ram[1266]), .A(ram[1202]), .S(n8550), .Y(n7916) );
  MUX2X1 U8923 ( .B(ram[1394]), .A(ram[1330]), .S(n8550), .Y(n7920) );
  MUX2X1 U8924 ( .B(ram[1522]), .A(ram[1458]), .S(n8550), .Y(n7919) );
  MUX2X1 U8925 ( .B(n7918), .A(n7915), .S(n8405), .Y(n7929) );
  MUX2X1 U8926 ( .B(ram[1650]), .A(ram[1586]), .S(n8550), .Y(n7923) );
  MUX2X1 U8927 ( .B(ram[1778]), .A(ram[1714]), .S(n8550), .Y(n7922) );
  MUX2X1 U8928 ( .B(ram[1906]), .A(ram[1842]), .S(n8550), .Y(n7926) );
  MUX2X1 U8929 ( .B(ram[2034]), .A(ram[1970]), .S(n8550), .Y(n7925) );
  MUX2X1 U8930 ( .B(n7924), .A(n7921), .S(n8398), .Y(n7928) );
  MUX2X1 U8931 ( .B(n7927), .A(n7912), .S(n8385), .Y(n8370) );
  MUX2X1 U8932 ( .B(ram[115]), .A(ram[51]), .S(n8550), .Y(n7932) );
  MUX2X1 U8933 ( .B(ram[243]), .A(ram[179]), .S(n8550), .Y(n7931) );
  MUX2X1 U8934 ( .B(ram[371]), .A(ram[307]), .S(n8550), .Y(n7935) );
  MUX2X1 U8935 ( .B(ram[499]), .A(ram[435]), .S(n8550), .Y(n7934) );
  MUX2X1 U8936 ( .B(n7933), .A(n7930), .S(n8407), .Y(n7944) );
  MUX2X1 U8937 ( .B(ram[627]), .A(ram[563]), .S(n8551), .Y(n7938) );
  MUX2X1 U8938 ( .B(ram[755]), .A(ram[691]), .S(n8551), .Y(n7937) );
  MUX2X1 U8939 ( .B(ram[883]), .A(ram[819]), .S(n8551), .Y(n7941) );
  MUX2X1 U8940 ( .B(ram[1011]), .A(ram[947]), .S(n8551), .Y(n7940) );
  MUX2X1 U8941 ( .B(n7939), .A(n7936), .S(n8401), .Y(n7943) );
  MUX2X1 U8942 ( .B(ram[1139]), .A(ram[1075]), .S(n8551), .Y(n7947) );
  MUX2X1 U8943 ( .B(ram[1267]), .A(ram[1203]), .S(n8551), .Y(n7946) );
  MUX2X1 U8944 ( .B(ram[1395]), .A(ram[1331]), .S(n8551), .Y(n7950) );
  MUX2X1 U8945 ( .B(ram[1523]), .A(ram[1459]), .S(n8551), .Y(n7949) );
  MUX2X1 U8946 ( .B(n7948), .A(n7945), .S(n8409), .Y(n7959) );
  MUX2X1 U8947 ( .B(ram[1651]), .A(ram[1587]), .S(n8551), .Y(n7953) );
  MUX2X1 U8948 ( .B(ram[1779]), .A(ram[1715]), .S(n8551), .Y(n7952) );
  MUX2X1 U8949 ( .B(ram[1907]), .A(ram[1843]), .S(n8551), .Y(n7956) );
  MUX2X1 U8950 ( .B(ram[2035]), .A(ram[1971]), .S(n8551), .Y(n7955) );
  MUX2X1 U8951 ( .B(n7954), .A(n7951), .S(n8408), .Y(n7958) );
  MUX2X1 U8952 ( .B(n7957), .A(n7942), .S(n8385), .Y(n8371) );
  MUX2X1 U8953 ( .B(ram[116]), .A(ram[52]), .S(n8552), .Y(n7962) );
  MUX2X1 U8954 ( .B(ram[244]), .A(ram[180]), .S(n8552), .Y(n7961) );
  MUX2X1 U8955 ( .B(ram[372]), .A(ram[308]), .S(n8552), .Y(n7965) );
  MUX2X1 U8956 ( .B(ram[500]), .A(ram[436]), .S(n8552), .Y(n7964) );
  MUX2X1 U8957 ( .B(n7963), .A(n7960), .S(n8408), .Y(n7974) );
  MUX2X1 U8958 ( .B(ram[628]), .A(ram[564]), .S(n8552), .Y(n7968) );
  MUX2X1 U8959 ( .B(ram[756]), .A(ram[692]), .S(n8552), .Y(n7967) );
  MUX2X1 U8960 ( .B(ram[884]), .A(ram[820]), .S(n8552), .Y(n7971) );
  MUX2X1 U8961 ( .B(ram[1012]), .A(ram[948]), .S(n8552), .Y(n7970) );
  MUX2X1 U8962 ( .B(n7969), .A(n7966), .S(n8408), .Y(n7973) );
  MUX2X1 U8963 ( .B(ram[1140]), .A(ram[1076]), .S(n8552), .Y(n7977) );
  MUX2X1 U8964 ( .B(ram[1268]), .A(ram[1204]), .S(n8552), .Y(n7976) );
  MUX2X1 U8965 ( .B(ram[1396]), .A(ram[1332]), .S(n8552), .Y(n7980) );
  MUX2X1 U8966 ( .B(ram[1524]), .A(ram[1460]), .S(n8552), .Y(n7979) );
  MUX2X1 U8967 ( .B(n7978), .A(n7975), .S(n8408), .Y(n7989) );
  MUX2X1 U8968 ( .B(ram[1652]), .A(ram[1588]), .S(n8553), .Y(n7983) );
  MUX2X1 U8969 ( .B(ram[1780]), .A(ram[1716]), .S(n8553), .Y(n7982) );
  MUX2X1 U8970 ( .B(ram[1908]), .A(ram[1844]), .S(n8553), .Y(n7986) );
  MUX2X1 U8971 ( .B(ram[2036]), .A(ram[1972]), .S(n8553), .Y(n7985) );
  MUX2X1 U8972 ( .B(n7984), .A(n7981), .S(n8408), .Y(n7988) );
  MUX2X1 U8973 ( .B(n7987), .A(n7972), .S(n8385), .Y(n8372) );
  MUX2X1 U8974 ( .B(ram[117]), .A(ram[53]), .S(n8553), .Y(n7992) );
  MUX2X1 U8975 ( .B(ram[245]), .A(ram[181]), .S(n8553), .Y(n7991) );
  MUX2X1 U8976 ( .B(ram[373]), .A(ram[309]), .S(n8553), .Y(n7995) );
  MUX2X1 U8977 ( .B(ram[501]), .A(ram[437]), .S(n8553), .Y(n7994) );
  MUX2X1 U8978 ( .B(n7993), .A(n7990), .S(n8408), .Y(n8004) );
  MUX2X1 U8979 ( .B(ram[629]), .A(ram[565]), .S(n8553), .Y(n7998) );
  MUX2X1 U8980 ( .B(ram[757]), .A(ram[693]), .S(n8553), .Y(n7997) );
  MUX2X1 U8981 ( .B(ram[885]), .A(ram[821]), .S(n8553), .Y(n8001) );
  MUX2X1 U8982 ( .B(ram[1013]), .A(ram[949]), .S(n8553), .Y(n8000) );
  MUX2X1 U8983 ( .B(n7999), .A(n7996), .S(n8408), .Y(n8003) );
  MUX2X1 U8984 ( .B(ram[1141]), .A(ram[1077]), .S(n8554), .Y(n8007) );
  MUX2X1 U8985 ( .B(ram[1269]), .A(ram[1205]), .S(n8554), .Y(n8006) );
  MUX2X1 U8986 ( .B(ram[1397]), .A(ram[1333]), .S(n8554), .Y(n8010) );
  MUX2X1 U8987 ( .B(ram[1525]), .A(ram[1461]), .S(n8554), .Y(n8009) );
  MUX2X1 U8988 ( .B(n8008), .A(n8005), .S(n8408), .Y(n8019) );
  MUX2X1 U8989 ( .B(ram[1653]), .A(ram[1589]), .S(n8554), .Y(n8013) );
  MUX2X1 U8990 ( .B(ram[1781]), .A(ram[1717]), .S(n8554), .Y(n8012) );
  MUX2X1 U8991 ( .B(ram[1909]), .A(ram[1845]), .S(n8554), .Y(n8016) );
  MUX2X1 U8992 ( .B(ram[2037]), .A(ram[1973]), .S(n8554), .Y(n8015) );
  MUX2X1 U8993 ( .B(n8014), .A(n8011), .S(n8408), .Y(n8018) );
  MUX2X1 U8994 ( .B(n8017), .A(n8002), .S(n8385), .Y(n8373) );
  MUX2X1 U8995 ( .B(ram[118]), .A(ram[54]), .S(n8554), .Y(n8022) );
  MUX2X1 U8996 ( .B(ram[246]), .A(ram[182]), .S(n8554), .Y(n8021) );
  MUX2X1 U8997 ( .B(ram[374]), .A(ram[310]), .S(n8554), .Y(n8025) );
  MUX2X1 U8998 ( .B(ram[502]), .A(ram[438]), .S(n8554), .Y(n8024) );
  MUX2X1 U8999 ( .B(n8023), .A(n8020), .S(n8408), .Y(n8034) );
  MUX2X1 U9000 ( .B(ram[630]), .A(ram[566]), .S(n8555), .Y(n8028) );
  MUX2X1 U9001 ( .B(ram[758]), .A(ram[694]), .S(n8555), .Y(n8027) );
  MUX2X1 U9002 ( .B(ram[886]), .A(ram[822]), .S(n8555), .Y(n8031) );
  MUX2X1 U9003 ( .B(ram[1014]), .A(ram[950]), .S(n8555), .Y(n8030) );
  MUX2X1 U9004 ( .B(n8029), .A(n8026), .S(n8408), .Y(n8033) );
  MUX2X1 U9005 ( .B(ram[1142]), .A(ram[1078]), .S(n8555), .Y(n8037) );
  MUX2X1 U9006 ( .B(ram[1270]), .A(ram[1206]), .S(n8555), .Y(n8036) );
  MUX2X1 U9007 ( .B(ram[1398]), .A(ram[1334]), .S(n8555), .Y(n8040) );
  MUX2X1 U9008 ( .B(ram[1526]), .A(ram[1462]), .S(n8555), .Y(n8039) );
  MUX2X1 U9009 ( .B(n8038), .A(n8035), .S(n8408), .Y(n8049) );
  MUX2X1 U9010 ( .B(ram[1654]), .A(ram[1590]), .S(n8555), .Y(n8043) );
  MUX2X1 U9011 ( .B(ram[1782]), .A(ram[1718]), .S(n8555), .Y(n8042) );
  MUX2X1 U9012 ( .B(ram[1910]), .A(ram[1846]), .S(n8555), .Y(n8046) );
  MUX2X1 U9013 ( .B(ram[2038]), .A(ram[1974]), .S(n8555), .Y(n8045) );
  MUX2X1 U9014 ( .B(n8044), .A(n8041), .S(n8408), .Y(n8048) );
  MUX2X1 U9015 ( .B(n8047), .A(n8032), .S(n8385), .Y(n8374) );
  MUX2X1 U9016 ( .B(ram[119]), .A(ram[55]), .S(n8556), .Y(n8052) );
  MUX2X1 U9017 ( .B(ram[247]), .A(ram[183]), .S(n8556), .Y(n8051) );
  MUX2X1 U9018 ( .B(ram[375]), .A(ram[311]), .S(n8556), .Y(n8055) );
  MUX2X1 U9019 ( .B(ram[503]), .A(ram[439]), .S(n8556), .Y(n8054) );
  MUX2X1 U9020 ( .B(n8053), .A(n8050), .S(n8409), .Y(n8064) );
  MUX2X1 U9021 ( .B(ram[631]), .A(ram[567]), .S(n8556), .Y(n8058) );
  MUX2X1 U9022 ( .B(ram[759]), .A(ram[695]), .S(n8556), .Y(n8057) );
  MUX2X1 U9023 ( .B(ram[887]), .A(ram[823]), .S(n8556), .Y(n8061) );
  MUX2X1 U9024 ( .B(ram[1015]), .A(ram[951]), .S(n8556), .Y(n8060) );
  MUX2X1 U9025 ( .B(n8059), .A(n8056), .S(n8409), .Y(n8063) );
  MUX2X1 U9026 ( .B(ram[1143]), .A(ram[1079]), .S(n8556), .Y(n8067) );
  MUX2X1 U9027 ( .B(ram[1271]), .A(ram[1207]), .S(n8556), .Y(n8066) );
  MUX2X1 U9028 ( .B(ram[1399]), .A(ram[1335]), .S(n8556), .Y(n8070) );
  MUX2X1 U9029 ( .B(ram[1527]), .A(ram[1463]), .S(n8556), .Y(n8069) );
  MUX2X1 U9030 ( .B(n8068), .A(n8065), .S(n8409), .Y(n8079) );
  MUX2X1 U9031 ( .B(ram[1655]), .A(ram[1591]), .S(n8557), .Y(n8073) );
  MUX2X1 U9032 ( .B(ram[1783]), .A(ram[1719]), .S(n8557), .Y(n8072) );
  MUX2X1 U9033 ( .B(ram[1911]), .A(ram[1847]), .S(n8557), .Y(n8076) );
  MUX2X1 U9034 ( .B(ram[2039]), .A(ram[1975]), .S(n8557), .Y(n8075) );
  MUX2X1 U9035 ( .B(n8074), .A(n8071), .S(n8409), .Y(n8078) );
  MUX2X1 U9036 ( .B(n8077), .A(n8062), .S(n8385), .Y(n8375) );
  MUX2X1 U9037 ( .B(ram[120]), .A(ram[56]), .S(n8557), .Y(n8082) );
  MUX2X1 U9038 ( .B(ram[248]), .A(ram[184]), .S(n8557), .Y(n8081) );
  MUX2X1 U9039 ( .B(ram[376]), .A(ram[312]), .S(n8557), .Y(n8085) );
  MUX2X1 U9040 ( .B(ram[504]), .A(ram[440]), .S(n8557), .Y(n8084) );
  MUX2X1 U9041 ( .B(n8083), .A(n8080), .S(n8409), .Y(n8094) );
  MUX2X1 U9042 ( .B(ram[632]), .A(ram[568]), .S(n8557), .Y(n8088) );
  MUX2X1 U9043 ( .B(ram[760]), .A(ram[696]), .S(n8557), .Y(n8087) );
  MUX2X1 U9044 ( .B(ram[888]), .A(ram[824]), .S(n8557), .Y(n8091) );
  MUX2X1 U9045 ( .B(ram[1016]), .A(ram[952]), .S(n8557), .Y(n8090) );
  MUX2X1 U9046 ( .B(n8089), .A(n8086), .S(n8409), .Y(n8093) );
  MUX2X1 U9047 ( .B(ram[1144]), .A(ram[1080]), .S(n8558), .Y(n8097) );
  MUX2X1 U9048 ( .B(ram[1272]), .A(ram[1208]), .S(n8558), .Y(n8096) );
  MUX2X1 U9049 ( .B(ram[1400]), .A(ram[1336]), .S(n8558), .Y(n8100) );
  MUX2X1 U9050 ( .B(ram[1528]), .A(ram[1464]), .S(n8558), .Y(n8099) );
  MUX2X1 U9051 ( .B(n8098), .A(n8095), .S(n8409), .Y(n8109) );
  MUX2X1 U9052 ( .B(ram[1656]), .A(ram[1592]), .S(n8558), .Y(n8103) );
  MUX2X1 U9053 ( .B(ram[1784]), .A(ram[1720]), .S(n8558), .Y(n8102) );
  MUX2X1 U9054 ( .B(ram[1912]), .A(ram[1848]), .S(n8558), .Y(n8106) );
  MUX2X1 U9055 ( .B(ram[2040]), .A(ram[1976]), .S(n8558), .Y(n8105) );
  MUX2X1 U9056 ( .B(n8104), .A(n8101), .S(n8409), .Y(n8108) );
  MUX2X1 U9057 ( .B(n8107), .A(n8092), .S(n8385), .Y(n8376) );
  MUX2X1 U9058 ( .B(ram[121]), .A(ram[57]), .S(n8558), .Y(n8112) );
  MUX2X1 U9059 ( .B(ram[249]), .A(ram[185]), .S(n8558), .Y(n8111) );
  MUX2X1 U9060 ( .B(ram[377]), .A(ram[313]), .S(n8558), .Y(n8115) );
  MUX2X1 U9061 ( .B(ram[505]), .A(ram[441]), .S(n8558), .Y(n8114) );
  MUX2X1 U9062 ( .B(n8113), .A(n8110), .S(n8409), .Y(n8124) );
  MUX2X1 U9063 ( .B(ram[633]), .A(ram[569]), .S(n8559), .Y(n8118) );
  MUX2X1 U9064 ( .B(ram[761]), .A(ram[697]), .S(n8559), .Y(n8117) );
  MUX2X1 U9065 ( .B(ram[889]), .A(ram[825]), .S(n8559), .Y(n8121) );
  MUX2X1 U9066 ( .B(ram[1017]), .A(ram[953]), .S(n8559), .Y(n8120) );
  MUX2X1 U9067 ( .B(n8119), .A(n8116), .S(n8409), .Y(n8123) );
  MUX2X1 U9068 ( .B(ram[1145]), .A(ram[1081]), .S(n8559), .Y(n8127) );
  MUX2X1 U9069 ( .B(ram[1273]), .A(ram[1209]), .S(n8559), .Y(n8126) );
  MUX2X1 U9070 ( .B(ram[1401]), .A(ram[1337]), .S(n8559), .Y(n8130) );
  MUX2X1 U9071 ( .B(ram[1529]), .A(ram[1465]), .S(n8559), .Y(n8129) );
  MUX2X1 U9072 ( .B(n8128), .A(n8125), .S(n8409), .Y(n8139) );
  MUX2X1 U9073 ( .B(ram[1657]), .A(ram[1593]), .S(n8559), .Y(n8133) );
  MUX2X1 U9074 ( .B(ram[1785]), .A(ram[1721]), .S(n8559), .Y(n8132) );
  MUX2X1 U9075 ( .B(ram[1913]), .A(ram[1849]), .S(n8559), .Y(n8136) );
  MUX2X1 U9076 ( .B(ram[2041]), .A(ram[1977]), .S(n8559), .Y(n8135) );
  MUX2X1 U9077 ( .B(n8134), .A(n8131), .S(n8409), .Y(n8138) );
  MUX2X1 U9078 ( .B(n8137), .A(n8122), .S(n8385), .Y(n8377) );
  MUX2X1 U9079 ( .B(ram[122]), .A(ram[58]), .S(n8560), .Y(n8142) );
  MUX2X1 U9080 ( .B(ram[250]), .A(ram[186]), .S(n8560), .Y(n8141) );
  MUX2X1 U9081 ( .B(ram[378]), .A(ram[314]), .S(n8560), .Y(n8145) );
  MUX2X1 U9082 ( .B(ram[506]), .A(ram[442]), .S(n8560), .Y(n8144) );
  MUX2X1 U9083 ( .B(n8143), .A(n8140), .S(n8410), .Y(n8154) );
  MUX2X1 U9084 ( .B(ram[634]), .A(ram[570]), .S(n8560), .Y(n8148) );
  MUX2X1 U9085 ( .B(ram[762]), .A(ram[698]), .S(n8560), .Y(n8147) );
  MUX2X1 U9086 ( .B(ram[890]), .A(ram[826]), .S(n8560), .Y(n8151) );
  MUX2X1 U9087 ( .B(ram[1018]), .A(ram[954]), .S(n8560), .Y(n8150) );
  MUX2X1 U9088 ( .B(n8149), .A(n8146), .S(n8410), .Y(n8153) );
  MUX2X1 U9089 ( .B(ram[1146]), .A(ram[1082]), .S(n8560), .Y(n8157) );
  MUX2X1 U9090 ( .B(ram[1274]), .A(ram[1210]), .S(n8560), .Y(n8156) );
  MUX2X1 U9091 ( .B(ram[1402]), .A(ram[1338]), .S(n8560), .Y(n8160) );
  MUX2X1 U9092 ( .B(ram[1530]), .A(ram[1466]), .S(n8560), .Y(n8159) );
  MUX2X1 U9093 ( .B(n8158), .A(n8155), .S(n8410), .Y(n8169) );
  MUX2X1 U9094 ( .B(ram[1658]), .A(ram[1594]), .S(n8561), .Y(n8163) );
  MUX2X1 U9095 ( .B(ram[1786]), .A(ram[1722]), .S(n8561), .Y(n8162) );
  MUX2X1 U9096 ( .B(ram[1914]), .A(ram[1850]), .S(n8561), .Y(n8166) );
  MUX2X1 U9097 ( .B(ram[2042]), .A(ram[1978]), .S(n8561), .Y(n8165) );
  MUX2X1 U9098 ( .B(n8164), .A(n8161), .S(n8410), .Y(n8168) );
  MUX2X1 U9099 ( .B(n8167), .A(n8152), .S(n8385), .Y(n8378) );
  MUX2X1 U9100 ( .B(ram[123]), .A(ram[59]), .S(n8561), .Y(n8172) );
  MUX2X1 U9101 ( .B(ram[251]), .A(ram[187]), .S(n8561), .Y(n8171) );
  MUX2X1 U9102 ( .B(ram[379]), .A(ram[315]), .S(n8561), .Y(n8175) );
  MUX2X1 U9103 ( .B(ram[507]), .A(ram[443]), .S(n8561), .Y(n8174) );
  MUX2X1 U9104 ( .B(n8173), .A(n8170), .S(n8410), .Y(n8184) );
  MUX2X1 U9105 ( .B(ram[635]), .A(ram[571]), .S(n8561), .Y(n8178) );
  MUX2X1 U9106 ( .B(ram[763]), .A(ram[699]), .S(n8561), .Y(n8177) );
  MUX2X1 U9107 ( .B(ram[891]), .A(ram[827]), .S(n8561), .Y(n8181) );
  MUX2X1 U9108 ( .B(ram[1019]), .A(ram[955]), .S(n8561), .Y(n8180) );
  MUX2X1 U9109 ( .B(n8179), .A(n8176), .S(n8410), .Y(n8183) );
  MUX2X1 U9110 ( .B(ram[1147]), .A(ram[1083]), .S(n8562), .Y(n8187) );
  MUX2X1 U9111 ( .B(ram[1275]), .A(ram[1211]), .S(n8562), .Y(n8186) );
  MUX2X1 U9112 ( .B(ram[1403]), .A(ram[1339]), .S(n8562), .Y(n8190) );
  MUX2X1 U9113 ( .B(ram[1531]), .A(ram[1467]), .S(n8562), .Y(n8189) );
  MUX2X1 U9114 ( .B(n8188), .A(n8185), .S(n8410), .Y(n8199) );
  MUX2X1 U9115 ( .B(ram[1659]), .A(ram[1595]), .S(n8562), .Y(n8193) );
  MUX2X1 U9116 ( .B(ram[1787]), .A(ram[1723]), .S(n8562), .Y(n8192) );
  MUX2X1 U9117 ( .B(ram[1915]), .A(ram[1851]), .S(n8562), .Y(n8196) );
  MUX2X1 U9118 ( .B(ram[2043]), .A(ram[1979]), .S(n8562), .Y(n8195) );
  MUX2X1 U9119 ( .B(n8194), .A(n8191), .S(n8410), .Y(n8198) );
  MUX2X1 U9120 ( .B(n8197), .A(n8182), .S(n8385), .Y(n8379) );
  MUX2X1 U9121 ( .B(ram[124]), .A(ram[60]), .S(n8562), .Y(n8202) );
  MUX2X1 U9122 ( .B(ram[252]), .A(ram[188]), .S(n8562), .Y(n8201) );
  MUX2X1 U9123 ( .B(ram[380]), .A(ram[316]), .S(n8562), .Y(n8205) );
  MUX2X1 U9124 ( .B(ram[508]), .A(ram[444]), .S(n8562), .Y(n8204) );
  MUX2X1 U9125 ( .B(n8203), .A(n8200), .S(n8410), .Y(n8214) );
  MUX2X1 U9126 ( .B(ram[636]), .A(ram[572]), .S(n8563), .Y(n8208) );
  MUX2X1 U9127 ( .B(ram[764]), .A(ram[700]), .S(n8563), .Y(n8207) );
  MUX2X1 U9128 ( .B(ram[892]), .A(ram[828]), .S(n8563), .Y(n8211) );
  MUX2X1 U9129 ( .B(ram[1020]), .A(ram[956]), .S(n8563), .Y(n8210) );
  MUX2X1 U9130 ( .B(n8209), .A(n8206), .S(n8410), .Y(n8213) );
  MUX2X1 U9131 ( .B(ram[1148]), .A(ram[1084]), .S(n8563), .Y(n8217) );
  MUX2X1 U9132 ( .B(ram[1276]), .A(ram[1212]), .S(n8563), .Y(n8216) );
  MUX2X1 U9133 ( .B(ram[1404]), .A(ram[1340]), .S(n8563), .Y(n8220) );
  MUX2X1 U9134 ( .B(ram[1532]), .A(ram[1468]), .S(n8563), .Y(n8219) );
  MUX2X1 U9135 ( .B(n8218), .A(n8215), .S(n8410), .Y(n8229) );
  MUX2X1 U9136 ( .B(ram[1660]), .A(ram[1596]), .S(n8563), .Y(n8223) );
  MUX2X1 U9137 ( .B(ram[1788]), .A(ram[1724]), .S(n8563), .Y(n8222) );
  MUX2X1 U9138 ( .B(ram[1916]), .A(ram[1852]), .S(n8563), .Y(n8226) );
  MUX2X1 U9139 ( .B(ram[2044]), .A(ram[1980]), .S(n8563), .Y(n8225) );
  MUX2X1 U9140 ( .B(n8224), .A(n8221), .S(n8410), .Y(n8228) );
  MUX2X1 U9141 ( .B(n8227), .A(n8212), .S(n8386), .Y(n8380) );
  MUX2X1 U9142 ( .B(ram[125]), .A(ram[61]), .S(n8564), .Y(n8232) );
  MUX2X1 U9143 ( .B(ram[253]), .A(ram[189]), .S(n8564), .Y(n8231) );
  MUX2X1 U9144 ( .B(ram[381]), .A(ram[317]), .S(n8564), .Y(n8235) );
  MUX2X1 U9145 ( .B(ram[509]), .A(ram[445]), .S(n8564), .Y(n8234) );
  MUX2X1 U9146 ( .B(n8233), .A(n8230), .S(n8405), .Y(n8244) );
  MUX2X1 U9147 ( .B(ram[637]), .A(ram[573]), .S(n8564), .Y(n8238) );
  MUX2X1 U9148 ( .B(ram[765]), .A(ram[701]), .S(n8564), .Y(n8237) );
  MUX2X1 U9149 ( .B(ram[893]), .A(ram[829]), .S(n8564), .Y(n8241) );
  MUX2X1 U9150 ( .B(ram[1021]), .A(ram[957]), .S(n8564), .Y(n8240) );
  MUX2X1 U9151 ( .B(n8239), .A(n8236), .S(n8406), .Y(n8243) );
  MUX2X1 U9152 ( .B(ram[1149]), .A(ram[1085]), .S(n8564), .Y(n8247) );
  MUX2X1 U9153 ( .B(ram[1277]), .A(ram[1213]), .S(n8564), .Y(n8246) );
  MUX2X1 U9154 ( .B(ram[1405]), .A(ram[1341]), .S(n8564), .Y(n8250) );
  MUX2X1 U9155 ( .B(ram[1533]), .A(ram[1469]), .S(n8564), .Y(n8249) );
  MUX2X1 U9156 ( .B(n8248), .A(n8245), .S(n8407), .Y(n8259) );
  MUX2X1 U9157 ( .B(ram[1661]), .A(ram[1597]), .S(n8565), .Y(n8253) );
  MUX2X1 U9158 ( .B(ram[1789]), .A(ram[1725]), .S(n8565), .Y(n8252) );
  MUX2X1 U9159 ( .B(ram[1917]), .A(ram[1853]), .S(n8565), .Y(n8256) );
  MUX2X1 U9160 ( .B(ram[2045]), .A(ram[1981]), .S(n8565), .Y(n8255) );
  MUX2X1 U9161 ( .B(n8254), .A(n8251), .S(n8408), .Y(n8258) );
  MUX2X1 U9162 ( .B(n8257), .A(n8242), .S(n8386), .Y(n8381) );
  MUX2X1 U9163 ( .B(ram[126]), .A(ram[62]), .S(n8565), .Y(n8262) );
  MUX2X1 U9164 ( .B(ram[254]), .A(ram[190]), .S(n8565), .Y(n8261) );
  MUX2X1 U9165 ( .B(ram[382]), .A(ram[318]), .S(n8565), .Y(n8265) );
  MUX2X1 U9166 ( .B(ram[510]), .A(ram[446]), .S(n8565), .Y(n8264) );
  MUX2X1 U9167 ( .B(n8263), .A(n8260), .S(n8408), .Y(n8274) );
  MUX2X1 U9168 ( .B(ram[638]), .A(ram[574]), .S(n8565), .Y(n8268) );
  MUX2X1 U9169 ( .B(ram[766]), .A(ram[702]), .S(n8565), .Y(n8267) );
  MUX2X1 U9170 ( .B(ram[894]), .A(ram[830]), .S(n8565), .Y(n8271) );
  MUX2X1 U9171 ( .B(ram[1022]), .A(ram[958]), .S(n8565), .Y(n8270) );
  MUX2X1 U9172 ( .B(n8269), .A(n8266), .S(n8402), .Y(n8273) );
  MUX2X1 U9173 ( .B(ram[1150]), .A(ram[1086]), .S(n8566), .Y(n8277) );
  MUX2X1 U9174 ( .B(ram[1278]), .A(ram[1214]), .S(n8566), .Y(n8276) );
  MUX2X1 U9175 ( .B(ram[1406]), .A(ram[1342]), .S(n8566), .Y(n8280) );
  MUX2X1 U9176 ( .B(ram[1534]), .A(ram[1470]), .S(n8566), .Y(n8279) );
  MUX2X1 U9177 ( .B(n8278), .A(n8275), .S(n8410), .Y(n8289) );
  MUX2X1 U9178 ( .B(ram[1662]), .A(ram[1598]), .S(n8566), .Y(n8283) );
  MUX2X1 U9179 ( .B(ram[1790]), .A(ram[1726]), .S(n8566), .Y(n8282) );
  MUX2X1 U9180 ( .B(ram[1918]), .A(ram[1854]), .S(n8566), .Y(n8286) );
  MUX2X1 U9181 ( .B(ram[2046]), .A(ram[1982]), .S(n8566), .Y(n8285) );
  MUX2X1 U9182 ( .B(n8284), .A(n8281), .S(n8409), .Y(n8288) );
  MUX2X1 U9183 ( .B(n8287), .A(n8272), .S(n8385), .Y(n8382) );
  MUX2X1 U9184 ( .B(ram[127]), .A(ram[63]), .S(n8566), .Y(n8292) );
  MUX2X1 U9185 ( .B(ram[255]), .A(ram[191]), .S(n8566), .Y(n8291) );
  MUX2X1 U9186 ( .B(ram[383]), .A(ram[319]), .S(n8566), .Y(n8295) );
  MUX2X1 U9187 ( .B(ram[511]), .A(ram[447]), .S(n8566), .Y(n8294) );
  MUX2X1 U9188 ( .B(n8293), .A(n8290), .S(n8404), .Y(n8304) );
  MUX2X1 U9189 ( .B(ram[639]), .A(ram[575]), .S(n8567), .Y(n8298) );
  MUX2X1 U9190 ( .B(ram[767]), .A(ram[703]), .S(n8567), .Y(n8297) );
  MUX2X1 U9191 ( .B(ram[895]), .A(ram[831]), .S(n8567), .Y(n8301) );
  MUX2X1 U9192 ( .B(ram[1023]), .A(ram[959]), .S(n8567), .Y(n8300) );
  MUX2X1 U9193 ( .B(n8299), .A(n8296), .S(n8405), .Y(n8303) );
  MUX2X1 U9194 ( .B(ram[1151]), .A(ram[1087]), .S(n8567), .Y(n8307) );
  MUX2X1 U9195 ( .B(ram[1279]), .A(ram[1215]), .S(n8567), .Y(n8306) );
  MUX2X1 U9196 ( .B(ram[1407]), .A(ram[1343]), .S(n8567), .Y(n8310) );
  MUX2X1 U9197 ( .B(ram[1535]), .A(ram[1471]), .S(n8567), .Y(n8309) );
  MUX2X1 U9198 ( .B(n8308), .A(n8305), .S(n8401), .Y(n8319) );
  MUX2X1 U9199 ( .B(ram[1663]), .A(ram[1599]), .S(n8567), .Y(n8313) );
  MUX2X1 U9200 ( .B(ram[1791]), .A(ram[1727]), .S(n8567), .Y(n8312) );
  MUX2X1 U9201 ( .B(ram[1919]), .A(ram[1855]), .S(n8567), .Y(n8316) );
  MUX2X1 U9202 ( .B(ram[2047]), .A(ram[1983]), .S(n8567), .Y(n8315) );
  MUX2X1 U9203 ( .B(n8314), .A(n8311), .S(n8398), .Y(n8318) );
  MUX2X1 U9204 ( .B(n8317), .A(n8302), .S(n8386), .Y(n8383) );
  MUX2X1 U9205 ( .B(n8577), .A(n8578), .S(n10590), .Y(n8576) );
  MUX2X1 U9206 ( .B(n8580), .A(n8581), .S(n10590), .Y(n8579) );
  MUX2X1 U9207 ( .B(n8583), .A(n8584), .S(n10590), .Y(n8582) );
  MUX2X1 U9208 ( .B(n8586), .A(n8587), .S(n10590), .Y(n8585) );
  MUX2X1 U9209 ( .B(n8589), .A(n8590), .S(n10564), .Y(n8588) );
  MUX2X1 U9210 ( .B(n8592), .A(n8593), .S(n10590), .Y(n8591) );
  MUX2X1 U9211 ( .B(n8595), .A(n8596), .S(n10590), .Y(n8594) );
  MUX2X1 U9212 ( .B(n8598), .A(n8599), .S(n10590), .Y(n8597) );
  MUX2X1 U9213 ( .B(n8601), .A(n8602), .S(n10590), .Y(n8600) );
  MUX2X1 U9214 ( .B(n8604), .A(n8605), .S(read2_addr[1]), .Y(n8603) );
  MUX2X1 U9215 ( .B(n8607), .A(n8608), .S(n10591), .Y(n8606) );
  MUX2X1 U9216 ( .B(n8610), .A(n8611), .S(n10591), .Y(n8609) );
  MUX2X1 U9217 ( .B(n8613), .A(n8614), .S(n10591), .Y(n8612) );
  MUX2X1 U9218 ( .B(n8616), .A(n8617), .S(n10591), .Y(n8615) );
  MUX2X1 U9219 ( .B(n8619), .A(n8620), .S(n10563), .Y(n8618) );
  MUX2X1 U9220 ( .B(n8622), .A(n8623), .S(n10591), .Y(n8621) );
  MUX2X1 U9221 ( .B(n8625), .A(n8626), .S(n10591), .Y(n8624) );
  MUX2X1 U9222 ( .B(n8628), .A(n8629), .S(n10591), .Y(n8627) );
  MUX2X1 U9223 ( .B(n8631), .A(n8632), .S(n10591), .Y(n8630) );
  MUX2X1 U9224 ( .B(n8634), .A(n8635), .S(n10565), .Y(n8633) );
  MUX2X1 U9225 ( .B(n8637), .A(n8638), .S(n10591), .Y(n8636) );
  MUX2X1 U9226 ( .B(n8640), .A(n8641), .S(n10591), .Y(n8639) );
  MUX2X1 U9227 ( .B(n8643), .A(n8644), .S(n10591), .Y(n8642) );
  MUX2X1 U9228 ( .B(n8646), .A(n8647), .S(n10591), .Y(n8645) );
  MUX2X1 U9229 ( .B(n8649), .A(n8650), .S(n10565), .Y(n8648) );
  MUX2X1 U9230 ( .B(n8652), .A(n8653), .S(n10592), .Y(n8651) );
  MUX2X1 U9231 ( .B(n8655), .A(n8656), .S(n10592), .Y(n8654) );
  MUX2X1 U9232 ( .B(n8658), .A(n8659), .S(n10592), .Y(n8657) );
  MUX2X1 U9233 ( .B(n8661), .A(n8662), .S(n10592), .Y(n8660) );
  MUX2X1 U9234 ( .B(n8664), .A(n8665), .S(n10565), .Y(n8663) );
  MUX2X1 U9235 ( .B(n8667), .A(n8668), .S(n10592), .Y(n8666) );
  MUX2X1 U9236 ( .B(n8670), .A(n8671), .S(n10592), .Y(n8669) );
  MUX2X1 U9237 ( .B(n8673), .A(n8674), .S(n10592), .Y(n8672) );
  MUX2X1 U9238 ( .B(n8676), .A(n8677), .S(n10592), .Y(n8675) );
  MUX2X1 U9239 ( .B(n8679), .A(n8680), .S(read2_addr[1]), .Y(n8678) );
  MUX2X1 U9240 ( .B(n8682), .A(n8683), .S(n10592), .Y(n8681) );
  MUX2X1 U9241 ( .B(n8685), .A(n8686), .S(n10592), .Y(n8684) );
  MUX2X1 U9242 ( .B(n8688), .A(n8689), .S(n10592), .Y(n8687) );
  MUX2X1 U9243 ( .B(n8691), .A(n8692), .S(n10592), .Y(n8690) );
  MUX2X1 U9244 ( .B(n8694), .A(n8695), .S(n10564), .Y(n8693) );
  MUX2X1 U9245 ( .B(n8697), .A(n8698), .S(n10593), .Y(n8696) );
  MUX2X1 U9246 ( .B(n8700), .A(n8701), .S(n10593), .Y(n8699) );
  MUX2X1 U9247 ( .B(n8703), .A(n8704), .S(n10593), .Y(n8702) );
  MUX2X1 U9248 ( .B(n8706), .A(n8707), .S(n10593), .Y(n8705) );
  MUX2X1 U9249 ( .B(n8709), .A(n8710), .S(n10563), .Y(n8708) );
  MUX2X1 U9250 ( .B(n8712), .A(n8713), .S(n10593), .Y(n8711) );
  MUX2X1 U9251 ( .B(n8715), .A(n8716), .S(n10593), .Y(n8714) );
  MUX2X1 U9252 ( .B(n8718), .A(n8719), .S(n10593), .Y(n8717) );
  MUX2X1 U9253 ( .B(n8721), .A(n8722), .S(n10593), .Y(n8720) );
  MUX2X1 U9254 ( .B(n8724), .A(n8725), .S(n10563), .Y(n8723) );
  MUX2X1 U9255 ( .B(n8727), .A(n8728), .S(n10593), .Y(n8726) );
  MUX2X1 U9256 ( .B(n8730), .A(n8731), .S(n10593), .Y(n8729) );
  MUX2X1 U9257 ( .B(n8733), .A(n8734), .S(n10593), .Y(n8732) );
  MUX2X1 U9258 ( .B(n8736), .A(n8737), .S(n10593), .Y(n8735) );
  MUX2X1 U9259 ( .B(n8739), .A(n8740), .S(n10563), .Y(n8738) );
  MUX2X1 U9260 ( .B(n8742), .A(n8743), .S(n10594), .Y(n8741) );
  MUX2X1 U9261 ( .B(n8745), .A(n8746), .S(n10594), .Y(n8744) );
  MUX2X1 U9262 ( .B(n8748), .A(n8749), .S(n10594), .Y(n8747) );
  MUX2X1 U9263 ( .B(n8751), .A(n8752), .S(n10594), .Y(n8750) );
  MUX2X1 U9264 ( .B(n8754), .A(n8755), .S(n10563), .Y(n8753) );
  MUX2X1 U9265 ( .B(n8757), .A(n8758), .S(n10594), .Y(n8756) );
  MUX2X1 U9266 ( .B(n8760), .A(n8761), .S(n10594), .Y(n8759) );
  MUX2X1 U9267 ( .B(n8763), .A(n8764), .S(n10594), .Y(n8762) );
  MUX2X1 U9268 ( .B(n8766), .A(n8767), .S(n10594), .Y(n8765) );
  MUX2X1 U9269 ( .B(n8769), .A(n8770), .S(n10563), .Y(n8768) );
  MUX2X1 U9270 ( .B(n8772), .A(n8773), .S(n10594), .Y(n8771) );
  MUX2X1 U9271 ( .B(n8775), .A(n8776), .S(n10594), .Y(n8774) );
  MUX2X1 U9272 ( .B(n8778), .A(n8779), .S(n10594), .Y(n8777) );
  MUX2X1 U9273 ( .B(n8781), .A(n8782), .S(n10594), .Y(n8780) );
  MUX2X1 U9274 ( .B(n8784), .A(n8785), .S(n10563), .Y(n8783) );
  MUX2X1 U9275 ( .B(n8787), .A(n8788), .S(n10595), .Y(n8786) );
  MUX2X1 U9276 ( .B(n8790), .A(n8791), .S(n10595), .Y(n8789) );
  MUX2X1 U9277 ( .B(n8793), .A(n8794), .S(n10595), .Y(n8792) );
  MUX2X1 U9278 ( .B(n8796), .A(n8797), .S(n10595), .Y(n8795) );
  MUX2X1 U9279 ( .B(n8799), .A(n8800), .S(n10563), .Y(n8798) );
  MUX2X1 U9280 ( .B(n8802), .A(n8803), .S(n10595), .Y(n8801) );
  MUX2X1 U9281 ( .B(n8805), .A(n8806), .S(n10595), .Y(n8804) );
  MUX2X1 U9282 ( .B(n8808), .A(n8809), .S(n10595), .Y(n8807) );
  MUX2X1 U9283 ( .B(n8811), .A(n8812), .S(n10595), .Y(n8810) );
  MUX2X1 U9284 ( .B(n8814), .A(n8815), .S(n10563), .Y(n8813) );
  MUX2X1 U9285 ( .B(n8817), .A(n8818), .S(n10595), .Y(n8816) );
  MUX2X1 U9286 ( .B(n8820), .A(n8821), .S(n10595), .Y(n8819) );
  MUX2X1 U9287 ( .B(n8823), .A(n8824), .S(n10595), .Y(n8822) );
  MUX2X1 U9288 ( .B(n8826), .A(n8827), .S(n10595), .Y(n8825) );
  MUX2X1 U9289 ( .B(n8829), .A(n8830), .S(n10563), .Y(n8828) );
  MUX2X1 U9290 ( .B(n8832), .A(n8833), .S(n10596), .Y(n8831) );
  MUX2X1 U9291 ( .B(n8835), .A(n8836), .S(n10596), .Y(n8834) );
  MUX2X1 U9292 ( .B(n8838), .A(n8839), .S(n10596), .Y(n8837) );
  MUX2X1 U9293 ( .B(n8841), .A(n8842), .S(n10596), .Y(n8840) );
  MUX2X1 U9294 ( .B(n8844), .A(n8845), .S(n10563), .Y(n8843) );
  MUX2X1 U9295 ( .B(n8847), .A(n8848), .S(n10596), .Y(n8846) );
  MUX2X1 U9296 ( .B(n8850), .A(n8851), .S(n10596), .Y(n8849) );
  MUX2X1 U9297 ( .B(n8853), .A(n8854), .S(n10596), .Y(n8852) );
  MUX2X1 U9298 ( .B(n8856), .A(n8857), .S(n10596), .Y(n8855) );
  MUX2X1 U9299 ( .B(n8859), .A(n8860), .S(n10563), .Y(n8858) );
  MUX2X1 U9300 ( .B(n8862), .A(n8863), .S(n10596), .Y(n8861) );
  MUX2X1 U9301 ( .B(n8865), .A(n8866), .S(n10596), .Y(n8864) );
  MUX2X1 U9302 ( .B(n8868), .A(n8869), .S(n10596), .Y(n8867) );
  MUX2X1 U9303 ( .B(n8871), .A(n8872), .S(n10596), .Y(n8870) );
  MUX2X1 U9304 ( .B(n8874), .A(n8875), .S(n10563), .Y(n8873) );
  MUX2X1 U9305 ( .B(n8877), .A(n8878), .S(n10597), .Y(n8876) );
  MUX2X1 U9306 ( .B(n8880), .A(n8881), .S(n10597), .Y(n8879) );
  MUX2X1 U9307 ( .B(n8883), .A(n8884), .S(n10597), .Y(n8882) );
  MUX2X1 U9308 ( .B(n8886), .A(n8887), .S(n10597), .Y(n8885) );
  MUX2X1 U9309 ( .B(n8889), .A(n8890), .S(n10564), .Y(n8888) );
  MUX2X1 U9310 ( .B(n8892), .A(n8893), .S(n10597), .Y(n8891) );
  MUX2X1 U9311 ( .B(n8895), .A(n8896), .S(n10597), .Y(n8894) );
  MUX2X1 U9312 ( .B(n8898), .A(n8899), .S(n10597), .Y(n8897) );
  MUX2X1 U9313 ( .B(n8901), .A(n8902), .S(n10597), .Y(n8900) );
  MUX2X1 U9314 ( .B(n8904), .A(n8905), .S(n10564), .Y(n8903) );
  MUX2X1 U9315 ( .B(n8907), .A(n8908), .S(n10597), .Y(n8906) );
  MUX2X1 U9316 ( .B(n8910), .A(n8911), .S(n10597), .Y(n8909) );
  MUX2X1 U9317 ( .B(n8913), .A(n8914), .S(n10597), .Y(n8912) );
  MUX2X1 U9318 ( .B(n8916), .A(n8917), .S(n10597), .Y(n8915) );
  MUX2X1 U9319 ( .B(n8919), .A(n8920), .S(n10564), .Y(n8918) );
  MUX2X1 U9320 ( .B(n8922), .A(n8923), .S(n10598), .Y(n8921) );
  MUX2X1 U9321 ( .B(n8925), .A(n8926), .S(n10598), .Y(n8924) );
  MUX2X1 U9322 ( .B(n8928), .A(n8929), .S(n10598), .Y(n8927) );
  MUX2X1 U9323 ( .B(n8931), .A(n8932), .S(n10598), .Y(n8930) );
  MUX2X1 U9324 ( .B(n8934), .A(n8935), .S(n10564), .Y(n8933) );
  MUX2X1 U9325 ( .B(n8937), .A(n8938), .S(n10598), .Y(n8936) );
  MUX2X1 U9326 ( .B(n8940), .A(n8941), .S(n10598), .Y(n8939) );
  MUX2X1 U9327 ( .B(n8943), .A(n8944), .S(n10598), .Y(n8942) );
  MUX2X1 U9328 ( .B(n8946), .A(n8947), .S(n10598), .Y(n8945) );
  MUX2X1 U9329 ( .B(n8949), .A(n8950), .S(n10564), .Y(n8948) );
  MUX2X1 U9330 ( .B(n8952), .A(n8953), .S(n10598), .Y(n8951) );
  MUX2X1 U9331 ( .B(n8955), .A(n8956), .S(n10598), .Y(n8954) );
  MUX2X1 U9332 ( .B(n8958), .A(n8959), .S(n10598), .Y(n8957) );
  MUX2X1 U9333 ( .B(n8961), .A(n8962), .S(n10598), .Y(n8960) );
  MUX2X1 U9334 ( .B(n8964), .A(n8965), .S(n10564), .Y(n8963) );
  MUX2X1 U9335 ( .B(n8967), .A(n8968), .S(n10599), .Y(n8966) );
  MUX2X1 U9336 ( .B(n8970), .A(n8971), .S(n10599), .Y(n8969) );
  MUX2X1 U9337 ( .B(n8973), .A(n8974), .S(n10599), .Y(n8972) );
  MUX2X1 U9338 ( .B(n8976), .A(n8977), .S(n10599), .Y(n8975) );
  MUX2X1 U9339 ( .B(n8979), .A(n8980), .S(n10564), .Y(n8978) );
  MUX2X1 U9340 ( .B(n8982), .A(n8983), .S(n10599), .Y(n8981) );
  MUX2X1 U9341 ( .B(n8985), .A(n8986), .S(n10599), .Y(n8984) );
  MUX2X1 U9342 ( .B(n8988), .A(n8989), .S(n10599), .Y(n8987) );
  MUX2X1 U9343 ( .B(n8991), .A(n8992), .S(n10599), .Y(n8990) );
  MUX2X1 U9344 ( .B(n8994), .A(n8995), .S(n10564), .Y(n8993) );
  MUX2X1 U9345 ( .B(n8997), .A(n8998), .S(n10599), .Y(n8996) );
  MUX2X1 U9346 ( .B(n9000), .A(n9001), .S(n10599), .Y(n8999) );
  MUX2X1 U9347 ( .B(n9003), .A(n9004), .S(n10599), .Y(n9002) );
  MUX2X1 U9348 ( .B(n9006), .A(n9007), .S(n10599), .Y(n9005) );
  MUX2X1 U9349 ( .B(n9009), .A(n9010), .S(n10564), .Y(n9008) );
  MUX2X1 U9350 ( .B(n9012), .A(n9013), .S(n10600), .Y(n9011) );
  MUX2X1 U9351 ( .B(n9015), .A(n9016), .S(n10600), .Y(n9014) );
  MUX2X1 U9352 ( .B(n9018), .A(n9019), .S(n10600), .Y(n9017) );
  MUX2X1 U9353 ( .B(n9021), .A(n9022), .S(n10600), .Y(n9020) );
  MUX2X1 U9354 ( .B(n9024), .A(n9025), .S(n10564), .Y(n9023) );
  MUX2X1 U9355 ( .B(n9027), .A(n9028), .S(n10600), .Y(n9026) );
  MUX2X1 U9356 ( .B(n9030), .A(n9031), .S(n10600), .Y(n9029) );
  MUX2X1 U9357 ( .B(n9033), .A(n9034), .S(n10600), .Y(n9032) );
  MUX2X1 U9358 ( .B(n9036), .A(n9037), .S(n10600), .Y(n9035) );
  MUX2X1 U9359 ( .B(n9039), .A(n9040), .S(n10564), .Y(n9038) );
  MUX2X1 U9360 ( .B(n9042), .A(n9043), .S(n10600), .Y(n9041) );
  MUX2X1 U9361 ( .B(n9045), .A(n9046), .S(n10600), .Y(n9044) );
  MUX2X1 U9362 ( .B(n9048), .A(n9049), .S(n10600), .Y(n9047) );
  MUX2X1 U9363 ( .B(n9051), .A(n9052), .S(n10600), .Y(n9050) );
  MUX2X1 U9364 ( .B(n9054), .A(n9055), .S(n10564), .Y(n9053) );
  MUX2X1 U9365 ( .B(n9057), .A(n9058), .S(n10601), .Y(n9056) );
  MUX2X1 U9366 ( .B(n9060), .A(n9061), .S(n10601), .Y(n9059) );
  MUX2X1 U9367 ( .B(n9063), .A(n9064), .S(n10601), .Y(n9062) );
  MUX2X1 U9368 ( .B(n9066), .A(n9067), .S(n10601), .Y(n9065) );
  MUX2X1 U9369 ( .B(n9069), .A(n9070), .S(n10565), .Y(n9068) );
  MUX2X1 U9370 ( .B(n9072), .A(n9073), .S(n10601), .Y(n9071) );
  MUX2X1 U9371 ( .B(n9075), .A(n9076), .S(n10601), .Y(n9074) );
  MUX2X1 U9372 ( .B(n9078), .A(n9079), .S(n10601), .Y(n9077) );
  MUX2X1 U9373 ( .B(n9081), .A(n9082), .S(n10601), .Y(n9080) );
  MUX2X1 U9374 ( .B(n9084), .A(n9085), .S(n10565), .Y(n9083) );
  MUX2X1 U9375 ( .B(n9087), .A(n9088), .S(n10601), .Y(n9086) );
  MUX2X1 U9376 ( .B(n9090), .A(n9091), .S(n10601), .Y(n9089) );
  MUX2X1 U9377 ( .B(n9093), .A(n9094), .S(n10601), .Y(n9092) );
  MUX2X1 U9378 ( .B(n9096), .A(n9097), .S(n10601), .Y(n9095) );
  MUX2X1 U9379 ( .B(n9099), .A(n9100), .S(n10565), .Y(n9098) );
  MUX2X1 U9380 ( .B(n9102), .A(n9103), .S(n10602), .Y(n9101) );
  MUX2X1 U9381 ( .B(n9105), .A(n9106), .S(n10602), .Y(n9104) );
  MUX2X1 U9382 ( .B(n9108), .A(n9109), .S(n10602), .Y(n9107) );
  MUX2X1 U9383 ( .B(n9111), .A(n9112), .S(n10602), .Y(n9110) );
  MUX2X1 U9384 ( .B(n9114), .A(n9115), .S(n10565), .Y(n9113) );
  MUX2X1 U9385 ( .B(n9117), .A(n9118), .S(n10602), .Y(n9116) );
  MUX2X1 U9386 ( .B(n9120), .A(n9121), .S(n10602), .Y(n9119) );
  MUX2X1 U9387 ( .B(n9123), .A(n9124), .S(n10602), .Y(n9122) );
  MUX2X1 U9388 ( .B(n9126), .A(n9127), .S(n10602), .Y(n9125) );
  MUX2X1 U9389 ( .B(n9129), .A(n9130), .S(n10565), .Y(n9128) );
  MUX2X1 U9390 ( .B(n9132), .A(n9133), .S(n10602), .Y(n9131) );
  MUX2X1 U9391 ( .B(n9135), .A(n9136), .S(n10602), .Y(n9134) );
  MUX2X1 U9392 ( .B(n9138), .A(n9139), .S(n10602), .Y(n9137) );
  MUX2X1 U9393 ( .B(n9141), .A(n9142), .S(n10602), .Y(n9140) );
  MUX2X1 U9394 ( .B(n9144), .A(n9145), .S(n10565), .Y(n9143) );
  MUX2X1 U9395 ( .B(n9147), .A(n9148), .S(n10603), .Y(n9146) );
  MUX2X1 U9396 ( .B(n9150), .A(n9151), .S(n10603), .Y(n9149) );
  MUX2X1 U9397 ( .B(n9153), .A(n9154), .S(n10603), .Y(n9152) );
  MUX2X1 U9398 ( .B(n9156), .A(n9157), .S(n10603), .Y(n9155) );
  MUX2X1 U9399 ( .B(n9159), .A(n9160), .S(n10565), .Y(n9158) );
  MUX2X1 U9400 ( .B(n9162), .A(n9163), .S(n10603), .Y(n9161) );
  MUX2X1 U9401 ( .B(n9165), .A(n9166), .S(n10603), .Y(n9164) );
  MUX2X1 U9402 ( .B(n9168), .A(n9169), .S(n10603), .Y(n9167) );
  MUX2X1 U9403 ( .B(n9171), .A(n9172), .S(n10603), .Y(n9170) );
  MUX2X1 U9404 ( .B(n9174), .A(n9175), .S(n10565), .Y(n9173) );
  MUX2X1 U9405 ( .B(n9177), .A(n9178), .S(n10603), .Y(n9176) );
  MUX2X1 U9406 ( .B(n9180), .A(n9181), .S(n10603), .Y(n9179) );
  MUX2X1 U9407 ( .B(n9183), .A(n9184), .S(n10603), .Y(n9182) );
  MUX2X1 U9408 ( .B(n9186), .A(n9187), .S(n10603), .Y(n9185) );
  MUX2X1 U9409 ( .B(n9189), .A(n9190), .S(n10565), .Y(n9188) );
  MUX2X1 U9410 ( .B(n9192), .A(n9193), .S(n10604), .Y(n9191) );
  MUX2X1 U9411 ( .B(n9195), .A(n9196), .S(n10604), .Y(n9194) );
  MUX2X1 U9412 ( .B(n9198), .A(n9199), .S(n10604), .Y(n9197) );
  MUX2X1 U9413 ( .B(n9201), .A(n9202), .S(n10604), .Y(n9200) );
  MUX2X1 U9414 ( .B(n9204), .A(n9205), .S(n10565), .Y(n9203) );
  MUX2X1 U9415 ( .B(n9207), .A(n9208), .S(n10604), .Y(n9206) );
  MUX2X1 U9416 ( .B(n9210), .A(n9211), .S(n10604), .Y(n9209) );
  MUX2X1 U9417 ( .B(n9213), .A(n9214), .S(n10604), .Y(n9212) );
  MUX2X1 U9418 ( .B(n9216), .A(n9217), .S(n10604), .Y(n9215) );
  MUX2X1 U9419 ( .B(n9219), .A(n9220), .S(n10565), .Y(n9218) );
  MUX2X1 U9420 ( .B(n9222), .A(n9223), .S(n10604), .Y(n9221) );
  MUX2X1 U9421 ( .B(n9225), .A(n9226), .S(n10604), .Y(n9224) );
  MUX2X1 U9422 ( .B(n9228), .A(n9229), .S(n10604), .Y(n9227) );
  MUX2X1 U9423 ( .B(n9231), .A(n9232), .S(n10604), .Y(n9230) );
  MUX2X1 U9424 ( .B(n9234), .A(n9235), .S(n10565), .Y(n9233) );
  MUX2X1 U9425 ( .B(n9237), .A(n9238), .S(n10605), .Y(n9236) );
  MUX2X1 U9426 ( .B(n9240), .A(n9241), .S(n10605), .Y(n9239) );
  MUX2X1 U9427 ( .B(n9243), .A(n9244), .S(n10605), .Y(n9242) );
  MUX2X1 U9428 ( .B(n9246), .A(n9247), .S(n10605), .Y(n9245) );
  MUX2X1 U9429 ( .B(n9249), .A(n9250), .S(read2_addr[1]), .Y(n9248) );
  MUX2X1 U9430 ( .B(n9252), .A(n9253), .S(n10605), .Y(n9251) );
  MUX2X1 U9431 ( .B(n9255), .A(n9256), .S(n10605), .Y(n9254) );
  MUX2X1 U9432 ( .B(n9258), .A(n9259), .S(n10605), .Y(n9257) );
  MUX2X1 U9433 ( .B(n9261), .A(n9262), .S(n10605), .Y(n9260) );
  MUX2X1 U9434 ( .B(n9264), .A(n9265), .S(read2_addr[1]), .Y(n9263) );
  MUX2X1 U9435 ( .B(n9267), .A(n9268), .S(n10605), .Y(n9266) );
  MUX2X1 U9436 ( .B(n9270), .A(n9271), .S(n10605), .Y(n9269) );
  MUX2X1 U9437 ( .B(n9273), .A(n9274), .S(n10605), .Y(n9272) );
  MUX2X1 U9438 ( .B(n9276), .A(n9277), .S(n10605), .Y(n9275) );
  MUX2X1 U9439 ( .B(n9279), .A(n9280), .S(read2_addr[1]), .Y(n9278) );
  MUX2X1 U9440 ( .B(n9282), .A(n9283), .S(n10606), .Y(n9281) );
  MUX2X1 U9441 ( .B(n9285), .A(n9286), .S(n10606), .Y(n9284) );
  MUX2X1 U9442 ( .B(n9288), .A(n9289), .S(n10606), .Y(n9287) );
  MUX2X1 U9443 ( .B(n9291), .A(n9292), .S(n10606), .Y(n9290) );
  MUX2X1 U9444 ( .B(n9294), .A(n9295), .S(read2_addr[1]), .Y(n9293) );
  MUX2X1 U9445 ( .B(n9297), .A(n9298), .S(n10606), .Y(n9296) );
  MUX2X1 U9446 ( .B(n9300), .A(n9301), .S(n10606), .Y(n9299) );
  MUX2X1 U9447 ( .B(n9303), .A(n9304), .S(n10606), .Y(n9302) );
  MUX2X1 U9448 ( .B(n9306), .A(n9307), .S(n10606), .Y(n9305) );
  MUX2X1 U9449 ( .B(n9309), .A(n9310), .S(read2_addr[1]), .Y(n9308) );
  MUX2X1 U9450 ( .B(n9312), .A(n9313), .S(n10606), .Y(n9311) );
  MUX2X1 U9451 ( .B(n9315), .A(n9316), .S(n10606), .Y(n9314) );
  MUX2X1 U9452 ( .B(n9318), .A(n9319), .S(n10606), .Y(n9317) );
  MUX2X1 U9453 ( .B(n9321), .A(n9322), .S(n10606), .Y(n9320) );
  MUX2X1 U9454 ( .B(n9324), .A(n9325), .S(read2_addr[1]), .Y(n9323) );
  MUX2X1 U9455 ( .B(n9327), .A(n9328), .S(n10607), .Y(n9326) );
  MUX2X1 U9456 ( .B(n9330), .A(n9331), .S(n10607), .Y(n9329) );
  MUX2X1 U9457 ( .B(n9333), .A(n9334), .S(n10607), .Y(n9332) );
  MUX2X1 U9458 ( .B(n9336), .A(n9337), .S(n10607), .Y(n9335) );
  MUX2X1 U9459 ( .B(n9339), .A(n9340), .S(read2_addr[1]), .Y(n9338) );
  MUX2X1 U9460 ( .B(n9342), .A(n9343), .S(n10607), .Y(n9341) );
  MUX2X1 U9461 ( .B(n9345), .A(n9346), .S(n10607), .Y(n9344) );
  MUX2X1 U9462 ( .B(n9348), .A(n9349), .S(n10607), .Y(n9347) );
  MUX2X1 U9463 ( .B(n9351), .A(n9352), .S(n10607), .Y(n9350) );
  MUX2X1 U9464 ( .B(n9354), .A(n9355), .S(read2_addr[1]), .Y(n9353) );
  MUX2X1 U9465 ( .B(n9357), .A(n9358), .S(n10607), .Y(n9356) );
  MUX2X1 U9466 ( .B(n9360), .A(n9361), .S(n10607), .Y(n9359) );
  MUX2X1 U9467 ( .B(n9363), .A(n9364), .S(n10607), .Y(n9362) );
  MUX2X1 U9468 ( .B(n9366), .A(n9367), .S(n10607), .Y(n9365) );
  MUX2X1 U9469 ( .B(n9369), .A(n9370), .S(read2_addr[1]), .Y(n9368) );
  MUX2X1 U9470 ( .B(n9372), .A(n9373), .S(n10608), .Y(n9371) );
  MUX2X1 U9471 ( .B(n9375), .A(n9376), .S(n10608), .Y(n9374) );
  MUX2X1 U9472 ( .B(n9378), .A(n9379), .S(n10608), .Y(n9377) );
  MUX2X1 U9473 ( .B(n9381), .A(n9382), .S(n10608), .Y(n9380) );
  MUX2X1 U9474 ( .B(n9384), .A(n9385), .S(read2_addr[1]), .Y(n9383) );
  MUX2X1 U9475 ( .B(n9387), .A(n9388), .S(n10608), .Y(n9386) );
  MUX2X1 U9476 ( .B(n9390), .A(n9391), .S(n10608), .Y(n9389) );
  MUX2X1 U9477 ( .B(n9393), .A(n9394), .S(n10608), .Y(n9392) );
  MUX2X1 U9478 ( .B(n9396), .A(n9397), .S(n10608), .Y(n9395) );
  MUX2X1 U9479 ( .B(n9399), .A(n9400), .S(read2_addr[1]), .Y(n9398) );
  MUX2X1 U9480 ( .B(n9402), .A(n9403), .S(n10608), .Y(n9401) );
  MUX2X1 U9481 ( .B(n9405), .A(n9406), .S(n10608), .Y(n9404) );
  MUX2X1 U9482 ( .B(n9408), .A(n9409), .S(n10608), .Y(n9407) );
  MUX2X1 U9483 ( .B(n9411), .A(n9412), .S(n10608), .Y(n9410) );
  MUX2X1 U9484 ( .B(n9414), .A(n9415), .S(read2_addr[1]), .Y(n9413) );
  MUX2X1 U9485 ( .B(n9417), .A(n9418), .S(n10609), .Y(n9416) );
  MUX2X1 U9486 ( .B(n9420), .A(n9421), .S(n10609), .Y(n9419) );
  MUX2X1 U9487 ( .B(n9423), .A(n9424), .S(n10609), .Y(n9422) );
  MUX2X1 U9488 ( .B(n9426), .A(n9427), .S(n10609), .Y(n9425) );
  MUX2X1 U9489 ( .B(n9429), .A(n9430), .S(n10565), .Y(n9428) );
  MUX2X1 U9490 ( .B(n9432), .A(n9433), .S(n10609), .Y(n9431) );
  MUX2X1 U9491 ( .B(n9435), .A(n9436), .S(n10609), .Y(n9434) );
  MUX2X1 U9492 ( .B(n9438), .A(n9439), .S(n10609), .Y(n9437) );
  MUX2X1 U9493 ( .B(n9441), .A(n9442), .S(n10609), .Y(n9440) );
  MUX2X1 U9494 ( .B(n9444), .A(n9445), .S(n10564), .Y(n9443) );
  MUX2X1 U9495 ( .B(n9447), .A(n9448), .S(n10609), .Y(n9446) );
  MUX2X1 U9496 ( .B(n9450), .A(n9451), .S(n10609), .Y(n9449) );
  MUX2X1 U9497 ( .B(n9453), .A(n9454), .S(n10609), .Y(n9452) );
  MUX2X1 U9498 ( .B(n9456), .A(n9457), .S(n10609), .Y(n9455) );
  MUX2X1 U9499 ( .B(n9459), .A(n9460), .S(n10563), .Y(n9458) );
  MUX2X1 U9500 ( .B(n9462), .A(n9463), .S(n10610), .Y(n9461) );
  MUX2X1 U9501 ( .B(n9465), .A(n9466), .S(n10610), .Y(n9464) );
  MUX2X1 U9502 ( .B(n9468), .A(n9469), .S(n10610), .Y(n9467) );
  MUX2X1 U9503 ( .B(n9471), .A(n9472), .S(n10610), .Y(n9470) );
  MUX2X1 U9504 ( .B(n9474), .A(n9475), .S(read2_addr[1]), .Y(n9473) );
  MUX2X1 U9505 ( .B(n9477), .A(n9478), .S(n10610), .Y(n9476) );
  MUX2X1 U9506 ( .B(n9480), .A(n9481), .S(n10610), .Y(n9479) );
  MUX2X1 U9507 ( .B(n9483), .A(n9484), .S(n10610), .Y(n9482) );
  MUX2X1 U9508 ( .B(n9486), .A(n9487), .S(n10610), .Y(n9485) );
  MUX2X1 U9509 ( .B(n9489), .A(n9490), .S(n10564), .Y(n9488) );
  MUX2X1 U9510 ( .B(n9492), .A(n9493), .S(n10610), .Y(n9491) );
  MUX2X1 U9511 ( .B(n9495), .A(n9496), .S(n10610), .Y(n9494) );
  MUX2X1 U9512 ( .B(n9498), .A(n9499), .S(n10610), .Y(n9497) );
  MUX2X1 U9513 ( .B(n9501), .A(n9502), .S(n10610), .Y(n9500) );
  MUX2X1 U9514 ( .B(n9504), .A(n9505), .S(n10565), .Y(n9503) );
  MUX2X1 U9515 ( .B(n9507), .A(n9508), .S(n10611), .Y(n9506) );
  MUX2X1 U9516 ( .B(n9510), .A(n9511), .S(n10611), .Y(n9509) );
  MUX2X1 U9517 ( .B(n9513), .A(n9514), .S(n10611), .Y(n9512) );
  MUX2X1 U9518 ( .B(n9516), .A(n9517), .S(n10611), .Y(n9515) );
  MUX2X1 U9519 ( .B(n9519), .A(n9520), .S(read2_addr[1]), .Y(n9518) );
  MUX2X1 U9520 ( .B(n9522), .A(n9523), .S(n10611), .Y(n9521) );
  MUX2X1 U9521 ( .B(n9525), .A(n9526), .S(n10611), .Y(n9524) );
  MUX2X1 U9522 ( .B(n9528), .A(n9529), .S(n10611), .Y(n9527) );
  MUX2X1 U9523 ( .B(n9531), .A(n9532), .S(n10611), .Y(n9530) );
  MUX2X1 U9524 ( .B(n9534), .A(n9535), .S(n10563), .Y(n9533) );
  MUX2X1 U9525 ( .B(n9537), .A(n9538), .S(n10611), .Y(n9536) );
  MUX2X1 U9526 ( .B(n9540), .A(n9541), .S(n10611), .Y(n9539) );
  MUX2X1 U9527 ( .B(n9543), .A(n9544), .S(n10611), .Y(n9542) );
  MUX2X1 U9528 ( .B(n9546), .A(n9547), .S(n10611), .Y(n9545) );
  MUX2X1 U9529 ( .B(n9549), .A(n9550), .S(n10565), .Y(n9548) );
  MUX2X1 U9530 ( .B(n9552), .A(n9553), .S(n10612), .Y(n9551) );
  MUX2X1 U9531 ( .B(n9555), .A(n9556), .S(n10612), .Y(n9554) );
  MUX2X1 U9532 ( .B(n9558), .A(n9559), .S(n10612), .Y(n9557) );
  MUX2X1 U9533 ( .B(n9561), .A(n9562), .S(n10612), .Y(n9560) );
  MUX2X1 U9534 ( .B(n9564), .A(n9565), .S(n10564), .Y(n9563) );
  MUX2X1 U9535 ( .B(n9567), .A(n9568), .S(n10612), .Y(n9566) );
  MUX2X1 U9536 ( .B(n9570), .A(n9571), .S(n10612), .Y(n9569) );
  MUX2X1 U9537 ( .B(n9573), .A(n9574), .S(n10612), .Y(n9572) );
  MUX2X1 U9538 ( .B(n9576), .A(n9577), .S(n10612), .Y(n9575) );
  MUX2X1 U9539 ( .B(n9579), .A(n9580), .S(n10563), .Y(n9578) );
  MUX2X1 U9540 ( .B(n9582), .A(n9583), .S(n10612), .Y(n9581) );
  MUX2X1 U9541 ( .B(n9585), .A(n9586), .S(n10612), .Y(n9584) );
  MUX2X1 U9542 ( .B(n9588), .A(n9589), .S(n10612), .Y(n9587) );
  MUX2X1 U9543 ( .B(n9591), .A(n9592), .S(n10612), .Y(n9590) );
  MUX2X1 U9544 ( .B(n9594), .A(n9595), .S(read2_addr[1]), .Y(n9593) );
  MUX2X1 U9545 ( .B(n9597), .A(n9598), .S(n10613), .Y(n9596) );
  MUX2X1 U9546 ( .B(n9600), .A(n9601), .S(n10613), .Y(n9599) );
  MUX2X1 U9547 ( .B(n9603), .A(n9604), .S(n10613), .Y(n9602) );
  MUX2X1 U9548 ( .B(n9606), .A(n9607), .S(n10613), .Y(n9605) );
  MUX2X1 U9549 ( .B(n9609), .A(n9610), .S(n10563), .Y(n9608) );
  MUX2X1 U9550 ( .B(n9612), .A(n9613), .S(n10613), .Y(n9611) );
  MUX2X1 U9551 ( .B(n9615), .A(n9616), .S(n10613), .Y(n9614) );
  MUX2X1 U9552 ( .B(n9618), .A(n9619), .S(n10613), .Y(n9617) );
  MUX2X1 U9553 ( .B(n9621), .A(n9622), .S(n10613), .Y(n9620) );
  MUX2X1 U9554 ( .B(n9624), .A(n9625), .S(read2_addr[1]), .Y(n9623) );
  MUX2X1 U9555 ( .B(n9627), .A(n9628), .S(n10613), .Y(n9626) );
  MUX2X1 U9556 ( .B(n9630), .A(n9631), .S(n10613), .Y(n9629) );
  MUX2X1 U9557 ( .B(n9633), .A(n9634), .S(n10613), .Y(n9632) );
  MUX2X1 U9558 ( .B(n9636), .A(n9637), .S(n10613), .Y(n9635) );
  MUX2X1 U9559 ( .B(n9639), .A(n9640), .S(read2_addr[1]), .Y(n9638) );
  MUX2X1 U9560 ( .B(n9642), .A(n9643), .S(n10614), .Y(n9641) );
  MUX2X1 U9561 ( .B(n9645), .A(n9646), .S(n10614), .Y(n9644) );
  MUX2X1 U9562 ( .B(n9648), .A(n9649), .S(n10614), .Y(n9647) );
  MUX2X1 U9563 ( .B(n9651), .A(n9652), .S(n10614), .Y(n9650) );
  MUX2X1 U9564 ( .B(n9654), .A(n9655), .S(read2_addr[1]), .Y(n9653) );
  MUX2X1 U9565 ( .B(n9657), .A(n9658), .S(n10614), .Y(n9656) );
  MUX2X1 U9566 ( .B(n9660), .A(n9661), .S(n10614), .Y(n9659) );
  MUX2X1 U9567 ( .B(n9663), .A(n9664), .S(n10614), .Y(n9662) );
  MUX2X1 U9568 ( .B(n9666), .A(n9667), .S(n10614), .Y(n9665) );
  MUX2X1 U9569 ( .B(n9669), .A(n9670), .S(n10565), .Y(n9668) );
  MUX2X1 U9570 ( .B(n9672), .A(n9673), .S(n10614), .Y(n9671) );
  MUX2X1 U9571 ( .B(n9675), .A(n9676), .S(n10614), .Y(n9674) );
  MUX2X1 U9572 ( .B(n9678), .A(n9679), .S(n10614), .Y(n9677) );
  MUX2X1 U9573 ( .B(n9681), .A(n9682), .S(n10614), .Y(n9680) );
  MUX2X1 U9574 ( .B(n9684), .A(n9685), .S(n10565), .Y(n9683) );
  MUX2X1 U9575 ( .B(n9687), .A(n9688), .S(n10615), .Y(n9686) );
  MUX2X1 U9576 ( .B(n9690), .A(n9691), .S(n10615), .Y(n9689) );
  MUX2X1 U9577 ( .B(n9693), .A(n9694), .S(n10615), .Y(n9692) );
  MUX2X1 U9578 ( .B(n9696), .A(n9697), .S(n10615), .Y(n9695) );
  MUX2X1 U9579 ( .B(n9699), .A(n9700), .S(n10563), .Y(n9698) );
  MUX2X1 U9580 ( .B(n9702), .A(n9703), .S(n10615), .Y(n9701) );
  MUX2X1 U9581 ( .B(n9705), .A(n9706), .S(n10615), .Y(n9704) );
  MUX2X1 U9582 ( .B(n9708), .A(n9709), .S(n10615), .Y(n9707) );
  MUX2X1 U9583 ( .B(n9711), .A(n9712), .S(n10615), .Y(n9710) );
  MUX2X1 U9584 ( .B(n9714), .A(n9715), .S(n10563), .Y(n9713) );
  MUX2X1 U9585 ( .B(n9717), .A(n9718), .S(n10615), .Y(n9716) );
  MUX2X1 U9586 ( .B(n9720), .A(n9721), .S(n10615), .Y(n9719) );
  MUX2X1 U9587 ( .B(n9723), .A(n9724), .S(n10615), .Y(n9722) );
  MUX2X1 U9588 ( .B(n9726), .A(n9727), .S(n10615), .Y(n9725) );
  MUX2X1 U9589 ( .B(n9729), .A(n9730), .S(n10564), .Y(n9728) );
  MUX2X1 U9590 ( .B(n9732), .A(n9733), .S(n10616), .Y(n9731) );
  MUX2X1 U9591 ( .B(n9735), .A(n9736), .S(n10616), .Y(n9734) );
  MUX2X1 U9592 ( .B(n9738), .A(n9739), .S(n10616), .Y(n9737) );
  MUX2X1 U9593 ( .B(n9741), .A(n9742), .S(n10616), .Y(n9740) );
  MUX2X1 U9594 ( .B(n9744), .A(n9745), .S(n10563), .Y(n9743) );
  MUX2X1 U9595 ( .B(n9747), .A(n9748), .S(n10616), .Y(n9746) );
  MUX2X1 U9596 ( .B(n9750), .A(n9751), .S(n10616), .Y(n9749) );
  MUX2X1 U9597 ( .B(n9753), .A(n9754), .S(n10616), .Y(n9752) );
  MUX2X1 U9598 ( .B(n9756), .A(n9757), .S(n10616), .Y(n9755) );
  MUX2X1 U9599 ( .B(n9759), .A(n9760), .S(n10564), .Y(n9758) );
  MUX2X1 U9600 ( .B(n9762), .A(n9763), .S(n10616), .Y(n9761) );
  MUX2X1 U9601 ( .B(n9765), .A(n9766), .S(n10616), .Y(n9764) );
  MUX2X1 U9602 ( .B(n9768), .A(n9769), .S(n10616), .Y(n9767) );
  MUX2X1 U9603 ( .B(n9771), .A(n9772), .S(n10616), .Y(n9770) );
  MUX2X1 U9604 ( .B(n9774), .A(n9775), .S(n10564), .Y(n9773) );
  MUX2X1 U9605 ( .B(n9777), .A(n9778), .S(n10617), .Y(n9776) );
  MUX2X1 U9606 ( .B(n9780), .A(n9781), .S(n10617), .Y(n9779) );
  MUX2X1 U9607 ( .B(n9783), .A(n9784), .S(n10617), .Y(n9782) );
  MUX2X1 U9608 ( .B(n9786), .A(n9787), .S(n10617), .Y(n9785) );
  MUX2X1 U9609 ( .B(n9789), .A(n9790), .S(n10564), .Y(n9788) );
  MUX2X1 U9610 ( .B(n9792), .A(n9793), .S(n10617), .Y(n9791) );
  MUX2X1 U9611 ( .B(n9795), .A(n9796), .S(n10617), .Y(n9794) );
  MUX2X1 U9612 ( .B(n9798), .A(n9799), .S(n10617), .Y(n9797) );
  MUX2X1 U9613 ( .B(n9801), .A(n9802), .S(n10617), .Y(n9800) );
  MUX2X1 U9614 ( .B(n9804), .A(n9805), .S(n10563), .Y(n9803) );
  MUX2X1 U9615 ( .B(n9807), .A(n9808), .S(n10617), .Y(n9806) );
  MUX2X1 U9616 ( .B(n9810), .A(n9811), .S(n10617), .Y(n9809) );
  MUX2X1 U9617 ( .B(n9813), .A(n9814), .S(n10617), .Y(n9812) );
  MUX2X1 U9618 ( .B(n9816), .A(n9817), .S(n10617), .Y(n9815) );
  MUX2X1 U9619 ( .B(n9819), .A(n9820), .S(n10563), .Y(n9818) );
  MUX2X1 U9620 ( .B(n9822), .A(n9823), .S(n10618), .Y(n9821) );
  MUX2X1 U9621 ( .B(n9825), .A(n9826), .S(n10618), .Y(n9824) );
  MUX2X1 U9622 ( .B(n9828), .A(n9829), .S(n10618), .Y(n9827) );
  MUX2X1 U9623 ( .B(n9831), .A(n9832), .S(n10618), .Y(n9830) );
  MUX2X1 U9624 ( .B(n9834), .A(n9835), .S(n10563), .Y(n9833) );
  MUX2X1 U9625 ( .B(n9837), .A(n9838), .S(n10618), .Y(n9836) );
  MUX2X1 U9626 ( .B(n9840), .A(n9841), .S(n10618), .Y(n9839) );
  MUX2X1 U9627 ( .B(n9843), .A(n9844), .S(n10618), .Y(n9842) );
  MUX2X1 U9628 ( .B(n9846), .A(n9847), .S(n10618), .Y(n9845) );
  MUX2X1 U9629 ( .B(n9849), .A(n9850), .S(n10563), .Y(n9848) );
  MUX2X1 U9630 ( .B(n9852), .A(n9853), .S(n10618), .Y(n9851) );
  MUX2X1 U9631 ( .B(n9855), .A(n9856), .S(n10618), .Y(n9854) );
  MUX2X1 U9632 ( .B(n9858), .A(n9859), .S(n10618), .Y(n9857) );
  MUX2X1 U9633 ( .B(n9861), .A(n9862), .S(n10618), .Y(n9860) );
  MUX2X1 U9634 ( .B(n9864), .A(n9865), .S(n10564), .Y(n9863) );
  MUX2X1 U9635 ( .B(n9867), .A(n9868), .S(n10619), .Y(n9866) );
  MUX2X1 U9636 ( .B(n9870), .A(n9871), .S(n10619), .Y(n9869) );
  MUX2X1 U9637 ( .B(n9873), .A(n9874), .S(n10619), .Y(n9872) );
  MUX2X1 U9638 ( .B(n9876), .A(n9877), .S(n10619), .Y(n9875) );
  MUX2X1 U9639 ( .B(n9879), .A(n9880), .S(read2_addr[1]), .Y(n9878) );
  MUX2X1 U9640 ( .B(n9882), .A(n9883), .S(n10619), .Y(n9881) );
  MUX2X1 U9641 ( .B(n9885), .A(n9886), .S(n10619), .Y(n9884) );
  MUX2X1 U9642 ( .B(n9888), .A(n9889), .S(n10619), .Y(n9887) );
  MUX2X1 U9643 ( .B(n9891), .A(n9892), .S(n10619), .Y(n9890) );
  MUX2X1 U9644 ( .B(n9894), .A(n9895), .S(n10564), .Y(n9893) );
  MUX2X1 U9645 ( .B(n9897), .A(n9898), .S(n10619), .Y(n9896) );
  MUX2X1 U9646 ( .B(n9900), .A(n9901), .S(n10619), .Y(n9899) );
  MUX2X1 U9647 ( .B(n9903), .A(n9904), .S(n10619), .Y(n9902) );
  MUX2X1 U9648 ( .B(n9906), .A(n9907), .S(n10619), .Y(n9905) );
  MUX2X1 U9649 ( .B(n9909), .A(n9910), .S(n10565), .Y(n9908) );
  MUX2X1 U9650 ( .B(n9912), .A(n9913), .S(n10620), .Y(n9911) );
  MUX2X1 U9651 ( .B(n9915), .A(n9916), .S(n10620), .Y(n9914) );
  MUX2X1 U9652 ( .B(n9918), .A(n9919), .S(n10620), .Y(n9917) );
  MUX2X1 U9653 ( .B(n9921), .A(n9922), .S(n10620), .Y(n9920) );
  MUX2X1 U9654 ( .B(n9924), .A(n9925), .S(n10563), .Y(n9923) );
  MUX2X1 U9655 ( .B(n9927), .A(n9928), .S(n10620), .Y(n9926) );
  MUX2X1 U9656 ( .B(n9930), .A(n9931), .S(n10620), .Y(n9929) );
  MUX2X1 U9657 ( .B(n9933), .A(n9934), .S(n10620), .Y(n9932) );
  MUX2X1 U9658 ( .B(n9936), .A(n9937), .S(n10620), .Y(n9935) );
  MUX2X1 U9659 ( .B(n9939), .A(n9940), .S(n10565), .Y(n9938) );
  MUX2X1 U9660 ( .B(n9942), .A(n9943), .S(n10620), .Y(n9941) );
  MUX2X1 U9661 ( .B(n9945), .A(n9946), .S(n10620), .Y(n9944) );
  MUX2X1 U9662 ( .B(n9948), .A(n9949), .S(n10620), .Y(n9947) );
  MUX2X1 U9663 ( .B(n9951), .A(n9952), .S(n10620), .Y(n9950) );
  MUX2X1 U9664 ( .B(n9954), .A(n9955), .S(read2_addr[1]), .Y(n9953) );
  MUX2X1 U9665 ( .B(n9957), .A(n9958), .S(n10621), .Y(n9956) );
  MUX2X1 U9666 ( .B(n9960), .A(n9961), .S(n10621), .Y(n9959) );
  MUX2X1 U9667 ( .B(n9963), .A(n9964), .S(n10621), .Y(n9962) );
  MUX2X1 U9668 ( .B(n9966), .A(n9967), .S(n10621), .Y(n9965) );
  MUX2X1 U9669 ( .B(n9969), .A(n9970), .S(n10564), .Y(n9968) );
  MUX2X1 U9670 ( .B(n9972), .A(n9973), .S(n10621), .Y(n9971) );
  MUX2X1 U9671 ( .B(n9975), .A(n9976), .S(n10621), .Y(n9974) );
  MUX2X1 U9672 ( .B(n9978), .A(n9979), .S(n10621), .Y(n9977) );
  MUX2X1 U9673 ( .B(n9981), .A(n9982), .S(n10621), .Y(n9980) );
  MUX2X1 U9674 ( .B(n9984), .A(n9985), .S(read2_addr[1]), .Y(n9983) );
  MUX2X1 U9675 ( .B(n9987), .A(n9988), .S(n10621), .Y(n9986) );
  MUX2X1 U9676 ( .B(n9990), .A(n9991), .S(n10621), .Y(n9989) );
  MUX2X1 U9677 ( .B(n9993), .A(n9994), .S(n10621), .Y(n9992) );
  MUX2X1 U9678 ( .B(n9996), .A(n9997), .S(n10621), .Y(n9995) );
  MUX2X1 U9679 ( .B(n9999), .A(n10000), .S(n10565), .Y(n9998) );
  MUX2X1 U9680 ( .B(n10002), .A(n10003), .S(n10622), .Y(n10001) );
  MUX2X1 U9681 ( .B(n10005), .A(n10006), .S(n10622), .Y(n10004) );
  MUX2X1 U9682 ( .B(n10008), .A(n10009), .S(n10622), .Y(n10007) );
  MUX2X1 U9683 ( .B(n10011), .A(n10012), .S(n10622), .Y(n10010) );
  MUX2X1 U9684 ( .B(n10014), .A(n10015), .S(n10563), .Y(n10013) );
  MUX2X1 U9685 ( .B(n10017), .A(n10018), .S(n10622), .Y(n10016) );
  MUX2X1 U9686 ( .B(n10020), .A(n10021), .S(n10622), .Y(n10019) );
  MUX2X1 U9687 ( .B(n10023), .A(n10024), .S(n10622), .Y(n10022) );
  MUX2X1 U9688 ( .B(n10026), .A(n10027), .S(n10622), .Y(n10025) );
  MUX2X1 U9689 ( .B(n10029), .A(n10030), .S(n10564), .Y(n10028) );
  MUX2X1 U9690 ( .B(n10032), .A(n10033), .S(n10622), .Y(n10031) );
  MUX2X1 U9691 ( .B(n10035), .A(n10036), .S(n10622), .Y(n10034) );
  MUX2X1 U9692 ( .B(n10038), .A(n10039), .S(n10622), .Y(n10037) );
  MUX2X1 U9693 ( .B(n10041), .A(n10042), .S(n10622), .Y(n10040) );
  MUX2X1 U9694 ( .B(n10044), .A(n10045), .S(n10564), .Y(n10043) );
  MUX2X1 U9695 ( .B(n10047), .A(n10048), .S(n10623), .Y(n10046) );
  MUX2X1 U9696 ( .B(n10050), .A(n10051), .S(n10623), .Y(n10049) );
  MUX2X1 U9697 ( .B(n10053), .A(n10054), .S(n10623), .Y(n10052) );
  MUX2X1 U9698 ( .B(n10056), .A(n10057), .S(n10623), .Y(n10055) );
  MUX2X1 U9699 ( .B(n10059), .A(n10060), .S(n10563), .Y(n10058) );
  MUX2X1 U9700 ( .B(n10062), .A(n10063), .S(n10623), .Y(n10061) );
  MUX2X1 U9701 ( .B(n10065), .A(n10066), .S(n10623), .Y(n10064) );
  MUX2X1 U9702 ( .B(n10068), .A(n10069), .S(n10623), .Y(n10067) );
  MUX2X1 U9703 ( .B(n10071), .A(n10072), .S(n10623), .Y(n10070) );
  MUX2X1 U9704 ( .B(n10074), .A(n10075), .S(read2_addr[1]), .Y(n10073) );
  MUX2X1 U9705 ( .B(n10077), .A(n10078), .S(n10623), .Y(n10076) );
  MUX2X1 U9706 ( .B(n10080), .A(n10081), .S(n10623), .Y(n10079) );
  MUX2X1 U9707 ( .B(n10083), .A(n10084), .S(n10623), .Y(n10082) );
  MUX2X1 U9708 ( .B(n10086), .A(n10087), .S(n10623), .Y(n10085) );
  MUX2X1 U9709 ( .B(n10089), .A(n10090), .S(n10563), .Y(n10088) );
  MUX2X1 U9710 ( .B(n10092), .A(n10093), .S(n10624), .Y(n10091) );
  MUX2X1 U9711 ( .B(n10095), .A(n10096), .S(n10624), .Y(n10094) );
  MUX2X1 U9712 ( .B(n10098), .A(n10099), .S(n10624), .Y(n10097) );
  MUX2X1 U9713 ( .B(n10101), .A(n10102), .S(n10624), .Y(n10100) );
  MUX2X1 U9714 ( .B(n10104), .A(n10105), .S(n10565), .Y(n10103) );
  MUX2X1 U9715 ( .B(n10107), .A(n10108), .S(n10624), .Y(n10106) );
  MUX2X1 U9716 ( .B(n10110), .A(n10111), .S(n10624), .Y(n10109) );
  MUX2X1 U9717 ( .B(n10113), .A(n10114), .S(n10624), .Y(n10112) );
  MUX2X1 U9718 ( .B(n10116), .A(n10117), .S(n10624), .Y(n10115) );
  MUX2X1 U9719 ( .B(n10119), .A(n10120), .S(read2_addr[1]), .Y(n10118) );
  MUX2X1 U9720 ( .B(n10122), .A(n10123), .S(n10624), .Y(n10121) );
  MUX2X1 U9721 ( .B(n10125), .A(n10126), .S(n10624), .Y(n10124) );
  MUX2X1 U9722 ( .B(n10128), .A(n10129), .S(n10624), .Y(n10127) );
  MUX2X1 U9723 ( .B(n10131), .A(n10132), .S(n10624), .Y(n10130) );
  MUX2X1 U9724 ( .B(n10134), .A(n10135), .S(n10564), .Y(n10133) );
  MUX2X1 U9725 ( .B(n10137), .A(n10138), .S(n10625), .Y(n10136) );
  MUX2X1 U9726 ( .B(n10140), .A(n10141), .S(n10625), .Y(n10139) );
  MUX2X1 U9727 ( .B(n10143), .A(n10144), .S(n10625), .Y(n10142) );
  MUX2X1 U9728 ( .B(n10146), .A(n10147), .S(n10625), .Y(n10145) );
  MUX2X1 U9729 ( .B(n10149), .A(n10150), .S(read2_addr[1]), .Y(n10148) );
  MUX2X1 U9730 ( .B(n10152), .A(n10153), .S(n10625), .Y(n10151) );
  MUX2X1 U9731 ( .B(n10155), .A(n10156), .S(n10625), .Y(n10154) );
  MUX2X1 U9732 ( .B(n10158), .A(n10159), .S(n10625), .Y(n10157) );
  MUX2X1 U9733 ( .B(n10161), .A(n10162), .S(n10625), .Y(n10160) );
  MUX2X1 U9734 ( .B(n10164), .A(n10165), .S(n10564), .Y(n10163) );
  MUX2X1 U9735 ( .B(n10167), .A(n10168), .S(n10625), .Y(n10166) );
  MUX2X1 U9736 ( .B(n10170), .A(n10171), .S(n10625), .Y(n10169) );
  MUX2X1 U9737 ( .B(n10173), .A(n10174), .S(n10625), .Y(n10172) );
  MUX2X1 U9738 ( .B(n10176), .A(n10177), .S(n10625), .Y(n10175) );
  MUX2X1 U9739 ( .B(n10179), .A(n10180), .S(n10565), .Y(n10178) );
  MUX2X1 U9740 ( .B(n10182), .A(n10183), .S(n10626), .Y(n10181) );
  MUX2X1 U9741 ( .B(n10185), .A(n10186), .S(n10626), .Y(n10184) );
  MUX2X1 U9742 ( .B(n10188), .A(n10189), .S(n10626), .Y(n10187) );
  MUX2X1 U9743 ( .B(n10191), .A(n10192), .S(n10626), .Y(n10190) );
  MUX2X1 U9744 ( .B(n10194), .A(n10195), .S(n10564), .Y(n10193) );
  MUX2X1 U9745 ( .B(n10197), .A(n10198), .S(n10626), .Y(n10196) );
  MUX2X1 U9746 ( .B(n10200), .A(n10201), .S(n10626), .Y(n10199) );
  MUX2X1 U9747 ( .B(n10203), .A(n10204), .S(n10626), .Y(n10202) );
  MUX2X1 U9748 ( .B(n10206), .A(n10207), .S(n10626), .Y(n10205) );
  MUX2X1 U9749 ( .B(n10209), .A(n10210), .S(n10565), .Y(n10208) );
  MUX2X1 U9750 ( .B(n10212), .A(n10213), .S(n10626), .Y(n10211) );
  MUX2X1 U9751 ( .B(n10215), .A(n10216), .S(n10626), .Y(n10214) );
  MUX2X1 U9752 ( .B(n10218), .A(n10219), .S(n10626), .Y(n10217) );
  MUX2X1 U9753 ( .B(n10221), .A(n10222), .S(n10626), .Y(n10220) );
  MUX2X1 U9754 ( .B(n10224), .A(n10225), .S(read2_addr[1]), .Y(n10223) );
  MUX2X1 U9755 ( .B(n10227), .A(n10228), .S(n10627), .Y(n10226) );
  MUX2X1 U9756 ( .B(n10230), .A(n10231), .S(n10627), .Y(n10229) );
  MUX2X1 U9757 ( .B(n10233), .A(n10234), .S(n10627), .Y(n10232) );
  MUX2X1 U9758 ( .B(n10236), .A(n10237), .S(n10627), .Y(n10235) );
  MUX2X1 U9759 ( .B(n10239), .A(n10240), .S(n10565), .Y(n10238) );
  MUX2X1 U9760 ( .B(n10242), .A(n10243), .S(n10627), .Y(n10241) );
  MUX2X1 U9761 ( .B(n10245), .A(n10246), .S(n10627), .Y(n10244) );
  MUX2X1 U9762 ( .B(n10248), .A(n10249), .S(n10627), .Y(n10247) );
  MUX2X1 U9763 ( .B(n10251), .A(n10252), .S(n10627), .Y(n10250) );
  MUX2X1 U9764 ( .B(n10254), .A(n10255), .S(n10565), .Y(n10253) );
  MUX2X1 U9765 ( .B(n10257), .A(n10258), .S(n10627), .Y(n10256) );
  MUX2X1 U9766 ( .B(n10260), .A(n10261), .S(n10627), .Y(n10259) );
  MUX2X1 U9767 ( .B(n10263), .A(n10264), .S(n10627), .Y(n10262) );
  MUX2X1 U9768 ( .B(n10266), .A(n10267), .S(n10627), .Y(n10265) );
  MUX2X1 U9769 ( .B(n10269), .A(n10270), .S(n10564), .Y(n10268) );
  MUX2X1 U9770 ( .B(n10272), .A(n10273), .S(n10628), .Y(n10271) );
  MUX2X1 U9771 ( .B(n10275), .A(n10276), .S(n10628), .Y(n10274) );
  MUX2X1 U9772 ( .B(n10278), .A(n10279), .S(n10628), .Y(n10277) );
  MUX2X1 U9773 ( .B(n10281), .A(n10282), .S(n10628), .Y(n10280) );
  MUX2X1 U9774 ( .B(n10284), .A(n10285), .S(n10564), .Y(n10283) );
  MUX2X1 U9775 ( .B(n10287), .A(n10288), .S(n10628), .Y(n10286) );
  MUX2X1 U9776 ( .B(n10290), .A(n10291), .S(n10628), .Y(n10289) );
  MUX2X1 U9777 ( .B(n10293), .A(n10294), .S(n10628), .Y(n10292) );
  MUX2X1 U9778 ( .B(n10296), .A(n10297), .S(n10628), .Y(n10295) );
  MUX2X1 U9779 ( .B(n10299), .A(n10300), .S(n10563), .Y(n10298) );
  MUX2X1 U9780 ( .B(n10302), .A(n10303), .S(n10628), .Y(n10301) );
  MUX2X1 U9781 ( .B(n10305), .A(n10306), .S(n10628), .Y(n10304) );
  MUX2X1 U9782 ( .B(n10308), .A(n10309), .S(n10628), .Y(n10307) );
  MUX2X1 U9783 ( .B(n10311), .A(n10312), .S(n10628), .Y(n10310) );
  MUX2X1 U9784 ( .B(n10314), .A(n10315), .S(n10563), .Y(n10313) );
  MUX2X1 U9785 ( .B(n10317), .A(n10318), .S(n10629), .Y(n10316) );
  MUX2X1 U9786 ( .B(n10320), .A(n10321), .S(n10629), .Y(n10319) );
  MUX2X1 U9787 ( .B(n10323), .A(n10324), .S(n10629), .Y(n10322) );
  MUX2X1 U9788 ( .B(n10326), .A(n10327), .S(n10629), .Y(n10325) );
  MUX2X1 U9789 ( .B(n10329), .A(n10330), .S(read2_addr[1]), .Y(n10328) );
  MUX2X1 U9790 ( .B(n10332), .A(n10333), .S(n10629), .Y(n10331) );
  MUX2X1 U9791 ( .B(n10335), .A(n10336), .S(n10629), .Y(n10334) );
  MUX2X1 U9792 ( .B(n10338), .A(n10339), .S(n10629), .Y(n10337) );
  MUX2X1 U9793 ( .B(n10341), .A(n10342), .S(n10629), .Y(n10340) );
  MUX2X1 U9794 ( .B(n10344), .A(n10345), .S(read2_addr[1]), .Y(n10343) );
  MUX2X1 U9795 ( .B(n10347), .A(n10348), .S(n10629), .Y(n10346) );
  MUX2X1 U9796 ( .B(n10350), .A(n10351), .S(n10629), .Y(n10349) );
  MUX2X1 U9797 ( .B(n10353), .A(n10354), .S(n10629), .Y(n10352) );
  MUX2X1 U9798 ( .B(n10356), .A(n10357), .S(n10629), .Y(n10355) );
  MUX2X1 U9799 ( .B(n10359), .A(n10360), .S(read2_addr[1]), .Y(n10358) );
  MUX2X1 U9800 ( .B(n10362), .A(n10363), .S(n10630), .Y(n10361) );
  MUX2X1 U9801 ( .B(n10365), .A(n10366), .S(n10630), .Y(n10364) );
  MUX2X1 U9802 ( .B(n10368), .A(n10369), .S(n10630), .Y(n10367) );
  MUX2X1 U9803 ( .B(n10371), .A(n10372), .S(n10630), .Y(n10370) );
  MUX2X1 U9804 ( .B(n10374), .A(n10375), .S(read2_addr[1]), .Y(n10373) );
  MUX2X1 U9805 ( .B(n10377), .A(n10378), .S(n10630), .Y(n10376) );
  MUX2X1 U9806 ( .B(n10380), .A(n10381), .S(n10630), .Y(n10379) );
  MUX2X1 U9807 ( .B(n10383), .A(n10384), .S(n10630), .Y(n10382) );
  MUX2X1 U9808 ( .B(n10386), .A(n10387), .S(n10630), .Y(n10385) );
  MUX2X1 U9809 ( .B(n10389), .A(n10390), .S(n10565), .Y(n10388) );
  MUX2X1 U9810 ( .B(n10392), .A(n10393), .S(n10630), .Y(n10391) );
  MUX2X1 U9811 ( .B(n10395), .A(n10396), .S(n10630), .Y(n10394) );
  MUX2X1 U9812 ( .B(n10398), .A(n10399), .S(n10630), .Y(n10397) );
  MUX2X1 U9813 ( .B(n10401), .A(n10402), .S(n10630), .Y(n10400) );
  MUX2X1 U9814 ( .B(n10404), .A(n10405), .S(n10565), .Y(n10403) );
  MUX2X1 U9815 ( .B(n10407), .A(n10408), .S(n10631), .Y(n10406) );
  MUX2X1 U9816 ( .B(n10410), .A(n10411), .S(n10631), .Y(n10409) );
  MUX2X1 U9817 ( .B(n10413), .A(n10414), .S(n10631), .Y(n10412) );
  MUX2X1 U9818 ( .B(n10416), .A(n10417), .S(n10631), .Y(n10415) );
  MUX2X1 U9819 ( .B(n10419), .A(n10420), .S(n10565), .Y(n10418) );
  MUX2X1 U9820 ( .B(n10422), .A(n10423), .S(n10631), .Y(n10421) );
  MUX2X1 U9821 ( .B(n10425), .A(n10426), .S(n10631), .Y(n10424) );
  MUX2X1 U9822 ( .B(n10428), .A(n10429), .S(n10631), .Y(n10427) );
  MUX2X1 U9823 ( .B(n10431), .A(n10432), .S(n10631), .Y(n10430) );
  MUX2X1 U9824 ( .B(n10434), .A(n10435), .S(n10564), .Y(n10433) );
  MUX2X1 U9825 ( .B(n10437), .A(n10438), .S(n10631), .Y(n10436) );
  MUX2X1 U9826 ( .B(n10440), .A(n10441), .S(n10631), .Y(n10439) );
  MUX2X1 U9827 ( .B(n10443), .A(n10444), .S(n10631), .Y(n10442) );
  MUX2X1 U9828 ( .B(n10446), .A(n10447), .S(n10631), .Y(n10445) );
  MUX2X1 U9829 ( .B(n10449), .A(n10450), .S(n10563), .Y(n10448) );
  MUX2X1 U9830 ( .B(n10452), .A(n10453), .S(n10632), .Y(n10451) );
  MUX2X1 U9831 ( .B(n10455), .A(n10456), .S(n10632), .Y(n10454) );
  MUX2X1 U9832 ( .B(n10458), .A(n10459), .S(n10632), .Y(n10457) );
  MUX2X1 U9833 ( .B(n10461), .A(n10462), .S(n10632), .Y(n10460) );
  MUX2X1 U9834 ( .B(n10464), .A(n10465), .S(read2_addr[1]), .Y(n10463) );
  MUX2X1 U9835 ( .B(n10467), .A(n10468), .S(n10632), .Y(n10466) );
  MUX2X1 U9836 ( .B(n10470), .A(n10471), .S(n10632), .Y(n10469) );
  MUX2X1 U9837 ( .B(n10473), .A(n10474), .S(n10632), .Y(n10472) );
  MUX2X1 U9838 ( .B(n10476), .A(n10477), .S(n10632), .Y(n10475) );
  MUX2X1 U9839 ( .B(n10479), .A(n10480), .S(n10565), .Y(n10478) );
  MUX2X1 U9840 ( .B(n10482), .A(n10483), .S(n10632), .Y(n10481) );
  MUX2X1 U9841 ( .B(n10485), .A(n10486), .S(n10632), .Y(n10484) );
  MUX2X1 U9842 ( .B(n10488), .A(n10489), .S(n10632), .Y(n10487) );
  MUX2X1 U9843 ( .B(n10491), .A(n10492), .S(n10632), .Y(n10490) );
  MUX2X1 U9844 ( .B(n10494), .A(n10495), .S(n10563), .Y(n10493) );
  MUX2X1 U9845 ( .B(ram[64]), .A(ram[0]), .S(n10657), .Y(n8578) );
  MUX2X1 U9846 ( .B(ram[192]), .A(ram[128]), .S(n10657), .Y(n8577) );
  MUX2X1 U9847 ( .B(ram[320]), .A(ram[256]), .S(n10657), .Y(n8581) );
  MUX2X1 U9848 ( .B(ram[448]), .A(ram[384]), .S(n10657), .Y(n8580) );
  MUX2X1 U9849 ( .B(n8579), .A(n8576), .S(n10572), .Y(n8590) );
  MUX2X1 U9850 ( .B(ram[576]), .A(ram[512]), .S(n10658), .Y(n8584) );
  MUX2X1 U9851 ( .B(ram[704]), .A(ram[640]), .S(n10658), .Y(n8583) );
  MUX2X1 U9852 ( .B(ram[832]), .A(ram[768]), .S(n10658), .Y(n8587) );
  MUX2X1 U9853 ( .B(ram[960]), .A(ram[896]), .S(n10658), .Y(n8586) );
  MUX2X1 U9854 ( .B(n8585), .A(n8582), .S(n10571), .Y(n8589) );
  MUX2X1 U9855 ( .B(ram[1088]), .A(ram[1024]), .S(n10658), .Y(n8593) );
  MUX2X1 U9856 ( .B(ram[1216]), .A(ram[1152]), .S(n10658), .Y(n8592) );
  MUX2X1 U9857 ( .B(ram[1344]), .A(ram[1280]), .S(n10658), .Y(n8596) );
  MUX2X1 U9858 ( .B(ram[1472]), .A(ram[1408]), .S(n10658), .Y(n8595) );
  MUX2X1 U9859 ( .B(n8594), .A(n8591), .S(n10574), .Y(n8605) );
  MUX2X1 U9860 ( .B(ram[1600]), .A(ram[1536]), .S(n10658), .Y(n8599) );
  MUX2X1 U9861 ( .B(ram[1728]), .A(ram[1664]), .S(n10658), .Y(n8598) );
  MUX2X1 U9862 ( .B(ram[1856]), .A(ram[1792]), .S(n10658), .Y(n8602) );
  MUX2X1 U9863 ( .B(ram[1984]), .A(ram[1920]), .S(n10658), .Y(n8601) );
  MUX2X1 U9864 ( .B(n8600), .A(n8597), .S(n10582), .Y(n8604) );
  MUX2X1 U9865 ( .B(n8603), .A(n8588), .S(n10562), .Y(n10496) );
  MUX2X1 U9866 ( .B(ram[65]), .A(ram[1]), .S(n10659), .Y(n8608) );
  MUX2X1 U9867 ( .B(ram[193]), .A(ram[129]), .S(n10659), .Y(n8607) );
  MUX2X1 U9868 ( .B(ram[321]), .A(ram[257]), .S(n10659), .Y(n8611) );
  MUX2X1 U9869 ( .B(ram[449]), .A(ram[385]), .S(n10659), .Y(n8610) );
  MUX2X1 U9870 ( .B(n8609), .A(n8606), .S(n10568), .Y(n8620) );
  MUX2X1 U9871 ( .B(ram[577]), .A(ram[513]), .S(n10659), .Y(n8614) );
  MUX2X1 U9872 ( .B(ram[705]), .A(ram[641]), .S(n10659), .Y(n8613) );
  MUX2X1 U9873 ( .B(ram[833]), .A(ram[769]), .S(n10659), .Y(n8617) );
  MUX2X1 U9874 ( .B(ram[961]), .A(ram[897]), .S(n10659), .Y(n8616) );
  MUX2X1 U9875 ( .B(n8615), .A(n8612), .S(n10568), .Y(n8619) );
  MUX2X1 U9876 ( .B(ram[1089]), .A(ram[1025]), .S(n10659), .Y(n8623) );
  MUX2X1 U9877 ( .B(ram[1217]), .A(ram[1153]), .S(n10659), .Y(n8622) );
  MUX2X1 U9878 ( .B(ram[1345]), .A(ram[1281]), .S(n10659), .Y(n8626) );
  MUX2X1 U9879 ( .B(ram[1473]), .A(ram[1409]), .S(n10659), .Y(n8625) );
  MUX2X1 U9880 ( .B(n8624), .A(n8621), .S(n10568), .Y(n8635) );
  MUX2X1 U9881 ( .B(ram[1601]), .A(ram[1537]), .S(n10660), .Y(n8629) );
  MUX2X1 U9882 ( .B(ram[1729]), .A(ram[1665]), .S(n10660), .Y(n8628) );
  MUX2X1 U9883 ( .B(ram[1857]), .A(ram[1793]), .S(n10660), .Y(n8632) );
  MUX2X1 U9884 ( .B(ram[1985]), .A(ram[1921]), .S(n10660), .Y(n8631) );
  MUX2X1 U9885 ( .B(n8630), .A(n8627), .S(n10568), .Y(n8634) );
  MUX2X1 U9886 ( .B(n8633), .A(n8618), .S(n10562), .Y(n10497) );
  MUX2X1 U9887 ( .B(ram[66]), .A(ram[2]), .S(n10660), .Y(n8638) );
  MUX2X1 U9888 ( .B(ram[194]), .A(ram[130]), .S(n10660), .Y(n8637) );
  MUX2X1 U9889 ( .B(ram[322]), .A(ram[258]), .S(n10660), .Y(n8641) );
  MUX2X1 U9890 ( .B(ram[450]), .A(ram[386]), .S(n10660), .Y(n8640) );
  MUX2X1 U9891 ( .B(n8639), .A(n8636), .S(n10568), .Y(n8650) );
  MUX2X1 U9892 ( .B(ram[578]), .A(ram[514]), .S(n10660), .Y(n8644) );
  MUX2X1 U9893 ( .B(ram[706]), .A(ram[642]), .S(n10660), .Y(n8643) );
  MUX2X1 U9894 ( .B(ram[834]), .A(ram[770]), .S(n10660), .Y(n8647) );
  MUX2X1 U9895 ( .B(ram[962]), .A(ram[898]), .S(n10660), .Y(n8646) );
  MUX2X1 U9896 ( .B(n8645), .A(n8642), .S(n10568), .Y(n8649) );
  MUX2X1 U9897 ( .B(ram[1090]), .A(ram[1026]), .S(n10661), .Y(n8653) );
  MUX2X1 U9898 ( .B(ram[1218]), .A(ram[1154]), .S(n10661), .Y(n8652) );
  MUX2X1 U9899 ( .B(ram[1346]), .A(ram[1282]), .S(n10661), .Y(n8656) );
  MUX2X1 U9900 ( .B(ram[1474]), .A(ram[1410]), .S(n10661), .Y(n8655) );
  MUX2X1 U9901 ( .B(n8654), .A(n8651), .S(n10568), .Y(n8665) );
  MUX2X1 U9902 ( .B(ram[1602]), .A(ram[1538]), .S(n10661), .Y(n8659) );
  MUX2X1 U9903 ( .B(ram[1730]), .A(ram[1666]), .S(n10661), .Y(n8658) );
  MUX2X1 U9904 ( .B(ram[1858]), .A(ram[1794]), .S(n10661), .Y(n8662) );
  MUX2X1 U9905 ( .B(ram[1986]), .A(ram[1922]), .S(n10661), .Y(n8661) );
  MUX2X1 U9906 ( .B(n8660), .A(n8657), .S(n10568), .Y(n8664) );
  MUX2X1 U9907 ( .B(n8663), .A(n8648), .S(n10562), .Y(n10498) );
  MUX2X1 U9908 ( .B(ram[67]), .A(ram[3]), .S(n10661), .Y(n8668) );
  MUX2X1 U9909 ( .B(ram[195]), .A(ram[131]), .S(n10661), .Y(n8667) );
  MUX2X1 U9910 ( .B(ram[323]), .A(ram[259]), .S(n10661), .Y(n8671) );
  MUX2X1 U9911 ( .B(ram[451]), .A(ram[387]), .S(n10661), .Y(n8670) );
  MUX2X1 U9912 ( .B(n8669), .A(n8666), .S(n10568), .Y(n8680) );
  MUX2X1 U9913 ( .B(ram[579]), .A(ram[515]), .S(n10662), .Y(n8674) );
  MUX2X1 U9914 ( .B(ram[707]), .A(ram[643]), .S(n10662), .Y(n8673) );
  MUX2X1 U9915 ( .B(ram[835]), .A(ram[771]), .S(n10662), .Y(n8677) );
  MUX2X1 U9916 ( .B(ram[963]), .A(ram[899]), .S(n10662), .Y(n8676) );
  MUX2X1 U9917 ( .B(n8675), .A(n8672), .S(n10568), .Y(n8679) );
  MUX2X1 U9918 ( .B(ram[1091]), .A(ram[1027]), .S(n10662), .Y(n8683) );
  MUX2X1 U9919 ( .B(ram[1219]), .A(ram[1155]), .S(n10662), .Y(n8682) );
  MUX2X1 U9920 ( .B(ram[1347]), .A(ram[1283]), .S(n10662), .Y(n8686) );
  MUX2X1 U9921 ( .B(ram[1475]), .A(ram[1411]), .S(n10662), .Y(n8685) );
  MUX2X1 U9922 ( .B(n8684), .A(n8681), .S(n10568), .Y(n8695) );
  MUX2X1 U9923 ( .B(ram[1603]), .A(ram[1539]), .S(n10662), .Y(n8689) );
  MUX2X1 U9924 ( .B(ram[1731]), .A(ram[1667]), .S(n10662), .Y(n8688) );
  MUX2X1 U9925 ( .B(ram[1859]), .A(ram[1795]), .S(n10662), .Y(n8692) );
  MUX2X1 U9926 ( .B(ram[1987]), .A(ram[1923]), .S(n10662), .Y(n8691) );
  MUX2X1 U9927 ( .B(n8690), .A(n8687), .S(n10568), .Y(n8694) );
  MUX2X1 U9928 ( .B(n8693), .A(n8678), .S(n10562), .Y(n10499) );
  MUX2X1 U9929 ( .B(ram[68]), .A(ram[4]), .S(n10663), .Y(n8698) );
  MUX2X1 U9930 ( .B(ram[196]), .A(ram[132]), .S(n10663), .Y(n8697) );
  MUX2X1 U9931 ( .B(ram[324]), .A(ram[260]), .S(n10663), .Y(n8701) );
  MUX2X1 U9932 ( .B(ram[452]), .A(ram[388]), .S(n10663), .Y(n8700) );
  MUX2X1 U9933 ( .B(n8699), .A(n8696), .S(n10569), .Y(n8710) );
  MUX2X1 U9934 ( .B(ram[580]), .A(ram[516]), .S(n10663), .Y(n8704) );
  MUX2X1 U9935 ( .B(ram[708]), .A(ram[644]), .S(n10663), .Y(n8703) );
  MUX2X1 U9936 ( .B(ram[836]), .A(ram[772]), .S(n10663), .Y(n8707) );
  MUX2X1 U9937 ( .B(ram[964]), .A(ram[900]), .S(n10663), .Y(n8706) );
  MUX2X1 U9938 ( .B(n8705), .A(n8702), .S(n10569), .Y(n8709) );
  MUX2X1 U9939 ( .B(ram[1092]), .A(ram[1028]), .S(n10663), .Y(n8713) );
  MUX2X1 U9940 ( .B(ram[1220]), .A(ram[1156]), .S(n10663), .Y(n8712) );
  MUX2X1 U9941 ( .B(ram[1348]), .A(ram[1284]), .S(n10663), .Y(n8716) );
  MUX2X1 U9942 ( .B(ram[1476]), .A(ram[1412]), .S(n10663), .Y(n8715) );
  MUX2X1 U9943 ( .B(n8714), .A(n8711), .S(n10569), .Y(n8725) );
  MUX2X1 U9944 ( .B(ram[1604]), .A(ram[1540]), .S(n10664), .Y(n8719) );
  MUX2X1 U9945 ( .B(ram[1732]), .A(ram[1668]), .S(n10664), .Y(n8718) );
  MUX2X1 U9946 ( .B(ram[1860]), .A(ram[1796]), .S(n10664), .Y(n8722) );
  MUX2X1 U9947 ( .B(ram[1988]), .A(ram[1924]), .S(n10664), .Y(n8721) );
  MUX2X1 U9948 ( .B(n8720), .A(n8717), .S(n10569), .Y(n8724) );
  MUX2X1 U9949 ( .B(n8723), .A(n8708), .S(n10562), .Y(n10500) );
  MUX2X1 U9950 ( .B(ram[69]), .A(ram[5]), .S(n10664), .Y(n8728) );
  MUX2X1 U9951 ( .B(ram[197]), .A(ram[133]), .S(n10664), .Y(n8727) );
  MUX2X1 U9952 ( .B(ram[325]), .A(ram[261]), .S(n10664), .Y(n8731) );
  MUX2X1 U9953 ( .B(ram[453]), .A(ram[389]), .S(n10664), .Y(n8730) );
  MUX2X1 U9954 ( .B(n8729), .A(n8726), .S(n10569), .Y(n8740) );
  MUX2X1 U9955 ( .B(ram[581]), .A(ram[517]), .S(n10664), .Y(n8734) );
  MUX2X1 U9956 ( .B(ram[709]), .A(ram[645]), .S(n10664), .Y(n8733) );
  MUX2X1 U9957 ( .B(ram[837]), .A(ram[773]), .S(n10664), .Y(n8737) );
  MUX2X1 U9958 ( .B(ram[965]), .A(ram[901]), .S(n10664), .Y(n8736) );
  MUX2X1 U9959 ( .B(n8735), .A(n8732), .S(n10569), .Y(n8739) );
  MUX2X1 U9960 ( .B(ram[1093]), .A(ram[1029]), .S(n10665), .Y(n8743) );
  MUX2X1 U9961 ( .B(ram[1221]), .A(ram[1157]), .S(n10665), .Y(n8742) );
  MUX2X1 U9962 ( .B(ram[1349]), .A(ram[1285]), .S(n10665), .Y(n8746) );
  MUX2X1 U9963 ( .B(ram[1477]), .A(ram[1413]), .S(n10665), .Y(n8745) );
  MUX2X1 U9964 ( .B(n8744), .A(n8741), .S(n10569), .Y(n8755) );
  MUX2X1 U9965 ( .B(ram[1605]), .A(ram[1541]), .S(n10665), .Y(n8749) );
  MUX2X1 U9966 ( .B(ram[1733]), .A(ram[1669]), .S(n10665), .Y(n8748) );
  MUX2X1 U9967 ( .B(ram[1861]), .A(ram[1797]), .S(n10665), .Y(n8752) );
  MUX2X1 U9968 ( .B(ram[1989]), .A(ram[1925]), .S(n10665), .Y(n8751) );
  MUX2X1 U9969 ( .B(n8750), .A(n8747), .S(n10569), .Y(n8754) );
  MUX2X1 U9970 ( .B(n8753), .A(n8738), .S(n10562), .Y(n10501) );
  MUX2X1 U9971 ( .B(ram[70]), .A(ram[6]), .S(n10665), .Y(n8758) );
  MUX2X1 U9972 ( .B(ram[198]), .A(ram[134]), .S(n10665), .Y(n8757) );
  MUX2X1 U9973 ( .B(ram[326]), .A(ram[262]), .S(n10665), .Y(n8761) );
  MUX2X1 U9974 ( .B(ram[454]), .A(ram[390]), .S(n10665), .Y(n8760) );
  MUX2X1 U9975 ( .B(n8759), .A(n8756), .S(n10569), .Y(n8770) );
  MUX2X1 U9976 ( .B(ram[582]), .A(ram[518]), .S(n10666), .Y(n8764) );
  MUX2X1 U9977 ( .B(ram[710]), .A(ram[646]), .S(n10666), .Y(n8763) );
  MUX2X1 U9978 ( .B(ram[838]), .A(ram[774]), .S(n10666), .Y(n8767) );
  MUX2X1 U9979 ( .B(ram[966]), .A(ram[902]), .S(n10666), .Y(n8766) );
  MUX2X1 U9980 ( .B(n8765), .A(n8762), .S(n10569), .Y(n8769) );
  MUX2X1 U9981 ( .B(ram[1094]), .A(ram[1030]), .S(n10666), .Y(n8773) );
  MUX2X1 U9982 ( .B(ram[1222]), .A(ram[1158]), .S(n10666), .Y(n8772) );
  MUX2X1 U9983 ( .B(ram[1350]), .A(ram[1286]), .S(n10666), .Y(n8776) );
  MUX2X1 U9984 ( .B(ram[1478]), .A(ram[1414]), .S(n10666), .Y(n8775) );
  MUX2X1 U9985 ( .B(n8774), .A(n8771), .S(n10569), .Y(n8785) );
  MUX2X1 U9986 ( .B(ram[1606]), .A(ram[1542]), .S(n10666), .Y(n8779) );
  MUX2X1 U9987 ( .B(ram[1734]), .A(ram[1670]), .S(n10666), .Y(n8778) );
  MUX2X1 U9988 ( .B(ram[1862]), .A(ram[1798]), .S(n10666), .Y(n8782) );
  MUX2X1 U9989 ( .B(ram[1990]), .A(ram[1926]), .S(n10666), .Y(n8781) );
  MUX2X1 U9990 ( .B(n8780), .A(n8777), .S(n10569), .Y(n8784) );
  MUX2X1 U9991 ( .B(n8783), .A(n8768), .S(n10562), .Y(n10502) );
  MUX2X1 U9992 ( .B(ram[71]), .A(ram[7]), .S(n10667), .Y(n8788) );
  MUX2X1 U9993 ( .B(ram[199]), .A(ram[135]), .S(n10667), .Y(n8787) );
  MUX2X1 U9994 ( .B(ram[327]), .A(ram[263]), .S(n10667), .Y(n8791) );
  MUX2X1 U9995 ( .B(ram[455]), .A(ram[391]), .S(n10667), .Y(n8790) );
  MUX2X1 U9996 ( .B(n8789), .A(n8786), .S(n10570), .Y(n8800) );
  MUX2X1 U9997 ( .B(ram[583]), .A(ram[519]), .S(n10667), .Y(n8794) );
  MUX2X1 U9998 ( .B(ram[711]), .A(ram[647]), .S(n10667), .Y(n8793) );
  MUX2X1 U9999 ( .B(ram[839]), .A(ram[775]), .S(n10667), .Y(n8797) );
  MUX2X1 U10000 ( .B(ram[967]), .A(ram[903]), .S(n10667), .Y(n8796) );
  MUX2X1 U10001 ( .B(n8795), .A(n8792), .S(n10570), .Y(n8799) );
  MUX2X1 U10002 ( .B(ram[1095]), .A(ram[1031]), .S(n10667), .Y(n8803) );
  MUX2X1 U10003 ( .B(ram[1223]), .A(ram[1159]), .S(n10667), .Y(n8802) );
  MUX2X1 U10004 ( .B(ram[1351]), .A(ram[1287]), .S(n10667), .Y(n8806) );
  MUX2X1 U10005 ( .B(ram[1479]), .A(ram[1415]), .S(n10667), .Y(n8805) );
  MUX2X1 U10006 ( .B(n8804), .A(n8801), .S(n10570), .Y(n8815) );
  MUX2X1 U10007 ( .B(ram[1607]), .A(ram[1543]), .S(n10668), .Y(n8809) );
  MUX2X1 U10008 ( .B(ram[1735]), .A(ram[1671]), .S(n10668), .Y(n8808) );
  MUX2X1 U10009 ( .B(ram[1863]), .A(ram[1799]), .S(n10668), .Y(n8812) );
  MUX2X1 U10010 ( .B(ram[1991]), .A(ram[1927]), .S(n10668), .Y(n8811) );
  MUX2X1 U10011 ( .B(n8810), .A(n8807), .S(n10570), .Y(n8814) );
  MUX2X1 U10012 ( .B(n8813), .A(n8798), .S(n10562), .Y(n10503) );
  MUX2X1 U10013 ( .B(ram[72]), .A(ram[8]), .S(n10668), .Y(n8818) );
  MUX2X1 U10014 ( .B(ram[200]), .A(ram[136]), .S(n10668), .Y(n8817) );
  MUX2X1 U10015 ( .B(ram[328]), .A(ram[264]), .S(n10668), .Y(n8821) );
  MUX2X1 U10016 ( .B(ram[456]), .A(ram[392]), .S(n10668), .Y(n8820) );
  MUX2X1 U10017 ( .B(n8819), .A(n8816), .S(n10570), .Y(n8830) );
  MUX2X1 U10018 ( .B(ram[584]), .A(ram[520]), .S(n10668), .Y(n8824) );
  MUX2X1 U10019 ( .B(ram[712]), .A(ram[648]), .S(n10668), .Y(n8823) );
  MUX2X1 U10020 ( .B(ram[840]), .A(ram[776]), .S(n10668), .Y(n8827) );
  MUX2X1 U10021 ( .B(ram[968]), .A(ram[904]), .S(n10668), .Y(n8826) );
  MUX2X1 U10022 ( .B(n8825), .A(n8822), .S(n10570), .Y(n8829) );
  MUX2X1 U10023 ( .B(ram[1096]), .A(ram[1032]), .S(n10669), .Y(n8833) );
  MUX2X1 U10024 ( .B(ram[1224]), .A(ram[1160]), .S(n10669), .Y(n8832) );
  MUX2X1 U10025 ( .B(ram[1352]), .A(ram[1288]), .S(n10669), .Y(n8836) );
  MUX2X1 U10026 ( .B(ram[1480]), .A(ram[1416]), .S(n10669), .Y(n8835) );
  MUX2X1 U10027 ( .B(n8834), .A(n8831), .S(n10570), .Y(n8845) );
  MUX2X1 U10028 ( .B(ram[1608]), .A(ram[1544]), .S(n10669), .Y(n8839) );
  MUX2X1 U10029 ( .B(ram[1736]), .A(ram[1672]), .S(n10669), .Y(n8838) );
  MUX2X1 U10030 ( .B(ram[1864]), .A(ram[1800]), .S(n10669), .Y(n8842) );
  MUX2X1 U10031 ( .B(ram[1992]), .A(ram[1928]), .S(n10669), .Y(n8841) );
  MUX2X1 U10032 ( .B(n8840), .A(n8837), .S(n10570), .Y(n8844) );
  MUX2X1 U10033 ( .B(n8843), .A(n8828), .S(n10562), .Y(n10504) );
  MUX2X1 U10034 ( .B(ram[73]), .A(ram[9]), .S(n10669), .Y(n8848) );
  MUX2X1 U10035 ( .B(ram[201]), .A(ram[137]), .S(n10669), .Y(n8847) );
  MUX2X1 U10036 ( .B(ram[329]), .A(ram[265]), .S(n10669), .Y(n8851) );
  MUX2X1 U10037 ( .B(ram[457]), .A(ram[393]), .S(n10669), .Y(n8850) );
  MUX2X1 U10038 ( .B(n8849), .A(n8846), .S(n10570), .Y(n8860) );
  MUX2X1 U10039 ( .B(ram[585]), .A(ram[521]), .S(n10670), .Y(n8854) );
  MUX2X1 U10040 ( .B(ram[713]), .A(ram[649]), .S(n10670), .Y(n8853) );
  MUX2X1 U10041 ( .B(ram[841]), .A(ram[777]), .S(n10670), .Y(n8857) );
  MUX2X1 U10042 ( .B(ram[969]), .A(ram[905]), .S(n10670), .Y(n8856) );
  MUX2X1 U10043 ( .B(n8855), .A(n8852), .S(n10570), .Y(n8859) );
  MUX2X1 U10044 ( .B(ram[1097]), .A(ram[1033]), .S(n10670), .Y(n8863) );
  MUX2X1 U10045 ( .B(ram[1225]), .A(ram[1161]), .S(n10670), .Y(n8862) );
  MUX2X1 U10046 ( .B(ram[1353]), .A(ram[1289]), .S(n10670), .Y(n8866) );
  MUX2X1 U10047 ( .B(ram[1481]), .A(ram[1417]), .S(n10670), .Y(n8865) );
  MUX2X1 U10048 ( .B(n8864), .A(n8861), .S(n10570), .Y(n8875) );
  MUX2X1 U10049 ( .B(ram[1609]), .A(ram[1545]), .S(n10670), .Y(n8869) );
  MUX2X1 U10050 ( .B(ram[1737]), .A(ram[1673]), .S(n10670), .Y(n8868) );
  MUX2X1 U10051 ( .B(ram[1865]), .A(ram[1801]), .S(n10670), .Y(n8872) );
  MUX2X1 U10052 ( .B(ram[1993]), .A(ram[1929]), .S(n10670), .Y(n8871) );
  MUX2X1 U10053 ( .B(n8870), .A(n8867), .S(n10570), .Y(n8874) );
  MUX2X1 U10054 ( .B(n8873), .A(n8858), .S(n10562), .Y(n10505) );
  MUX2X1 U10055 ( .B(ram[74]), .A(ram[10]), .S(n10671), .Y(n8878) );
  MUX2X1 U10056 ( .B(ram[202]), .A(ram[138]), .S(n10671), .Y(n8877) );
  MUX2X1 U10057 ( .B(ram[330]), .A(ram[266]), .S(n10671), .Y(n8881) );
  MUX2X1 U10058 ( .B(ram[458]), .A(ram[394]), .S(n10671), .Y(n8880) );
  MUX2X1 U10059 ( .B(n8879), .A(n8876), .S(n10571), .Y(n8890) );
  MUX2X1 U10060 ( .B(ram[586]), .A(ram[522]), .S(n10671), .Y(n8884) );
  MUX2X1 U10061 ( .B(ram[714]), .A(ram[650]), .S(n10671), .Y(n8883) );
  MUX2X1 U10062 ( .B(ram[842]), .A(ram[778]), .S(n10671), .Y(n8887) );
  MUX2X1 U10063 ( .B(ram[970]), .A(ram[906]), .S(n10671), .Y(n8886) );
  MUX2X1 U10064 ( .B(n8885), .A(n8882), .S(n10571), .Y(n8889) );
  MUX2X1 U10065 ( .B(ram[1098]), .A(ram[1034]), .S(n10671), .Y(n8893) );
  MUX2X1 U10066 ( .B(ram[1226]), .A(ram[1162]), .S(n10671), .Y(n8892) );
  MUX2X1 U10067 ( .B(ram[1354]), .A(ram[1290]), .S(n10671), .Y(n8896) );
  MUX2X1 U10068 ( .B(ram[1482]), .A(ram[1418]), .S(n10671), .Y(n8895) );
  MUX2X1 U10069 ( .B(n8894), .A(n8891), .S(n10571), .Y(n8905) );
  MUX2X1 U10070 ( .B(ram[1610]), .A(ram[1546]), .S(n10672), .Y(n8899) );
  MUX2X1 U10071 ( .B(ram[1738]), .A(ram[1674]), .S(n10672), .Y(n8898) );
  MUX2X1 U10072 ( .B(ram[1866]), .A(ram[1802]), .S(n10672), .Y(n8902) );
  MUX2X1 U10073 ( .B(ram[1994]), .A(ram[1930]), .S(n10672), .Y(n8901) );
  MUX2X1 U10074 ( .B(n8900), .A(n8897), .S(n10571), .Y(n8904) );
  MUX2X1 U10075 ( .B(n8903), .A(n8888), .S(n10562), .Y(n10506) );
  MUX2X1 U10076 ( .B(ram[75]), .A(ram[11]), .S(n10672), .Y(n8908) );
  MUX2X1 U10077 ( .B(ram[203]), .A(ram[139]), .S(n10672), .Y(n8907) );
  MUX2X1 U10078 ( .B(ram[331]), .A(ram[267]), .S(n10672), .Y(n8911) );
  MUX2X1 U10079 ( .B(ram[459]), .A(ram[395]), .S(n10672), .Y(n8910) );
  MUX2X1 U10080 ( .B(n8909), .A(n8906), .S(n10571), .Y(n8920) );
  MUX2X1 U10081 ( .B(ram[587]), .A(ram[523]), .S(n10672), .Y(n8914) );
  MUX2X1 U10082 ( .B(ram[715]), .A(ram[651]), .S(n10672), .Y(n8913) );
  MUX2X1 U10083 ( .B(ram[843]), .A(ram[779]), .S(n10672), .Y(n8917) );
  MUX2X1 U10084 ( .B(ram[971]), .A(ram[907]), .S(n10672), .Y(n8916) );
  MUX2X1 U10085 ( .B(n8915), .A(n8912), .S(n10571), .Y(n8919) );
  MUX2X1 U10086 ( .B(ram[1099]), .A(ram[1035]), .S(n10673), .Y(n8923) );
  MUX2X1 U10087 ( .B(ram[1227]), .A(ram[1163]), .S(n10673), .Y(n8922) );
  MUX2X1 U10088 ( .B(ram[1355]), .A(ram[1291]), .S(n10673), .Y(n8926) );
  MUX2X1 U10089 ( .B(ram[1483]), .A(ram[1419]), .S(n10673), .Y(n8925) );
  MUX2X1 U10090 ( .B(n8924), .A(n8921), .S(n10571), .Y(n8935) );
  MUX2X1 U10091 ( .B(ram[1611]), .A(ram[1547]), .S(n10673), .Y(n8929) );
  MUX2X1 U10092 ( .B(ram[1739]), .A(ram[1675]), .S(n10673), .Y(n8928) );
  MUX2X1 U10093 ( .B(ram[1867]), .A(ram[1803]), .S(n10673), .Y(n8932) );
  MUX2X1 U10094 ( .B(ram[1995]), .A(ram[1931]), .S(n10673), .Y(n8931) );
  MUX2X1 U10095 ( .B(n8930), .A(n8927), .S(n10571), .Y(n8934) );
  MUX2X1 U10096 ( .B(n8933), .A(n8918), .S(n10562), .Y(n10507) );
  MUX2X1 U10097 ( .B(ram[76]), .A(ram[12]), .S(n10673), .Y(n8938) );
  MUX2X1 U10098 ( .B(ram[204]), .A(ram[140]), .S(n10673), .Y(n8937) );
  MUX2X1 U10099 ( .B(ram[332]), .A(ram[268]), .S(n10673), .Y(n8941) );
  MUX2X1 U10100 ( .B(ram[460]), .A(ram[396]), .S(n10673), .Y(n8940) );
  MUX2X1 U10101 ( .B(n8939), .A(n8936), .S(n10571), .Y(n8950) );
  MUX2X1 U10102 ( .B(ram[588]), .A(ram[524]), .S(n10674), .Y(n8944) );
  MUX2X1 U10103 ( .B(ram[716]), .A(ram[652]), .S(n10674), .Y(n8943) );
  MUX2X1 U10104 ( .B(ram[844]), .A(ram[780]), .S(n10674), .Y(n8947) );
  MUX2X1 U10105 ( .B(ram[972]), .A(ram[908]), .S(n10674), .Y(n8946) );
  MUX2X1 U10106 ( .B(n8945), .A(n8942), .S(n10571), .Y(n8949) );
  MUX2X1 U10107 ( .B(ram[1100]), .A(ram[1036]), .S(n10674), .Y(n8953) );
  MUX2X1 U10108 ( .B(ram[1228]), .A(ram[1164]), .S(n10674), .Y(n8952) );
  MUX2X1 U10109 ( .B(ram[1356]), .A(ram[1292]), .S(n10674), .Y(n8956) );
  MUX2X1 U10110 ( .B(ram[1484]), .A(ram[1420]), .S(n10674), .Y(n8955) );
  MUX2X1 U10111 ( .B(n8954), .A(n8951), .S(n10571), .Y(n8965) );
  MUX2X1 U10112 ( .B(ram[1612]), .A(ram[1548]), .S(n10674), .Y(n8959) );
  MUX2X1 U10113 ( .B(ram[1740]), .A(ram[1676]), .S(n10674), .Y(n8958) );
  MUX2X1 U10114 ( .B(ram[1868]), .A(ram[1804]), .S(n10674), .Y(n8962) );
  MUX2X1 U10115 ( .B(ram[1996]), .A(ram[1932]), .S(n10674), .Y(n8961) );
  MUX2X1 U10116 ( .B(n8960), .A(n8957), .S(n10571), .Y(n8964) );
  MUX2X1 U10117 ( .B(n8963), .A(n8948), .S(n10561), .Y(n10508) );
  MUX2X1 U10118 ( .B(ram[77]), .A(ram[13]), .S(n10675), .Y(n8968) );
  MUX2X1 U10119 ( .B(ram[205]), .A(ram[141]), .S(n10675), .Y(n8967) );
  MUX2X1 U10120 ( .B(ram[333]), .A(ram[269]), .S(n10675), .Y(n8971) );
  MUX2X1 U10121 ( .B(ram[461]), .A(ram[397]), .S(n10675), .Y(n8970) );
  MUX2X1 U10122 ( .B(n8969), .A(n8966), .S(n10572), .Y(n8980) );
  MUX2X1 U10123 ( .B(ram[589]), .A(ram[525]), .S(n10675), .Y(n8974) );
  MUX2X1 U10124 ( .B(ram[717]), .A(ram[653]), .S(n10675), .Y(n8973) );
  MUX2X1 U10125 ( .B(ram[845]), .A(ram[781]), .S(n10675), .Y(n8977) );
  MUX2X1 U10126 ( .B(ram[973]), .A(ram[909]), .S(n10675), .Y(n8976) );
  MUX2X1 U10127 ( .B(n8975), .A(n8972), .S(n10572), .Y(n8979) );
  MUX2X1 U10128 ( .B(ram[1101]), .A(ram[1037]), .S(n10675), .Y(n8983) );
  MUX2X1 U10129 ( .B(ram[1229]), .A(ram[1165]), .S(n10675), .Y(n8982) );
  MUX2X1 U10130 ( .B(ram[1357]), .A(ram[1293]), .S(n10675), .Y(n8986) );
  MUX2X1 U10131 ( .B(ram[1485]), .A(ram[1421]), .S(n10675), .Y(n8985) );
  MUX2X1 U10132 ( .B(n8984), .A(n8981), .S(n10572), .Y(n8995) );
  MUX2X1 U10133 ( .B(ram[1613]), .A(ram[1549]), .S(n10676), .Y(n8989) );
  MUX2X1 U10134 ( .B(ram[1741]), .A(ram[1677]), .S(n10676), .Y(n8988) );
  MUX2X1 U10135 ( .B(ram[1869]), .A(ram[1805]), .S(n10676), .Y(n8992) );
  MUX2X1 U10136 ( .B(ram[1997]), .A(ram[1933]), .S(n10676), .Y(n8991) );
  MUX2X1 U10137 ( .B(n8990), .A(n8987), .S(n10572), .Y(n8994) );
  MUX2X1 U10138 ( .B(n8993), .A(n8978), .S(n10561), .Y(n10509) );
  MUX2X1 U10139 ( .B(ram[78]), .A(ram[14]), .S(n10676), .Y(n8998) );
  MUX2X1 U10140 ( .B(ram[206]), .A(ram[142]), .S(n10676), .Y(n8997) );
  MUX2X1 U10141 ( .B(ram[334]), .A(ram[270]), .S(n10676), .Y(n9001) );
  MUX2X1 U10142 ( .B(ram[462]), .A(ram[398]), .S(n10676), .Y(n9000) );
  MUX2X1 U10143 ( .B(n8999), .A(n8996), .S(n10572), .Y(n9010) );
  MUX2X1 U10144 ( .B(ram[590]), .A(ram[526]), .S(n10676), .Y(n9004) );
  MUX2X1 U10145 ( .B(ram[718]), .A(ram[654]), .S(n10676), .Y(n9003) );
  MUX2X1 U10146 ( .B(ram[846]), .A(ram[782]), .S(n10676), .Y(n9007) );
  MUX2X1 U10147 ( .B(ram[974]), .A(ram[910]), .S(n10676), .Y(n9006) );
  MUX2X1 U10148 ( .B(n9005), .A(n9002), .S(n10572), .Y(n9009) );
  MUX2X1 U10149 ( .B(ram[1102]), .A(ram[1038]), .S(n10677), .Y(n9013) );
  MUX2X1 U10150 ( .B(ram[1230]), .A(ram[1166]), .S(n10677), .Y(n9012) );
  MUX2X1 U10151 ( .B(ram[1358]), .A(ram[1294]), .S(n10677), .Y(n9016) );
  MUX2X1 U10152 ( .B(ram[1486]), .A(ram[1422]), .S(n10677), .Y(n9015) );
  MUX2X1 U10153 ( .B(n9014), .A(n9011), .S(n10572), .Y(n9025) );
  MUX2X1 U10154 ( .B(ram[1614]), .A(ram[1550]), .S(n10677), .Y(n9019) );
  MUX2X1 U10155 ( .B(ram[1742]), .A(ram[1678]), .S(n10677), .Y(n9018) );
  MUX2X1 U10156 ( .B(ram[1870]), .A(ram[1806]), .S(n10677), .Y(n9022) );
  MUX2X1 U10157 ( .B(ram[1998]), .A(ram[1934]), .S(n10677), .Y(n9021) );
  MUX2X1 U10158 ( .B(n9020), .A(n9017), .S(n10572), .Y(n9024) );
  MUX2X1 U10159 ( .B(n9023), .A(n9008), .S(n10561), .Y(n10510) );
  MUX2X1 U10160 ( .B(ram[79]), .A(ram[15]), .S(n10677), .Y(n9028) );
  MUX2X1 U10161 ( .B(ram[207]), .A(ram[143]), .S(n10677), .Y(n9027) );
  MUX2X1 U10162 ( .B(ram[335]), .A(ram[271]), .S(n10677), .Y(n9031) );
  MUX2X1 U10163 ( .B(ram[463]), .A(ram[399]), .S(n10677), .Y(n9030) );
  MUX2X1 U10164 ( .B(n9029), .A(n9026), .S(n10572), .Y(n9040) );
  MUX2X1 U10165 ( .B(ram[591]), .A(ram[527]), .S(n10678), .Y(n9034) );
  MUX2X1 U10166 ( .B(ram[719]), .A(ram[655]), .S(n10678), .Y(n9033) );
  MUX2X1 U10167 ( .B(ram[847]), .A(ram[783]), .S(n10678), .Y(n9037) );
  MUX2X1 U10168 ( .B(ram[975]), .A(ram[911]), .S(n10678), .Y(n9036) );
  MUX2X1 U10169 ( .B(n9035), .A(n9032), .S(n10572), .Y(n9039) );
  MUX2X1 U10170 ( .B(ram[1103]), .A(ram[1039]), .S(n10678), .Y(n9043) );
  MUX2X1 U10171 ( .B(ram[1231]), .A(ram[1167]), .S(n10678), .Y(n9042) );
  MUX2X1 U10172 ( .B(ram[1359]), .A(ram[1295]), .S(n10678), .Y(n9046) );
  MUX2X1 U10173 ( .B(ram[1487]), .A(ram[1423]), .S(n10678), .Y(n9045) );
  MUX2X1 U10174 ( .B(n9044), .A(n9041), .S(n10572), .Y(n9055) );
  MUX2X1 U10175 ( .B(ram[1615]), .A(ram[1551]), .S(n10678), .Y(n9049) );
  MUX2X1 U10176 ( .B(ram[1743]), .A(ram[1679]), .S(n10678), .Y(n9048) );
  MUX2X1 U10177 ( .B(ram[1871]), .A(ram[1807]), .S(n10678), .Y(n9052) );
  MUX2X1 U10178 ( .B(ram[1999]), .A(ram[1935]), .S(n10678), .Y(n9051) );
  MUX2X1 U10179 ( .B(n9050), .A(n9047), .S(n10572), .Y(n9054) );
  MUX2X1 U10180 ( .B(n9053), .A(n9038), .S(n10561), .Y(n10511) );
  MUX2X1 U10181 ( .B(ram[80]), .A(ram[16]), .S(n10679), .Y(n9058) );
  MUX2X1 U10182 ( .B(ram[208]), .A(ram[144]), .S(n10679), .Y(n9057) );
  MUX2X1 U10183 ( .B(ram[336]), .A(ram[272]), .S(n10679), .Y(n9061) );
  MUX2X1 U10184 ( .B(ram[464]), .A(ram[400]), .S(n10679), .Y(n9060) );
  MUX2X1 U10185 ( .B(n9059), .A(n9056), .S(n10573), .Y(n9070) );
  MUX2X1 U10186 ( .B(ram[592]), .A(ram[528]), .S(n10679), .Y(n9064) );
  MUX2X1 U10187 ( .B(ram[720]), .A(ram[656]), .S(n10679), .Y(n9063) );
  MUX2X1 U10188 ( .B(ram[848]), .A(ram[784]), .S(n10679), .Y(n9067) );
  MUX2X1 U10189 ( .B(ram[976]), .A(ram[912]), .S(n10679), .Y(n9066) );
  MUX2X1 U10190 ( .B(n9065), .A(n9062), .S(n10573), .Y(n9069) );
  MUX2X1 U10191 ( .B(ram[1104]), .A(ram[1040]), .S(n10679), .Y(n9073) );
  MUX2X1 U10192 ( .B(ram[1232]), .A(ram[1168]), .S(n10679), .Y(n9072) );
  MUX2X1 U10193 ( .B(ram[1360]), .A(ram[1296]), .S(n10679), .Y(n9076) );
  MUX2X1 U10194 ( .B(ram[1488]), .A(ram[1424]), .S(n10679), .Y(n9075) );
  MUX2X1 U10195 ( .B(n9074), .A(n9071), .S(n10573), .Y(n9085) );
  MUX2X1 U10196 ( .B(ram[1616]), .A(ram[1552]), .S(n10680), .Y(n9079) );
  MUX2X1 U10197 ( .B(ram[1744]), .A(ram[1680]), .S(n10680), .Y(n9078) );
  MUX2X1 U10198 ( .B(ram[1872]), .A(ram[1808]), .S(n10680), .Y(n9082) );
  MUX2X1 U10199 ( .B(ram[2000]), .A(ram[1936]), .S(n10680), .Y(n9081) );
  MUX2X1 U10200 ( .B(n9080), .A(n9077), .S(n10573), .Y(n9084) );
  MUX2X1 U10201 ( .B(n9083), .A(n9068), .S(n10561), .Y(n10512) );
  MUX2X1 U10202 ( .B(ram[81]), .A(ram[17]), .S(n10680), .Y(n9088) );
  MUX2X1 U10203 ( .B(ram[209]), .A(ram[145]), .S(n10680), .Y(n9087) );
  MUX2X1 U10204 ( .B(ram[337]), .A(ram[273]), .S(n10680), .Y(n9091) );
  MUX2X1 U10205 ( .B(ram[465]), .A(ram[401]), .S(n10680), .Y(n9090) );
  MUX2X1 U10206 ( .B(n9089), .A(n9086), .S(n10573), .Y(n9100) );
  MUX2X1 U10207 ( .B(ram[593]), .A(ram[529]), .S(n10680), .Y(n9094) );
  MUX2X1 U10208 ( .B(ram[721]), .A(ram[657]), .S(n10680), .Y(n9093) );
  MUX2X1 U10209 ( .B(ram[849]), .A(ram[785]), .S(n10680), .Y(n9097) );
  MUX2X1 U10210 ( .B(ram[977]), .A(ram[913]), .S(n10680), .Y(n9096) );
  MUX2X1 U10211 ( .B(n9095), .A(n9092), .S(n10573), .Y(n9099) );
  MUX2X1 U10212 ( .B(ram[1105]), .A(ram[1041]), .S(n10681), .Y(n9103) );
  MUX2X1 U10213 ( .B(ram[1233]), .A(ram[1169]), .S(n10681), .Y(n9102) );
  MUX2X1 U10214 ( .B(ram[1361]), .A(ram[1297]), .S(n10681), .Y(n9106) );
  MUX2X1 U10215 ( .B(ram[1489]), .A(ram[1425]), .S(n10681), .Y(n9105) );
  MUX2X1 U10216 ( .B(n9104), .A(n9101), .S(n10573), .Y(n9115) );
  MUX2X1 U10217 ( .B(ram[1617]), .A(ram[1553]), .S(n10681), .Y(n9109) );
  MUX2X1 U10218 ( .B(ram[1745]), .A(ram[1681]), .S(n10681), .Y(n9108) );
  MUX2X1 U10219 ( .B(ram[1873]), .A(ram[1809]), .S(n10681), .Y(n9112) );
  MUX2X1 U10220 ( .B(ram[2001]), .A(ram[1937]), .S(n10681), .Y(n9111) );
  MUX2X1 U10221 ( .B(n9110), .A(n9107), .S(n10573), .Y(n9114) );
  MUX2X1 U10222 ( .B(n9113), .A(n9098), .S(n10561), .Y(n10513) );
  MUX2X1 U10223 ( .B(ram[82]), .A(ram[18]), .S(n10681), .Y(n9118) );
  MUX2X1 U10224 ( .B(ram[210]), .A(ram[146]), .S(n10681), .Y(n9117) );
  MUX2X1 U10225 ( .B(ram[338]), .A(ram[274]), .S(n10681), .Y(n9121) );
  MUX2X1 U10226 ( .B(ram[466]), .A(ram[402]), .S(n10681), .Y(n9120) );
  MUX2X1 U10227 ( .B(n9119), .A(n9116), .S(n10573), .Y(n9130) );
  MUX2X1 U10228 ( .B(ram[594]), .A(ram[530]), .S(n10682), .Y(n9124) );
  MUX2X1 U10229 ( .B(ram[722]), .A(ram[658]), .S(n10682), .Y(n9123) );
  MUX2X1 U10230 ( .B(ram[850]), .A(ram[786]), .S(n10682), .Y(n9127) );
  MUX2X1 U10231 ( .B(ram[978]), .A(ram[914]), .S(n10682), .Y(n9126) );
  MUX2X1 U10232 ( .B(n9125), .A(n9122), .S(n10573), .Y(n9129) );
  MUX2X1 U10233 ( .B(ram[1106]), .A(ram[1042]), .S(n10682), .Y(n9133) );
  MUX2X1 U10234 ( .B(ram[1234]), .A(ram[1170]), .S(n10682), .Y(n9132) );
  MUX2X1 U10235 ( .B(ram[1362]), .A(ram[1298]), .S(n10682), .Y(n9136) );
  MUX2X1 U10236 ( .B(ram[1490]), .A(ram[1426]), .S(n10682), .Y(n9135) );
  MUX2X1 U10237 ( .B(n9134), .A(n9131), .S(n10573), .Y(n9145) );
  MUX2X1 U10238 ( .B(ram[1618]), .A(ram[1554]), .S(n10682), .Y(n9139) );
  MUX2X1 U10239 ( .B(ram[1746]), .A(ram[1682]), .S(n10682), .Y(n9138) );
  MUX2X1 U10240 ( .B(ram[1874]), .A(ram[1810]), .S(n10682), .Y(n9142) );
  MUX2X1 U10241 ( .B(ram[2002]), .A(ram[1938]), .S(n10682), .Y(n9141) );
  MUX2X1 U10242 ( .B(n9140), .A(n9137), .S(n10573), .Y(n9144) );
  MUX2X1 U10243 ( .B(n9143), .A(n9128), .S(n10561), .Y(n10514) );
  MUX2X1 U10244 ( .B(ram[83]), .A(ram[19]), .S(n10683), .Y(n9148) );
  MUX2X1 U10245 ( .B(ram[211]), .A(ram[147]), .S(n10683), .Y(n9147) );
  MUX2X1 U10246 ( .B(ram[339]), .A(ram[275]), .S(n10683), .Y(n9151) );
  MUX2X1 U10247 ( .B(ram[467]), .A(ram[403]), .S(n10683), .Y(n9150) );
  MUX2X1 U10248 ( .B(n9149), .A(n9146), .S(n10574), .Y(n9160) );
  MUX2X1 U10249 ( .B(ram[595]), .A(ram[531]), .S(n10683), .Y(n9154) );
  MUX2X1 U10250 ( .B(ram[723]), .A(ram[659]), .S(n10683), .Y(n9153) );
  MUX2X1 U10251 ( .B(ram[851]), .A(ram[787]), .S(n10683), .Y(n9157) );
  MUX2X1 U10252 ( .B(ram[979]), .A(ram[915]), .S(n10683), .Y(n9156) );
  MUX2X1 U10253 ( .B(n9155), .A(n9152), .S(n10574), .Y(n9159) );
  MUX2X1 U10254 ( .B(ram[1107]), .A(ram[1043]), .S(n10683), .Y(n9163) );
  MUX2X1 U10255 ( .B(ram[1235]), .A(ram[1171]), .S(n10683), .Y(n9162) );
  MUX2X1 U10256 ( .B(ram[1363]), .A(ram[1299]), .S(n10683), .Y(n9166) );
  MUX2X1 U10257 ( .B(ram[1491]), .A(ram[1427]), .S(n10683), .Y(n9165) );
  MUX2X1 U10258 ( .B(n9164), .A(n9161), .S(n10574), .Y(n9175) );
  MUX2X1 U10259 ( .B(ram[1619]), .A(ram[1555]), .S(n10684), .Y(n9169) );
  MUX2X1 U10260 ( .B(ram[1747]), .A(ram[1683]), .S(n10684), .Y(n9168) );
  MUX2X1 U10261 ( .B(ram[1875]), .A(ram[1811]), .S(n10684), .Y(n9172) );
  MUX2X1 U10262 ( .B(ram[2003]), .A(ram[1939]), .S(n10684), .Y(n9171) );
  MUX2X1 U10263 ( .B(n9170), .A(n9167), .S(n10574), .Y(n9174) );
  MUX2X1 U10264 ( .B(n9173), .A(n9158), .S(n10561), .Y(n10515) );
  MUX2X1 U10265 ( .B(ram[84]), .A(ram[20]), .S(n10684), .Y(n9178) );
  MUX2X1 U10266 ( .B(ram[212]), .A(ram[148]), .S(n10684), .Y(n9177) );
  MUX2X1 U10267 ( .B(ram[340]), .A(ram[276]), .S(n10684), .Y(n9181) );
  MUX2X1 U10268 ( .B(ram[468]), .A(ram[404]), .S(n10684), .Y(n9180) );
  MUX2X1 U10269 ( .B(n9179), .A(n9176), .S(n10574), .Y(n9190) );
  MUX2X1 U10270 ( .B(ram[596]), .A(ram[532]), .S(n10684), .Y(n9184) );
  MUX2X1 U10271 ( .B(ram[724]), .A(ram[660]), .S(n10684), .Y(n9183) );
  MUX2X1 U10272 ( .B(ram[852]), .A(ram[788]), .S(n10684), .Y(n9187) );
  MUX2X1 U10273 ( .B(ram[980]), .A(ram[916]), .S(n10684), .Y(n9186) );
  MUX2X1 U10274 ( .B(n9185), .A(n9182), .S(n10574), .Y(n9189) );
  MUX2X1 U10275 ( .B(ram[1108]), .A(ram[1044]), .S(n10685), .Y(n9193) );
  MUX2X1 U10276 ( .B(ram[1236]), .A(ram[1172]), .S(n10685), .Y(n9192) );
  MUX2X1 U10277 ( .B(ram[1364]), .A(ram[1300]), .S(n10685), .Y(n9196) );
  MUX2X1 U10278 ( .B(ram[1492]), .A(ram[1428]), .S(n10685), .Y(n9195) );
  MUX2X1 U10279 ( .B(n9194), .A(n9191), .S(n10574), .Y(n9205) );
  MUX2X1 U10280 ( .B(ram[1620]), .A(ram[1556]), .S(n10685), .Y(n9199) );
  MUX2X1 U10281 ( .B(ram[1748]), .A(ram[1684]), .S(n10685), .Y(n9198) );
  MUX2X1 U10282 ( .B(ram[1876]), .A(ram[1812]), .S(n10685), .Y(n9202) );
  MUX2X1 U10283 ( .B(ram[2004]), .A(ram[1940]), .S(n10685), .Y(n9201) );
  MUX2X1 U10284 ( .B(n9200), .A(n9197), .S(n10574), .Y(n9204) );
  MUX2X1 U10285 ( .B(n9203), .A(n9188), .S(n10561), .Y(n10516) );
  MUX2X1 U10286 ( .B(ram[85]), .A(ram[21]), .S(n10685), .Y(n9208) );
  MUX2X1 U10287 ( .B(ram[213]), .A(ram[149]), .S(n10685), .Y(n9207) );
  MUX2X1 U10288 ( .B(ram[341]), .A(ram[277]), .S(n10685), .Y(n9211) );
  MUX2X1 U10289 ( .B(ram[469]), .A(ram[405]), .S(n10685), .Y(n9210) );
  MUX2X1 U10290 ( .B(n9209), .A(n9206), .S(n10574), .Y(n9220) );
  MUX2X1 U10291 ( .B(ram[597]), .A(ram[533]), .S(n10686), .Y(n9214) );
  MUX2X1 U10292 ( .B(ram[725]), .A(ram[661]), .S(n10686), .Y(n9213) );
  MUX2X1 U10293 ( .B(ram[853]), .A(ram[789]), .S(n10686), .Y(n9217) );
  MUX2X1 U10294 ( .B(ram[981]), .A(ram[917]), .S(n10686), .Y(n9216) );
  MUX2X1 U10295 ( .B(n9215), .A(n9212), .S(n10574), .Y(n9219) );
  MUX2X1 U10296 ( .B(ram[1109]), .A(ram[1045]), .S(n10686), .Y(n9223) );
  MUX2X1 U10297 ( .B(ram[1237]), .A(ram[1173]), .S(n10686), .Y(n9222) );
  MUX2X1 U10298 ( .B(ram[1365]), .A(ram[1301]), .S(n10686), .Y(n9226) );
  MUX2X1 U10299 ( .B(ram[1493]), .A(ram[1429]), .S(n10686), .Y(n9225) );
  MUX2X1 U10300 ( .B(n9224), .A(n9221), .S(n10574), .Y(n9235) );
  MUX2X1 U10301 ( .B(ram[1621]), .A(ram[1557]), .S(n10686), .Y(n9229) );
  MUX2X1 U10302 ( .B(ram[1749]), .A(ram[1685]), .S(n10686), .Y(n9228) );
  MUX2X1 U10303 ( .B(ram[1877]), .A(ram[1813]), .S(n10686), .Y(n9232) );
  MUX2X1 U10304 ( .B(ram[2005]), .A(ram[1941]), .S(n10686), .Y(n9231) );
  MUX2X1 U10305 ( .B(n9230), .A(n9227), .S(n10574), .Y(n9234) );
  MUX2X1 U10306 ( .B(n9233), .A(n9218), .S(n10561), .Y(n10517) );
  MUX2X1 U10307 ( .B(ram[86]), .A(ram[22]), .S(n10687), .Y(n9238) );
  MUX2X1 U10308 ( .B(ram[214]), .A(ram[150]), .S(n10687), .Y(n9237) );
  MUX2X1 U10309 ( .B(ram[342]), .A(ram[278]), .S(n10687), .Y(n9241) );
  MUX2X1 U10310 ( .B(ram[470]), .A(ram[406]), .S(n10687), .Y(n9240) );
  MUX2X1 U10311 ( .B(n9239), .A(n9236), .S(n10575), .Y(n9250) );
  MUX2X1 U10312 ( .B(ram[598]), .A(ram[534]), .S(n10687), .Y(n9244) );
  MUX2X1 U10313 ( .B(ram[726]), .A(ram[662]), .S(n10687), .Y(n9243) );
  MUX2X1 U10314 ( .B(ram[854]), .A(ram[790]), .S(n10687), .Y(n9247) );
  MUX2X1 U10315 ( .B(ram[982]), .A(ram[918]), .S(n10687), .Y(n9246) );
  MUX2X1 U10316 ( .B(n9245), .A(n9242), .S(n10575), .Y(n9249) );
  MUX2X1 U10317 ( .B(ram[1110]), .A(ram[1046]), .S(n10687), .Y(n9253) );
  MUX2X1 U10318 ( .B(ram[1238]), .A(ram[1174]), .S(n10687), .Y(n9252) );
  MUX2X1 U10319 ( .B(ram[1366]), .A(ram[1302]), .S(n10687), .Y(n9256) );
  MUX2X1 U10320 ( .B(ram[1494]), .A(ram[1430]), .S(n10687), .Y(n9255) );
  MUX2X1 U10321 ( .B(n9254), .A(n9251), .S(n10575), .Y(n9265) );
  MUX2X1 U10322 ( .B(ram[1622]), .A(ram[1558]), .S(n10688), .Y(n9259) );
  MUX2X1 U10323 ( .B(ram[1750]), .A(ram[1686]), .S(n10688), .Y(n9258) );
  MUX2X1 U10324 ( .B(ram[1878]), .A(ram[1814]), .S(n10688), .Y(n9262) );
  MUX2X1 U10325 ( .B(ram[2006]), .A(ram[1942]), .S(n10688), .Y(n9261) );
  MUX2X1 U10326 ( .B(n9260), .A(n9257), .S(n10575), .Y(n9264) );
  MUX2X1 U10327 ( .B(n9263), .A(n9248), .S(n10561), .Y(n10518) );
  MUX2X1 U10328 ( .B(ram[87]), .A(ram[23]), .S(n10688), .Y(n9268) );
  MUX2X1 U10329 ( .B(ram[215]), .A(ram[151]), .S(n10688), .Y(n9267) );
  MUX2X1 U10330 ( .B(ram[343]), .A(ram[279]), .S(n10688), .Y(n9271) );
  MUX2X1 U10331 ( .B(ram[471]), .A(ram[407]), .S(n10688), .Y(n9270) );
  MUX2X1 U10332 ( .B(n9269), .A(n9266), .S(n10575), .Y(n9280) );
  MUX2X1 U10333 ( .B(ram[599]), .A(ram[535]), .S(n10688), .Y(n9274) );
  MUX2X1 U10334 ( .B(ram[727]), .A(ram[663]), .S(n10688), .Y(n9273) );
  MUX2X1 U10335 ( .B(ram[855]), .A(ram[791]), .S(n10688), .Y(n9277) );
  MUX2X1 U10336 ( .B(ram[983]), .A(ram[919]), .S(n10688), .Y(n9276) );
  MUX2X1 U10337 ( .B(n9275), .A(n9272), .S(n10575), .Y(n9279) );
  MUX2X1 U10338 ( .B(ram[1111]), .A(ram[1047]), .S(n10689), .Y(n9283) );
  MUX2X1 U10339 ( .B(ram[1239]), .A(ram[1175]), .S(n10689), .Y(n9282) );
  MUX2X1 U10340 ( .B(ram[1367]), .A(ram[1303]), .S(n10689), .Y(n9286) );
  MUX2X1 U10341 ( .B(ram[1495]), .A(ram[1431]), .S(n10689), .Y(n9285) );
  MUX2X1 U10342 ( .B(n9284), .A(n9281), .S(n10575), .Y(n9295) );
  MUX2X1 U10343 ( .B(ram[1623]), .A(ram[1559]), .S(n10689), .Y(n9289) );
  MUX2X1 U10344 ( .B(ram[1751]), .A(ram[1687]), .S(n10689), .Y(n9288) );
  MUX2X1 U10345 ( .B(ram[1879]), .A(ram[1815]), .S(n10689), .Y(n9292) );
  MUX2X1 U10346 ( .B(ram[2007]), .A(ram[1943]), .S(n10689), .Y(n9291) );
  MUX2X1 U10347 ( .B(n9290), .A(n9287), .S(n10575), .Y(n9294) );
  MUX2X1 U10348 ( .B(n9293), .A(n9278), .S(n10561), .Y(n10519) );
  MUX2X1 U10349 ( .B(ram[88]), .A(ram[24]), .S(n10689), .Y(n9298) );
  MUX2X1 U10350 ( .B(ram[216]), .A(ram[152]), .S(n10689), .Y(n9297) );
  MUX2X1 U10351 ( .B(ram[344]), .A(ram[280]), .S(n10689), .Y(n9301) );
  MUX2X1 U10352 ( .B(ram[472]), .A(ram[408]), .S(n10689), .Y(n9300) );
  MUX2X1 U10353 ( .B(n9299), .A(n9296), .S(n10575), .Y(n9310) );
  MUX2X1 U10354 ( .B(ram[600]), .A(ram[536]), .S(n10690), .Y(n9304) );
  MUX2X1 U10355 ( .B(ram[728]), .A(ram[664]), .S(n10690), .Y(n9303) );
  MUX2X1 U10356 ( .B(ram[856]), .A(ram[792]), .S(n10690), .Y(n9307) );
  MUX2X1 U10357 ( .B(ram[984]), .A(ram[920]), .S(n10690), .Y(n9306) );
  MUX2X1 U10358 ( .B(n9305), .A(n9302), .S(n10575), .Y(n9309) );
  MUX2X1 U10359 ( .B(ram[1112]), .A(ram[1048]), .S(n10690), .Y(n9313) );
  MUX2X1 U10360 ( .B(ram[1240]), .A(ram[1176]), .S(n10690), .Y(n9312) );
  MUX2X1 U10361 ( .B(ram[1368]), .A(ram[1304]), .S(n10690), .Y(n9316) );
  MUX2X1 U10362 ( .B(ram[1496]), .A(ram[1432]), .S(n10690), .Y(n9315) );
  MUX2X1 U10363 ( .B(n9314), .A(n9311), .S(n10575), .Y(n9325) );
  MUX2X1 U10364 ( .B(ram[1624]), .A(ram[1560]), .S(n10690), .Y(n9319) );
  MUX2X1 U10365 ( .B(ram[1752]), .A(ram[1688]), .S(n10690), .Y(n9318) );
  MUX2X1 U10366 ( .B(ram[1880]), .A(ram[1816]), .S(n10690), .Y(n9322) );
  MUX2X1 U10367 ( .B(ram[2008]), .A(ram[1944]), .S(n10690), .Y(n9321) );
  MUX2X1 U10368 ( .B(n9320), .A(n9317), .S(n10575), .Y(n9324) );
  MUX2X1 U10369 ( .B(n9323), .A(n9308), .S(read2_addr[0]), .Y(n10520) );
  MUX2X1 U10370 ( .B(ram[89]), .A(ram[25]), .S(n10691), .Y(n9328) );
  MUX2X1 U10371 ( .B(ram[217]), .A(ram[153]), .S(n10691), .Y(n9327) );
  MUX2X1 U10372 ( .B(ram[345]), .A(ram[281]), .S(n10691), .Y(n9331) );
  MUX2X1 U10373 ( .B(ram[473]), .A(ram[409]), .S(n10691), .Y(n9330) );
  MUX2X1 U10374 ( .B(n9329), .A(n9326), .S(n10576), .Y(n9340) );
  MUX2X1 U10375 ( .B(ram[601]), .A(ram[537]), .S(n10691), .Y(n9334) );
  MUX2X1 U10376 ( .B(ram[729]), .A(ram[665]), .S(n10691), .Y(n9333) );
  MUX2X1 U10377 ( .B(ram[857]), .A(ram[793]), .S(n10691), .Y(n9337) );
  MUX2X1 U10378 ( .B(ram[985]), .A(ram[921]), .S(n10691), .Y(n9336) );
  MUX2X1 U10379 ( .B(n9335), .A(n9332), .S(n10576), .Y(n9339) );
  MUX2X1 U10380 ( .B(ram[1113]), .A(ram[1049]), .S(n10691), .Y(n9343) );
  MUX2X1 U10381 ( .B(ram[1241]), .A(ram[1177]), .S(n10691), .Y(n9342) );
  MUX2X1 U10382 ( .B(ram[1369]), .A(ram[1305]), .S(n10691), .Y(n9346) );
  MUX2X1 U10383 ( .B(ram[1497]), .A(ram[1433]), .S(n10691), .Y(n9345) );
  MUX2X1 U10384 ( .B(n9344), .A(n9341), .S(n10576), .Y(n9355) );
  MUX2X1 U10385 ( .B(ram[1625]), .A(ram[1561]), .S(n10692), .Y(n9349) );
  MUX2X1 U10386 ( .B(ram[1753]), .A(ram[1689]), .S(n10692), .Y(n9348) );
  MUX2X1 U10387 ( .B(ram[1881]), .A(ram[1817]), .S(n10692), .Y(n9352) );
  MUX2X1 U10388 ( .B(ram[2009]), .A(ram[1945]), .S(n10692), .Y(n9351) );
  MUX2X1 U10389 ( .B(n9350), .A(n9347), .S(n10576), .Y(n9354) );
  MUX2X1 U10390 ( .B(n9353), .A(n9338), .S(read2_addr[0]), .Y(n10521) );
  MUX2X1 U10391 ( .B(ram[90]), .A(ram[26]), .S(n10692), .Y(n9358) );
  MUX2X1 U10392 ( .B(ram[218]), .A(ram[154]), .S(n10692), .Y(n9357) );
  MUX2X1 U10393 ( .B(ram[346]), .A(ram[282]), .S(n10692), .Y(n9361) );
  MUX2X1 U10394 ( .B(ram[474]), .A(ram[410]), .S(n10692), .Y(n9360) );
  MUX2X1 U10395 ( .B(n9359), .A(n9356), .S(n10576), .Y(n9370) );
  MUX2X1 U10396 ( .B(ram[602]), .A(ram[538]), .S(n10692), .Y(n9364) );
  MUX2X1 U10397 ( .B(ram[730]), .A(ram[666]), .S(n10692), .Y(n9363) );
  MUX2X1 U10398 ( .B(ram[858]), .A(ram[794]), .S(n10692), .Y(n9367) );
  MUX2X1 U10399 ( .B(ram[986]), .A(ram[922]), .S(n10692), .Y(n9366) );
  MUX2X1 U10400 ( .B(n9365), .A(n9362), .S(n10576), .Y(n9369) );
  MUX2X1 U10401 ( .B(ram[1114]), .A(ram[1050]), .S(n10693), .Y(n9373) );
  MUX2X1 U10402 ( .B(ram[1242]), .A(ram[1178]), .S(n10693), .Y(n9372) );
  MUX2X1 U10403 ( .B(ram[1370]), .A(ram[1306]), .S(n10693), .Y(n9376) );
  MUX2X1 U10404 ( .B(ram[1498]), .A(ram[1434]), .S(n10693), .Y(n9375) );
  MUX2X1 U10405 ( .B(n9374), .A(n9371), .S(n10576), .Y(n9385) );
  MUX2X1 U10406 ( .B(ram[1626]), .A(ram[1562]), .S(n10693), .Y(n9379) );
  MUX2X1 U10407 ( .B(ram[1754]), .A(ram[1690]), .S(n10693), .Y(n9378) );
  MUX2X1 U10408 ( .B(ram[1882]), .A(ram[1818]), .S(n10693), .Y(n9382) );
  MUX2X1 U10409 ( .B(ram[2010]), .A(ram[1946]), .S(n10693), .Y(n9381) );
  MUX2X1 U10410 ( .B(n9380), .A(n9377), .S(n10576), .Y(n9384) );
  MUX2X1 U10411 ( .B(n9383), .A(n9368), .S(read2_addr[0]), .Y(n10522) );
  MUX2X1 U10412 ( .B(ram[91]), .A(ram[27]), .S(n10693), .Y(n9388) );
  MUX2X1 U10413 ( .B(ram[219]), .A(ram[155]), .S(n10693), .Y(n9387) );
  MUX2X1 U10414 ( .B(ram[347]), .A(ram[283]), .S(n10693), .Y(n9391) );
  MUX2X1 U10415 ( .B(ram[475]), .A(ram[411]), .S(n10693), .Y(n9390) );
  MUX2X1 U10416 ( .B(n9389), .A(n9386), .S(n10576), .Y(n9400) );
  MUX2X1 U10417 ( .B(ram[603]), .A(ram[539]), .S(n10694), .Y(n9394) );
  MUX2X1 U10418 ( .B(ram[731]), .A(ram[667]), .S(n10694), .Y(n9393) );
  MUX2X1 U10419 ( .B(ram[859]), .A(ram[795]), .S(n10694), .Y(n9397) );
  MUX2X1 U10420 ( .B(ram[987]), .A(ram[923]), .S(n10694), .Y(n9396) );
  MUX2X1 U10421 ( .B(n9395), .A(n9392), .S(n10576), .Y(n9399) );
  MUX2X1 U10422 ( .B(ram[1115]), .A(ram[1051]), .S(n10694), .Y(n9403) );
  MUX2X1 U10423 ( .B(ram[1243]), .A(ram[1179]), .S(n10694), .Y(n9402) );
  MUX2X1 U10424 ( .B(ram[1371]), .A(ram[1307]), .S(n10694), .Y(n9406) );
  MUX2X1 U10425 ( .B(ram[1499]), .A(ram[1435]), .S(n10694), .Y(n9405) );
  MUX2X1 U10426 ( .B(n9404), .A(n9401), .S(n10576), .Y(n9415) );
  MUX2X1 U10427 ( .B(ram[1627]), .A(ram[1563]), .S(n10694), .Y(n9409) );
  MUX2X1 U10428 ( .B(ram[1755]), .A(ram[1691]), .S(n10694), .Y(n9408) );
  MUX2X1 U10429 ( .B(ram[1883]), .A(ram[1819]), .S(n10694), .Y(n9412) );
  MUX2X1 U10430 ( .B(ram[2011]), .A(ram[1947]), .S(n10694), .Y(n9411) );
  MUX2X1 U10431 ( .B(n9410), .A(n9407), .S(n10576), .Y(n9414) );
  MUX2X1 U10432 ( .B(n9413), .A(n9398), .S(read2_addr[0]), .Y(n10523) );
  MUX2X1 U10433 ( .B(ram[92]), .A(ram[28]), .S(n10695), .Y(n9418) );
  MUX2X1 U10434 ( .B(ram[220]), .A(ram[156]), .S(n10695), .Y(n9417) );
  MUX2X1 U10435 ( .B(ram[348]), .A(ram[284]), .S(n10695), .Y(n9421) );
  MUX2X1 U10436 ( .B(ram[476]), .A(ram[412]), .S(n10695), .Y(n9420) );
  MUX2X1 U10437 ( .B(n9419), .A(n9416), .S(n10577), .Y(n9430) );
  MUX2X1 U10438 ( .B(ram[604]), .A(ram[540]), .S(n10695), .Y(n9424) );
  MUX2X1 U10439 ( .B(ram[732]), .A(ram[668]), .S(n10695), .Y(n9423) );
  MUX2X1 U10440 ( .B(ram[860]), .A(ram[796]), .S(n10695), .Y(n9427) );
  MUX2X1 U10441 ( .B(ram[988]), .A(ram[924]), .S(n10695), .Y(n9426) );
  MUX2X1 U10442 ( .B(n9425), .A(n9422), .S(n10577), .Y(n9429) );
  MUX2X1 U10443 ( .B(ram[1116]), .A(ram[1052]), .S(n10695), .Y(n9433) );
  MUX2X1 U10444 ( .B(ram[1244]), .A(ram[1180]), .S(n10695), .Y(n9432) );
  MUX2X1 U10445 ( .B(ram[1372]), .A(ram[1308]), .S(n10695), .Y(n9436) );
  MUX2X1 U10446 ( .B(ram[1500]), .A(ram[1436]), .S(n10695), .Y(n9435) );
  MUX2X1 U10447 ( .B(n9434), .A(n9431), .S(n10577), .Y(n9445) );
  MUX2X1 U10448 ( .B(ram[1628]), .A(ram[1564]), .S(n10696), .Y(n9439) );
  MUX2X1 U10449 ( .B(ram[1756]), .A(ram[1692]), .S(n10696), .Y(n9438) );
  MUX2X1 U10450 ( .B(ram[1884]), .A(ram[1820]), .S(n10696), .Y(n9442) );
  MUX2X1 U10451 ( .B(ram[2012]), .A(ram[1948]), .S(n10696), .Y(n9441) );
  MUX2X1 U10452 ( .B(n9440), .A(n9437), .S(n10577), .Y(n9444) );
  MUX2X1 U10453 ( .B(n9443), .A(n9428), .S(read2_addr[0]), .Y(n10524) );
  MUX2X1 U10454 ( .B(ram[93]), .A(ram[29]), .S(n10696), .Y(n9448) );
  MUX2X1 U10455 ( .B(ram[221]), .A(ram[157]), .S(n10696), .Y(n9447) );
  MUX2X1 U10456 ( .B(ram[349]), .A(ram[285]), .S(n10696), .Y(n9451) );
  MUX2X1 U10457 ( .B(ram[477]), .A(ram[413]), .S(n10696), .Y(n9450) );
  MUX2X1 U10458 ( .B(n9449), .A(n9446), .S(n10577), .Y(n9460) );
  MUX2X1 U10459 ( .B(ram[605]), .A(ram[541]), .S(n10696), .Y(n9454) );
  MUX2X1 U10460 ( .B(ram[733]), .A(ram[669]), .S(n10696), .Y(n9453) );
  MUX2X1 U10461 ( .B(ram[861]), .A(ram[797]), .S(n10696), .Y(n9457) );
  MUX2X1 U10462 ( .B(ram[989]), .A(ram[925]), .S(n10696), .Y(n9456) );
  MUX2X1 U10463 ( .B(n9455), .A(n9452), .S(n10577), .Y(n9459) );
  MUX2X1 U10464 ( .B(ram[1117]), .A(ram[1053]), .S(n10697), .Y(n9463) );
  MUX2X1 U10465 ( .B(ram[1245]), .A(ram[1181]), .S(n10697), .Y(n9462) );
  MUX2X1 U10466 ( .B(ram[1373]), .A(ram[1309]), .S(n10697), .Y(n9466) );
  MUX2X1 U10467 ( .B(ram[1501]), .A(ram[1437]), .S(n10697), .Y(n9465) );
  MUX2X1 U10468 ( .B(n9464), .A(n9461), .S(n10577), .Y(n9475) );
  MUX2X1 U10469 ( .B(ram[1629]), .A(ram[1565]), .S(n10697), .Y(n9469) );
  MUX2X1 U10470 ( .B(ram[1757]), .A(ram[1693]), .S(n10697), .Y(n9468) );
  MUX2X1 U10471 ( .B(ram[1885]), .A(ram[1821]), .S(n10697), .Y(n9472) );
  MUX2X1 U10472 ( .B(ram[2013]), .A(ram[1949]), .S(n10697), .Y(n9471) );
  MUX2X1 U10473 ( .B(n9470), .A(n9467), .S(n10577), .Y(n9474) );
  MUX2X1 U10474 ( .B(n9473), .A(n9458), .S(read2_addr[0]), .Y(n10525) );
  MUX2X1 U10475 ( .B(ram[94]), .A(ram[30]), .S(n10697), .Y(n9478) );
  MUX2X1 U10476 ( .B(ram[222]), .A(ram[158]), .S(n10697), .Y(n9477) );
  MUX2X1 U10477 ( .B(ram[350]), .A(ram[286]), .S(n10697), .Y(n9481) );
  MUX2X1 U10478 ( .B(ram[478]), .A(ram[414]), .S(n10697), .Y(n9480) );
  MUX2X1 U10479 ( .B(n9479), .A(n9476), .S(n10577), .Y(n9490) );
  MUX2X1 U10480 ( .B(ram[606]), .A(ram[542]), .S(n10698), .Y(n9484) );
  MUX2X1 U10481 ( .B(ram[734]), .A(ram[670]), .S(n10698), .Y(n9483) );
  MUX2X1 U10482 ( .B(ram[862]), .A(ram[798]), .S(n10698), .Y(n9487) );
  MUX2X1 U10483 ( .B(ram[990]), .A(ram[926]), .S(n10698), .Y(n9486) );
  MUX2X1 U10484 ( .B(n9485), .A(n9482), .S(n10577), .Y(n9489) );
  MUX2X1 U10485 ( .B(ram[1118]), .A(ram[1054]), .S(n10698), .Y(n9493) );
  MUX2X1 U10486 ( .B(ram[1246]), .A(ram[1182]), .S(n10698), .Y(n9492) );
  MUX2X1 U10487 ( .B(ram[1374]), .A(ram[1310]), .S(n10698), .Y(n9496) );
  MUX2X1 U10488 ( .B(ram[1502]), .A(ram[1438]), .S(n10698), .Y(n9495) );
  MUX2X1 U10489 ( .B(n9494), .A(n9491), .S(n10577), .Y(n9505) );
  MUX2X1 U10490 ( .B(ram[1630]), .A(ram[1566]), .S(n10698), .Y(n9499) );
  MUX2X1 U10491 ( .B(ram[1758]), .A(ram[1694]), .S(n10698), .Y(n9498) );
  MUX2X1 U10492 ( .B(ram[1886]), .A(ram[1822]), .S(n10698), .Y(n9502) );
  MUX2X1 U10493 ( .B(ram[2014]), .A(ram[1950]), .S(n10698), .Y(n9501) );
  MUX2X1 U10494 ( .B(n9500), .A(n9497), .S(n10577), .Y(n9504) );
  MUX2X1 U10495 ( .B(n9503), .A(n9488), .S(read2_addr[0]), .Y(n10526) );
  MUX2X1 U10496 ( .B(ram[95]), .A(ram[31]), .S(n10699), .Y(n9508) );
  MUX2X1 U10497 ( .B(ram[223]), .A(ram[159]), .S(n10699), .Y(n9507) );
  MUX2X1 U10498 ( .B(ram[351]), .A(ram[287]), .S(n10699), .Y(n9511) );
  MUX2X1 U10499 ( .B(ram[479]), .A(ram[415]), .S(n10699), .Y(n9510) );
  MUX2X1 U10500 ( .B(n9509), .A(n9506), .S(n10578), .Y(n9520) );
  MUX2X1 U10501 ( .B(ram[607]), .A(ram[543]), .S(n10699), .Y(n9514) );
  MUX2X1 U10502 ( .B(ram[735]), .A(ram[671]), .S(n10699), .Y(n9513) );
  MUX2X1 U10503 ( .B(ram[863]), .A(ram[799]), .S(n10699), .Y(n9517) );
  MUX2X1 U10504 ( .B(ram[991]), .A(ram[927]), .S(n10699), .Y(n9516) );
  MUX2X1 U10505 ( .B(n9515), .A(n9512), .S(n10578), .Y(n9519) );
  MUX2X1 U10506 ( .B(ram[1119]), .A(ram[1055]), .S(n10699), .Y(n9523) );
  MUX2X1 U10507 ( .B(ram[1247]), .A(ram[1183]), .S(n10699), .Y(n9522) );
  MUX2X1 U10508 ( .B(ram[1375]), .A(ram[1311]), .S(n10699), .Y(n9526) );
  MUX2X1 U10509 ( .B(ram[1503]), .A(ram[1439]), .S(n10699), .Y(n9525) );
  MUX2X1 U10510 ( .B(n9524), .A(n9521), .S(n10578), .Y(n9535) );
  MUX2X1 U10511 ( .B(ram[1631]), .A(ram[1567]), .S(n10700), .Y(n9529) );
  MUX2X1 U10512 ( .B(ram[1759]), .A(ram[1695]), .S(n10700), .Y(n9528) );
  MUX2X1 U10513 ( .B(ram[1887]), .A(ram[1823]), .S(n10700), .Y(n9532) );
  MUX2X1 U10514 ( .B(ram[2015]), .A(ram[1951]), .S(n10700), .Y(n9531) );
  MUX2X1 U10515 ( .B(n9530), .A(n9527), .S(n10578), .Y(n9534) );
  MUX2X1 U10516 ( .B(n9533), .A(n9518), .S(read2_addr[0]), .Y(n10527) );
  MUX2X1 U10517 ( .B(ram[96]), .A(ram[32]), .S(n10700), .Y(n9538) );
  MUX2X1 U10518 ( .B(ram[224]), .A(ram[160]), .S(n10700), .Y(n9537) );
  MUX2X1 U10519 ( .B(ram[352]), .A(ram[288]), .S(n10700), .Y(n9541) );
  MUX2X1 U10520 ( .B(ram[480]), .A(ram[416]), .S(n10700), .Y(n9540) );
  MUX2X1 U10521 ( .B(n9539), .A(n9536), .S(n10578), .Y(n9550) );
  MUX2X1 U10522 ( .B(ram[608]), .A(ram[544]), .S(n10700), .Y(n9544) );
  MUX2X1 U10523 ( .B(ram[736]), .A(ram[672]), .S(n10700), .Y(n9543) );
  MUX2X1 U10524 ( .B(ram[864]), .A(ram[800]), .S(n10700), .Y(n9547) );
  MUX2X1 U10525 ( .B(ram[992]), .A(ram[928]), .S(n10700), .Y(n9546) );
  MUX2X1 U10526 ( .B(n9545), .A(n9542), .S(n10578), .Y(n9549) );
  MUX2X1 U10527 ( .B(ram[1120]), .A(ram[1056]), .S(n10701), .Y(n9553) );
  MUX2X1 U10528 ( .B(ram[1248]), .A(ram[1184]), .S(n10701), .Y(n9552) );
  MUX2X1 U10529 ( .B(ram[1376]), .A(ram[1312]), .S(n10701), .Y(n9556) );
  MUX2X1 U10530 ( .B(ram[1504]), .A(ram[1440]), .S(n10701), .Y(n9555) );
  MUX2X1 U10531 ( .B(n9554), .A(n9551), .S(n10578), .Y(n9565) );
  MUX2X1 U10532 ( .B(ram[1632]), .A(ram[1568]), .S(n10701), .Y(n9559) );
  MUX2X1 U10533 ( .B(ram[1760]), .A(ram[1696]), .S(n10701), .Y(n9558) );
  MUX2X1 U10534 ( .B(ram[1888]), .A(ram[1824]), .S(n10701), .Y(n9562) );
  MUX2X1 U10535 ( .B(ram[2016]), .A(ram[1952]), .S(n10701), .Y(n9561) );
  MUX2X1 U10536 ( .B(n9560), .A(n9557), .S(n10578), .Y(n9564) );
  MUX2X1 U10537 ( .B(n9563), .A(n9548), .S(read2_addr[0]), .Y(n10528) );
  MUX2X1 U10538 ( .B(ram[97]), .A(ram[33]), .S(n10701), .Y(n9568) );
  MUX2X1 U10539 ( .B(ram[225]), .A(ram[161]), .S(n10701), .Y(n9567) );
  MUX2X1 U10540 ( .B(ram[353]), .A(ram[289]), .S(n10701), .Y(n9571) );
  MUX2X1 U10541 ( .B(ram[481]), .A(ram[417]), .S(n10701), .Y(n9570) );
  MUX2X1 U10542 ( .B(n9569), .A(n9566), .S(n10578), .Y(n9580) );
  MUX2X1 U10543 ( .B(ram[609]), .A(ram[545]), .S(n10702), .Y(n9574) );
  MUX2X1 U10544 ( .B(ram[737]), .A(ram[673]), .S(n10702), .Y(n9573) );
  MUX2X1 U10545 ( .B(ram[865]), .A(ram[801]), .S(n10702), .Y(n9577) );
  MUX2X1 U10546 ( .B(ram[993]), .A(ram[929]), .S(n10702), .Y(n9576) );
  MUX2X1 U10547 ( .B(n9575), .A(n9572), .S(n10578), .Y(n9579) );
  MUX2X1 U10548 ( .B(ram[1121]), .A(ram[1057]), .S(n10702), .Y(n9583) );
  MUX2X1 U10549 ( .B(ram[1249]), .A(ram[1185]), .S(n10702), .Y(n9582) );
  MUX2X1 U10550 ( .B(ram[1377]), .A(ram[1313]), .S(n10702), .Y(n9586) );
  MUX2X1 U10551 ( .B(ram[1505]), .A(ram[1441]), .S(n10702), .Y(n9585) );
  MUX2X1 U10552 ( .B(n9584), .A(n9581), .S(n10578), .Y(n9595) );
  MUX2X1 U10553 ( .B(ram[1633]), .A(ram[1569]), .S(n10702), .Y(n9589) );
  MUX2X1 U10554 ( .B(ram[1761]), .A(ram[1697]), .S(n10702), .Y(n9588) );
  MUX2X1 U10555 ( .B(ram[1889]), .A(ram[1825]), .S(n10702), .Y(n9592) );
  MUX2X1 U10556 ( .B(ram[2017]), .A(ram[1953]), .S(n10702), .Y(n9591) );
  MUX2X1 U10557 ( .B(n9590), .A(n9587), .S(n10578), .Y(n9594) );
  MUX2X1 U10558 ( .B(n9593), .A(n9578), .S(read2_addr[0]), .Y(n10529) );
  MUX2X1 U10559 ( .B(ram[98]), .A(ram[34]), .S(n10703), .Y(n9598) );
  MUX2X1 U10560 ( .B(ram[226]), .A(ram[162]), .S(n10703), .Y(n9597) );
  MUX2X1 U10561 ( .B(ram[354]), .A(ram[290]), .S(n10703), .Y(n9601) );
  MUX2X1 U10562 ( .B(ram[482]), .A(ram[418]), .S(n10703), .Y(n9600) );
  MUX2X1 U10563 ( .B(n9599), .A(n9596), .S(n10579), .Y(n9610) );
  MUX2X1 U10564 ( .B(ram[610]), .A(ram[546]), .S(n10703), .Y(n9604) );
  MUX2X1 U10565 ( .B(ram[738]), .A(ram[674]), .S(n10703), .Y(n9603) );
  MUX2X1 U10566 ( .B(ram[866]), .A(ram[802]), .S(n10703), .Y(n9607) );
  MUX2X1 U10567 ( .B(ram[994]), .A(ram[930]), .S(n10703), .Y(n9606) );
  MUX2X1 U10568 ( .B(n9605), .A(n9602), .S(n10579), .Y(n9609) );
  MUX2X1 U10569 ( .B(ram[1122]), .A(ram[1058]), .S(n10703), .Y(n9613) );
  MUX2X1 U10570 ( .B(ram[1250]), .A(ram[1186]), .S(n10703), .Y(n9612) );
  MUX2X1 U10571 ( .B(ram[1378]), .A(ram[1314]), .S(n10703), .Y(n9616) );
  MUX2X1 U10572 ( .B(ram[1506]), .A(ram[1442]), .S(n10703), .Y(n9615) );
  MUX2X1 U10573 ( .B(n9614), .A(n9611), .S(n10579), .Y(n9625) );
  MUX2X1 U10574 ( .B(ram[1634]), .A(ram[1570]), .S(n10704), .Y(n9619) );
  MUX2X1 U10575 ( .B(ram[1762]), .A(ram[1698]), .S(n10704), .Y(n9618) );
  MUX2X1 U10576 ( .B(ram[1890]), .A(ram[1826]), .S(n10704), .Y(n9622) );
  MUX2X1 U10577 ( .B(ram[2018]), .A(ram[1954]), .S(n10704), .Y(n9621) );
  MUX2X1 U10578 ( .B(n9620), .A(n9617), .S(n10579), .Y(n9624) );
  MUX2X1 U10579 ( .B(n9623), .A(n9608), .S(read2_addr[0]), .Y(n10530) );
  MUX2X1 U10580 ( .B(ram[99]), .A(ram[35]), .S(n10704), .Y(n9628) );
  MUX2X1 U10581 ( .B(ram[227]), .A(ram[163]), .S(n10704), .Y(n9627) );
  MUX2X1 U10582 ( .B(ram[355]), .A(ram[291]), .S(n10704), .Y(n9631) );
  MUX2X1 U10583 ( .B(ram[483]), .A(ram[419]), .S(n10704), .Y(n9630) );
  MUX2X1 U10584 ( .B(n9629), .A(n9626), .S(n10579), .Y(n9640) );
  MUX2X1 U10585 ( .B(ram[611]), .A(ram[547]), .S(n10704), .Y(n9634) );
  MUX2X1 U10586 ( .B(ram[739]), .A(ram[675]), .S(n10704), .Y(n9633) );
  MUX2X1 U10587 ( .B(ram[867]), .A(ram[803]), .S(n10704), .Y(n9637) );
  MUX2X1 U10588 ( .B(ram[995]), .A(ram[931]), .S(n10704), .Y(n9636) );
  MUX2X1 U10589 ( .B(n9635), .A(n9632), .S(n10579), .Y(n9639) );
  MUX2X1 U10590 ( .B(ram[1123]), .A(ram[1059]), .S(n10705), .Y(n9643) );
  MUX2X1 U10591 ( .B(ram[1251]), .A(ram[1187]), .S(n10705), .Y(n9642) );
  MUX2X1 U10592 ( .B(ram[1379]), .A(ram[1315]), .S(n10705), .Y(n9646) );
  MUX2X1 U10593 ( .B(ram[1507]), .A(ram[1443]), .S(n10705), .Y(n9645) );
  MUX2X1 U10594 ( .B(n9644), .A(n9641), .S(n10579), .Y(n9655) );
  MUX2X1 U10595 ( .B(ram[1635]), .A(ram[1571]), .S(n10705), .Y(n9649) );
  MUX2X1 U10596 ( .B(ram[1763]), .A(ram[1699]), .S(n10705), .Y(n9648) );
  MUX2X1 U10597 ( .B(ram[1891]), .A(ram[1827]), .S(n10705), .Y(n9652) );
  MUX2X1 U10598 ( .B(ram[2019]), .A(ram[1955]), .S(n10705), .Y(n9651) );
  MUX2X1 U10599 ( .B(n9650), .A(n9647), .S(n10579), .Y(n9654) );
  MUX2X1 U10600 ( .B(n9653), .A(n9638), .S(read2_addr[0]), .Y(n10531) );
  MUX2X1 U10601 ( .B(ram[100]), .A(ram[36]), .S(n10705), .Y(n9658) );
  MUX2X1 U10602 ( .B(ram[228]), .A(ram[164]), .S(n10705), .Y(n9657) );
  MUX2X1 U10603 ( .B(ram[356]), .A(ram[292]), .S(n10705), .Y(n9661) );
  MUX2X1 U10604 ( .B(ram[484]), .A(ram[420]), .S(n10705), .Y(n9660) );
  MUX2X1 U10605 ( .B(n9659), .A(n9656), .S(n10579), .Y(n9670) );
  MUX2X1 U10606 ( .B(ram[612]), .A(ram[548]), .S(n10706), .Y(n9664) );
  MUX2X1 U10607 ( .B(ram[740]), .A(ram[676]), .S(n10706), .Y(n9663) );
  MUX2X1 U10608 ( .B(ram[868]), .A(ram[804]), .S(n10706), .Y(n9667) );
  MUX2X1 U10609 ( .B(ram[996]), .A(ram[932]), .S(n10706), .Y(n9666) );
  MUX2X1 U10610 ( .B(n9665), .A(n9662), .S(n10579), .Y(n9669) );
  MUX2X1 U10611 ( .B(ram[1124]), .A(ram[1060]), .S(n10706), .Y(n9673) );
  MUX2X1 U10612 ( .B(ram[1252]), .A(ram[1188]), .S(n10706), .Y(n9672) );
  MUX2X1 U10613 ( .B(ram[1380]), .A(ram[1316]), .S(n10706), .Y(n9676) );
  MUX2X1 U10614 ( .B(ram[1508]), .A(ram[1444]), .S(n10706), .Y(n9675) );
  MUX2X1 U10615 ( .B(n9674), .A(n9671), .S(n10579), .Y(n9685) );
  MUX2X1 U10616 ( .B(ram[1636]), .A(ram[1572]), .S(n10706), .Y(n9679) );
  MUX2X1 U10617 ( .B(ram[1764]), .A(ram[1700]), .S(n10706), .Y(n9678) );
  MUX2X1 U10618 ( .B(ram[1892]), .A(ram[1828]), .S(n10706), .Y(n9682) );
  MUX2X1 U10619 ( .B(ram[2020]), .A(ram[1956]), .S(n10706), .Y(n9681) );
  MUX2X1 U10620 ( .B(n9680), .A(n9677), .S(n10579), .Y(n9684) );
  MUX2X1 U10621 ( .B(n9683), .A(n9668), .S(read2_addr[0]), .Y(n10532) );
  MUX2X1 U10622 ( .B(ram[101]), .A(ram[37]), .S(n10707), .Y(n9688) );
  MUX2X1 U10623 ( .B(ram[229]), .A(ram[165]), .S(n10707), .Y(n9687) );
  MUX2X1 U10624 ( .B(ram[357]), .A(ram[293]), .S(n10707), .Y(n9691) );
  MUX2X1 U10625 ( .B(ram[485]), .A(ram[421]), .S(n10707), .Y(n9690) );
  MUX2X1 U10626 ( .B(n9689), .A(n9686), .S(n10580), .Y(n9700) );
  MUX2X1 U10627 ( .B(ram[613]), .A(ram[549]), .S(n10707), .Y(n9694) );
  MUX2X1 U10628 ( .B(ram[741]), .A(ram[677]), .S(n10707), .Y(n9693) );
  MUX2X1 U10629 ( .B(ram[869]), .A(ram[805]), .S(n10707), .Y(n9697) );
  MUX2X1 U10630 ( .B(ram[997]), .A(ram[933]), .S(n10707), .Y(n9696) );
  MUX2X1 U10631 ( .B(n9695), .A(n9692), .S(n10580), .Y(n9699) );
  MUX2X1 U10632 ( .B(ram[1125]), .A(ram[1061]), .S(n10707), .Y(n9703) );
  MUX2X1 U10633 ( .B(ram[1253]), .A(ram[1189]), .S(n10707), .Y(n9702) );
  MUX2X1 U10634 ( .B(ram[1381]), .A(ram[1317]), .S(n10707), .Y(n9706) );
  MUX2X1 U10635 ( .B(ram[1509]), .A(ram[1445]), .S(n10707), .Y(n9705) );
  MUX2X1 U10636 ( .B(n9704), .A(n9701), .S(n10580), .Y(n9715) );
  MUX2X1 U10637 ( .B(ram[1637]), .A(ram[1573]), .S(n10708), .Y(n9709) );
  MUX2X1 U10638 ( .B(ram[1765]), .A(ram[1701]), .S(n10708), .Y(n9708) );
  MUX2X1 U10639 ( .B(ram[1893]), .A(ram[1829]), .S(n10708), .Y(n9712) );
  MUX2X1 U10640 ( .B(ram[2021]), .A(ram[1957]), .S(n10708), .Y(n9711) );
  MUX2X1 U10641 ( .B(n9710), .A(n9707), .S(n10580), .Y(n9714) );
  MUX2X1 U10642 ( .B(n9713), .A(n9698), .S(read2_addr[0]), .Y(n10533) );
  MUX2X1 U10643 ( .B(ram[102]), .A(ram[38]), .S(n10708), .Y(n9718) );
  MUX2X1 U10644 ( .B(ram[230]), .A(ram[166]), .S(n10708), .Y(n9717) );
  MUX2X1 U10645 ( .B(ram[358]), .A(ram[294]), .S(n10708), .Y(n9721) );
  MUX2X1 U10646 ( .B(ram[486]), .A(ram[422]), .S(n10708), .Y(n9720) );
  MUX2X1 U10647 ( .B(n9719), .A(n9716), .S(n10580), .Y(n9730) );
  MUX2X1 U10648 ( .B(ram[614]), .A(ram[550]), .S(n10708), .Y(n9724) );
  MUX2X1 U10649 ( .B(ram[742]), .A(ram[678]), .S(n10708), .Y(n9723) );
  MUX2X1 U10650 ( .B(ram[870]), .A(ram[806]), .S(n10708), .Y(n9727) );
  MUX2X1 U10651 ( .B(ram[998]), .A(ram[934]), .S(n10708), .Y(n9726) );
  MUX2X1 U10652 ( .B(n9725), .A(n9722), .S(n10580), .Y(n9729) );
  MUX2X1 U10653 ( .B(ram[1126]), .A(ram[1062]), .S(n10709), .Y(n9733) );
  MUX2X1 U10654 ( .B(ram[1254]), .A(ram[1190]), .S(n10709), .Y(n9732) );
  MUX2X1 U10655 ( .B(ram[1382]), .A(ram[1318]), .S(n10709), .Y(n9736) );
  MUX2X1 U10656 ( .B(ram[1510]), .A(ram[1446]), .S(n10709), .Y(n9735) );
  MUX2X1 U10657 ( .B(n9734), .A(n9731), .S(n10580), .Y(n9745) );
  MUX2X1 U10658 ( .B(ram[1638]), .A(ram[1574]), .S(n10709), .Y(n9739) );
  MUX2X1 U10659 ( .B(ram[1766]), .A(ram[1702]), .S(n10709), .Y(n9738) );
  MUX2X1 U10660 ( .B(ram[1894]), .A(ram[1830]), .S(n10709), .Y(n9742) );
  MUX2X1 U10661 ( .B(ram[2022]), .A(ram[1958]), .S(n10709), .Y(n9741) );
  MUX2X1 U10662 ( .B(n9740), .A(n9737), .S(n10580), .Y(n9744) );
  MUX2X1 U10663 ( .B(n9743), .A(n9728), .S(read2_addr[0]), .Y(n10534) );
  MUX2X1 U10664 ( .B(ram[103]), .A(ram[39]), .S(n10709), .Y(n9748) );
  MUX2X1 U10665 ( .B(ram[231]), .A(ram[167]), .S(n10709), .Y(n9747) );
  MUX2X1 U10666 ( .B(ram[359]), .A(ram[295]), .S(n10709), .Y(n9751) );
  MUX2X1 U10667 ( .B(ram[487]), .A(ram[423]), .S(n10709), .Y(n9750) );
  MUX2X1 U10668 ( .B(n9749), .A(n9746), .S(n10580), .Y(n9760) );
  MUX2X1 U10669 ( .B(ram[615]), .A(ram[551]), .S(n10710), .Y(n9754) );
  MUX2X1 U10670 ( .B(ram[743]), .A(ram[679]), .S(n10710), .Y(n9753) );
  MUX2X1 U10671 ( .B(ram[871]), .A(ram[807]), .S(n10710), .Y(n9757) );
  MUX2X1 U10672 ( .B(ram[999]), .A(ram[935]), .S(n10710), .Y(n9756) );
  MUX2X1 U10673 ( .B(n9755), .A(n9752), .S(n10580), .Y(n9759) );
  MUX2X1 U10674 ( .B(ram[1127]), .A(ram[1063]), .S(n10710), .Y(n9763) );
  MUX2X1 U10675 ( .B(ram[1255]), .A(ram[1191]), .S(n10710), .Y(n9762) );
  MUX2X1 U10676 ( .B(ram[1383]), .A(ram[1319]), .S(n10710), .Y(n9766) );
  MUX2X1 U10677 ( .B(ram[1511]), .A(ram[1447]), .S(n10710), .Y(n9765) );
  MUX2X1 U10678 ( .B(n9764), .A(n9761), .S(n10580), .Y(n9775) );
  MUX2X1 U10679 ( .B(ram[1639]), .A(ram[1575]), .S(n10710), .Y(n9769) );
  MUX2X1 U10680 ( .B(ram[1767]), .A(ram[1703]), .S(n10710), .Y(n9768) );
  MUX2X1 U10681 ( .B(ram[1895]), .A(ram[1831]), .S(n10710), .Y(n9772) );
  MUX2X1 U10682 ( .B(ram[2023]), .A(ram[1959]), .S(n10710), .Y(n9771) );
  MUX2X1 U10683 ( .B(n9770), .A(n9767), .S(n10580), .Y(n9774) );
  MUX2X1 U10684 ( .B(n9773), .A(n9758), .S(read2_addr[0]), .Y(n10535) );
  MUX2X1 U10685 ( .B(ram[104]), .A(ram[40]), .S(n10711), .Y(n9778) );
  MUX2X1 U10686 ( .B(ram[232]), .A(ram[168]), .S(n10711), .Y(n9777) );
  MUX2X1 U10687 ( .B(ram[360]), .A(ram[296]), .S(n10711), .Y(n9781) );
  MUX2X1 U10688 ( .B(ram[488]), .A(ram[424]), .S(n10711), .Y(n9780) );
  MUX2X1 U10689 ( .B(n9779), .A(n9776), .S(n10581), .Y(n9790) );
  MUX2X1 U10690 ( .B(ram[616]), .A(ram[552]), .S(n10711), .Y(n9784) );
  MUX2X1 U10691 ( .B(ram[744]), .A(ram[680]), .S(n10711), .Y(n9783) );
  MUX2X1 U10692 ( .B(ram[872]), .A(ram[808]), .S(n10711), .Y(n9787) );
  MUX2X1 U10693 ( .B(ram[1000]), .A(ram[936]), .S(n10711), .Y(n9786) );
  MUX2X1 U10694 ( .B(n9785), .A(n9782), .S(n10581), .Y(n9789) );
  MUX2X1 U10695 ( .B(ram[1128]), .A(ram[1064]), .S(n10711), .Y(n9793) );
  MUX2X1 U10696 ( .B(ram[1256]), .A(ram[1192]), .S(n10711), .Y(n9792) );
  MUX2X1 U10697 ( .B(ram[1384]), .A(ram[1320]), .S(n10711), .Y(n9796) );
  MUX2X1 U10698 ( .B(ram[1512]), .A(ram[1448]), .S(n10711), .Y(n9795) );
  MUX2X1 U10699 ( .B(n9794), .A(n9791), .S(n10581), .Y(n9805) );
  MUX2X1 U10700 ( .B(ram[1640]), .A(ram[1576]), .S(n10712), .Y(n9799) );
  MUX2X1 U10701 ( .B(ram[1768]), .A(ram[1704]), .S(n10712), .Y(n9798) );
  MUX2X1 U10702 ( .B(ram[1896]), .A(ram[1832]), .S(n10712), .Y(n9802) );
  MUX2X1 U10703 ( .B(ram[2024]), .A(ram[1960]), .S(n10712), .Y(n9801) );
  MUX2X1 U10704 ( .B(n9800), .A(n9797), .S(n10581), .Y(n9804) );
  MUX2X1 U10705 ( .B(n9803), .A(n9788), .S(read2_addr[0]), .Y(n10536) );
  MUX2X1 U10706 ( .B(ram[105]), .A(ram[41]), .S(n10712), .Y(n9808) );
  MUX2X1 U10707 ( .B(ram[233]), .A(ram[169]), .S(n10712), .Y(n9807) );
  MUX2X1 U10708 ( .B(ram[361]), .A(ram[297]), .S(n10712), .Y(n9811) );
  MUX2X1 U10709 ( .B(ram[489]), .A(ram[425]), .S(n10712), .Y(n9810) );
  MUX2X1 U10710 ( .B(n9809), .A(n9806), .S(n10581), .Y(n9820) );
  MUX2X1 U10711 ( .B(ram[617]), .A(ram[553]), .S(n10712), .Y(n9814) );
  MUX2X1 U10712 ( .B(ram[745]), .A(ram[681]), .S(n10712), .Y(n9813) );
  MUX2X1 U10713 ( .B(ram[873]), .A(ram[809]), .S(n10712), .Y(n9817) );
  MUX2X1 U10714 ( .B(ram[1001]), .A(ram[937]), .S(n10712), .Y(n9816) );
  MUX2X1 U10715 ( .B(n9815), .A(n9812), .S(n10581), .Y(n9819) );
  MUX2X1 U10716 ( .B(ram[1129]), .A(ram[1065]), .S(n10713), .Y(n9823) );
  MUX2X1 U10717 ( .B(ram[1257]), .A(ram[1193]), .S(n10713), .Y(n9822) );
  MUX2X1 U10718 ( .B(ram[1385]), .A(ram[1321]), .S(n10713), .Y(n9826) );
  MUX2X1 U10719 ( .B(ram[1513]), .A(ram[1449]), .S(n10713), .Y(n9825) );
  MUX2X1 U10720 ( .B(n9824), .A(n9821), .S(n10581), .Y(n9835) );
  MUX2X1 U10721 ( .B(ram[1641]), .A(ram[1577]), .S(n10713), .Y(n9829) );
  MUX2X1 U10722 ( .B(ram[1769]), .A(ram[1705]), .S(n10713), .Y(n9828) );
  MUX2X1 U10723 ( .B(ram[1897]), .A(ram[1833]), .S(n10713), .Y(n9832) );
  MUX2X1 U10724 ( .B(ram[2025]), .A(ram[1961]), .S(n10713), .Y(n9831) );
  MUX2X1 U10725 ( .B(n9830), .A(n9827), .S(n10581), .Y(n9834) );
  MUX2X1 U10726 ( .B(n9833), .A(n9818), .S(read2_addr[0]), .Y(n10537) );
  MUX2X1 U10727 ( .B(ram[106]), .A(ram[42]), .S(n10713), .Y(n9838) );
  MUX2X1 U10728 ( .B(ram[234]), .A(ram[170]), .S(n10713), .Y(n9837) );
  MUX2X1 U10729 ( .B(ram[362]), .A(ram[298]), .S(n10713), .Y(n9841) );
  MUX2X1 U10730 ( .B(ram[490]), .A(ram[426]), .S(n10713), .Y(n9840) );
  MUX2X1 U10731 ( .B(n9839), .A(n9836), .S(n10581), .Y(n9850) );
  MUX2X1 U10732 ( .B(ram[618]), .A(ram[554]), .S(n10714), .Y(n9844) );
  MUX2X1 U10733 ( .B(ram[746]), .A(ram[682]), .S(n10714), .Y(n9843) );
  MUX2X1 U10734 ( .B(ram[874]), .A(ram[810]), .S(n10714), .Y(n9847) );
  MUX2X1 U10735 ( .B(ram[1002]), .A(ram[938]), .S(n10714), .Y(n9846) );
  MUX2X1 U10736 ( .B(n9845), .A(n9842), .S(n10581), .Y(n9849) );
  MUX2X1 U10737 ( .B(ram[1130]), .A(ram[1066]), .S(n10714), .Y(n9853) );
  MUX2X1 U10738 ( .B(ram[1258]), .A(ram[1194]), .S(n10714), .Y(n9852) );
  MUX2X1 U10739 ( .B(ram[1386]), .A(ram[1322]), .S(n10714), .Y(n9856) );
  MUX2X1 U10740 ( .B(ram[1514]), .A(ram[1450]), .S(n10714), .Y(n9855) );
  MUX2X1 U10741 ( .B(n9854), .A(n9851), .S(n10581), .Y(n9865) );
  MUX2X1 U10742 ( .B(ram[1642]), .A(ram[1578]), .S(n10714), .Y(n9859) );
  MUX2X1 U10743 ( .B(ram[1770]), .A(ram[1706]), .S(n10714), .Y(n9858) );
  MUX2X1 U10744 ( .B(ram[1898]), .A(ram[1834]), .S(n10714), .Y(n9862) );
  MUX2X1 U10745 ( .B(ram[2026]), .A(ram[1962]), .S(n10714), .Y(n9861) );
  MUX2X1 U10746 ( .B(n9860), .A(n9857), .S(n10581), .Y(n9864) );
  MUX2X1 U10747 ( .B(n9863), .A(n9848), .S(read2_addr[0]), .Y(n10538) );
  MUX2X1 U10748 ( .B(ram[107]), .A(ram[43]), .S(n10715), .Y(n9868) );
  MUX2X1 U10749 ( .B(ram[235]), .A(ram[171]), .S(n10715), .Y(n9867) );
  MUX2X1 U10750 ( .B(ram[363]), .A(ram[299]), .S(n10715), .Y(n9871) );
  MUX2X1 U10751 ( .B(ram[491]), .A(ram[427]), .S(n10715), .Y(n9870) );
  MUX2X1 U10752 ( .B(n9869), .A(n9866), .S(n10582), .Y(n9880) );
  MUX2X1 U10753 ( .B(ram[619]), .A(ram[555]), .S(n10715), .Y(n9874) );
  MUX2X1 U10754 ( .B(ram[747]), .A(ram[683]), .S(n10715), .Y(n9873) );
  MUX2X1 U10755 ( .B(ram[875]), .A(ram[811]), .S(n10715), .Y(n9877) );
  MUX2X1 U10756 ( .B(ram[1003]), .A(ram[939]), .S(n10715), .Y(n9876) );
  MUX2X1 U10757 ( .B(n9875), .A(n9872), .S(n10582), .Y(n9879) );
  MUX2X1 U10758 ( .B(ram[1131]), .A(ram[1067]), .S(n10715), .Y(n9883) );
  MUX2X1 U10759 ( .B(ram[1259]), .A(ram[1195]), .S(n10715), .Y(n9882) );
  MUX2X1 U10760 ( .B(ram[1387]), .A(ram[1323]), .S(n10715), .Y(n9886) );
  MUX2X1 U10761 ( .B(ram[1515]), .A(ram[1451]), .S(n10715), .Y(n9885) );
  MUX2X1 U10762 ( .B(n9884), .A(n9881), .S(n10582), .Y(n9895) );
  MUX2X1 U10763 ( .B(ram[1643]), .A(ram[1579]), .S(n10716), .Y(n9889) );
  MUX2X1 U10764 ( .B(ram[1771]), .A(ram[1707]), .S(n10716), .Y(n9888) );
  MUX2X1 U10765 ( .B(ram[1899]), .A(ram[1835]), .S(n10716), .Y(n9892) );
  MUX2X1 U10766 ( .B(ram[2027]), .A(ram[1963]), .S(n10716), .Y(n9891) );
  MUX2X1 U10767 ( .B(n9890), .A(n9887), .S(n10582), .Y(n9894) );
  MUX2X1 U10768 ( .B(n9893), .A(n9878), .S(read2_addr[0]), .Y(n10539) );
  MUX2X1 U10769 ( .B(ram[108]), .A(ram[44]), .S(n10716), .Y(n9898) );
  MUX2X1 U10770 ( .B(ram[236]), .A(ram[172]), .S(n10716), .Y(n9897) );
  MUX2X1 U10771 ( .B(ram[364]), .A(ram[300]), .S(n10716), .Y(n9901) );
  MUX2X1 U10772 ( .B(ram[492]), .A(ram[428]), .S(n10716), .Y(n9900) );
  MUX2X1 U10773 ( .B(n9899), .A(n9896), .S(n10582), .Y(n9910) );
  MUX2X1 U10774 ( .B(ram[620]), .A(ram[556]), .S(n10716), .Y(n9904) );
  MUX2X1 U10775 ( .B(ram[748]), .A(ram[684]), .S(n10716), .Y(n9903) );
  MUX2X1 U10776 ( .B(ram[876]), .A(ram[812]), .S(n10716), .Y(n9907) );
  MUX2X1 U10777 ( .B(ram[1004]), .A(ram[940]), .S(n10716), .Y(n9906) );
  MUX2X1 U10778 ( .B(n9905), .A(n9902), .S(n10582), .Y(n9909) );
  MUX2X1 U10779 ( .B(ram[1132]), .A(ram[1068]), .S(n10717), .Y(n9913) );
  MUX2X1 U10780 ( .B(ram[1260]), .A(ram[1196]), .S(n10717), .Y(n9912) );
  MUX2X1 U10781 ( .B(ram[1388]), .A(ram[1324]), .S(n10717), .Y(n9916) );
  MUX2X1 U10782 ( .B(ram[1516]), .A(ram[1452]), .S(n10717), .Y(n9915) );
  MUX2X1 U10783 ( .B(n9914), .A(n9911), .S(n10582), .Y(n9925) );
  MUX2X1 U10784 ( .B(ram[1644]), .A(ram[1580]), .S(n10717), .Y(n9919) );
  MUX2X1 U10785 ( .B(ram[1772]), .A(ram[1708]), .S(n10717), .Y(n9918) );
  MUX2X1 U10786 ( .B(ram[1900]), .A(ram[1836]), .S(n10717), .Y(n9922) );
  MUX2X1 U10787 ( .B(ram[2028]), .A(ram[1964]), .S(n10717), .Y(n9921) );
  MUX2X1 U10788 ( .B(n9920), .A(n9917), .S(n10582), .Y(n9924) );
  MUX2X1 U10789 ( .B(n9923), .A(n9908), .S(read2_addr[0]), .Y(n10540) );
  MUX2X1 U10790 ( .B(ram[109]), .A(ram[45]), .S(n10717), .Y(n9928) );
  MUX2X1 U10791 ( .B(ram[237]), .A(ram[173]), .S(n10717), .Y(n9927) );
  MUX2X1 U10792 ( .B(ram[365]), .A(ram[301]), .S(n10717), .Y(n9931) );
  MUX2X1 U10793 ( .B(ram[493]), .A(ram[429]), .S(n10717), .Y(n9930) );
  MUX2X1 U10794 ( .B(n9929), .A(n9926), .S(n10582), .Y(n9940) );
  MUX2X1 U10795 ( .B(ram[621]), .A(ram[557]), .S(n10718), .Y(n9934) );
  MUX2X1 U10796 ( .B(ram[749]), .A(ram[685]), .S(n10718), .Y(n9933) );
  MUX2X1 U10797 ( .B(ram[877]), .A(ram[813]), .S(n10718), .Y(n9937) );
  MUX2X1 U10798 ( .B(ram[1005]), .A(ram[941]), .S(n10718), .Y(n9936) );
  MUX2X1 U10799 ( .B(n9935), .A(n9932), .S(n10582), .Y(n9939) );
  MUX2X1 U10800 ( .B(ram[1133]), .A(ram[1069]), .S(n10718), .Y(n9943) );
  MUX2X1 U10801 ( .B(ram[1261]), .A(ram[1197]), .S(n10718), .Y(n9942) );
  MUX2X1 U10802 ( .B(ram[1389]), .A(ram[1325]), .S(n10718), .Y(n9946) );
  MUX2X1 U10803 ( .B(ram[1517]), .A(ram[1453]), .S(n10718), .Y(n9945) );
  MUX2X1 U10804 ( .B(n9944), .A(n9941), .S(n10582), .Y(n9955) );
  MUX2X1 U10805 ( .B(ram[1645]), .A(ram[1581]), .S(n10718), .Y(n9949) );
  MUX2X1 U10806 ( .B(ram[1773]), .A(ram[1709]), .S(n10718), .Y(n9948) );
  MUX2X1 U10807 ( .B(ram[1901]), .A(ram[1837]), .S(n10718), .Y(n9952) );
  MUX2X1 U10808 ( .B(ram[2029]), .A(ram[1965]), .S(n10718), .Y(n9951) );
  MUX2X1 U10809 ( .B(n9950), .A(n9947), .S(n10582), .Y(n9954) );
  MUX2X1 U10810 ( .B(n9953), .A(n9938), .S(read2_addr[0]), .Y(n10541) );
  MUX2X1 U10811 ( .B(ram[110]), .A(ram[46]), .S(n10719), .Y(n9958) );
  MUX2X1 U10812 ( .B(ram[238]), .A(ram[174]), .S(n10719), .Y(n9957) );
  MUX2X1 U10813 ( .B(ram[366]), .A(ram[302]), .S(n10719), .Y(n9961) );
  MUX2X1 U10814 ( .B(ram[494]), .A(ram[430]), .S(n10719), .Y(n9960) );
  MUX2X1 U10815 ( .B(n9959), .A(n9956), .S(n10583), .Y(n9970) );
  MUX2X1 U10816 ( .B(ram[622]), .A(ram[558]), .S(n10719), .Y(n9964) );
  MUX2X1 U10817 ( .B(ram[750]), .A(ram[686]), .S(n10719), .Y(n9963) );
  MUX2X1 U10818 ( .B(ram[878]), .A(ram[814]), .S(n10719), .Y(n9967) );
  MUX2X1 U10819 ( .B(ram[1006]), .A(ram[942]), .S(n10719), .Y(n9966) );
  MUX2X1 U10820 ( .B(n9965), .A(n9962), .S(n10583), .Y(n9969) );
  MUX2X1 U10821 ( .B(ram[1134]), .A(ram[1070]), .S(n10719), .Y(n9973) );
  MUX2X1 U10822 ( .B(ram[1262]), .A(ram[1198]), .S(n10719), .Y(n9972) );
  MUX2X1 U10823 ( .B(ram[1390]), .A(ram[1326]), .S(n10719), .Y(n9976) );
  MUX2X1 U10824 ( .B(ram[1518]), .A(ram[1454]), .S(n10719), .Y(n9975) );
  MUX2X1 U10825 ( .B(n9974), .A(n9971), .S(n10583), .Y(n9985) );
  MUX2X1 U10826 ( .B(ram[1646]), .A(ram[1582]), .S(n10720), .Y(n9979) );
  MUX2X1 U10827 ( .B(ram[1774]), .A(ram[1710]), .S(n10720), .Y(n9978) );
  MUX2X1 U10828 ( .B(ram[1902]), .A(ram[1838]), .S(n10720), .Y(n9982) );
  MUX2X1 U10829 ( .B(ram[2030]), .A(ram[1966]), .S(n10720), .Y(n9981) );
  MUX2X1 U10830 ( .B(n9980), .A(n9977), .S(n10583), .Y(n9984) );
  MUX2X1 U10831 ( .B(n9983), .A(n9968), .S(read2_addr[0]), .Y(n10542) );
  MUX2X1 U10832 ( .B(ram[111]), .A(ram[47]), .S(n10720), .Y(n9988) );
  MUX2X1 U10833 ( .B(ram[239]), .A(ram[175]), .S(n10720), .Y(n9987) );
  MUX2X1 U10834 ( .B(ram[367]), .A(ram[303]), .S(n10720), .Y(n9991) );
  MUX2X1 U10835 ( .B(ram[495]), .A(ram[431]), .S(n10720), .Y(n9990) );
  MUX2X1 U10836 ( .B(n9989), .A(n9986), .S(n10583), .Y(n10000) );
  MUX2X1 U10837 ( .B(ram[623]), .A(ram[559]), .S(n10720), .Y(n9994) );
  MUX2X1 U10838 ( .B(ram[751]), .A(ram[687]), .S(n10720), .Y(n9993) );
  MUX2X1 U10839 ( .B(ram[879]), .A(ram[815]), .S(n10720), .Y(n9997) );
  MUX2X1 U10840 ( .B(ram[1007]), .A(ram[943]), .S(n10720), .Y(n9996) );
  MUX2X1 U10841 ( .B(n9995), .A(n9992), .S(n10583), .Y(n9999) );
  MUX2X1 U10842 ( .B(ram[1135]), .A(ram[1071]), .S(n10721), .Y(n10003) );
  MUX2X1 U10843 ( .B(ram[1263]), .A(ram[1199]), .S(n10721), .Y(n10002) );
  MUX2X1 U10844 ( .B(ram[1391]), .A(ram[1327]), .S(n10721), .Y(n10006) );
  MUX2X1 U10845 ( .B(ram[1519]), .A(ram[1455]), .S(n10721), .Y(n10005) );
  MUX2X1 U10846 ( .B(n10004), .A(n10001), .S(n10583), .Y(n10015) );
  MUX2X1 U10847 ( .B(ram[1647]), .A(ram[1583]), .S(n10721), .Y(n10009) );
  MUX2X1 U10848 ( .B(ram[1775]), .A(ram[1711]), .S(n10721), .Y(n10008) );
  MUX2X1 U10849 ( .B(ram[1903]), .A(ram[1839]), .S(n10721), .Y(n10012) );
  MUX2X1 U10850 ( .B(ram[2031]), .A(ram[1967]), .S(n10721), .Y(n10011) );
  MUX2X1 U10851 ( .B(n10010), .A(n10007), .S(n10583), .Y(n10014) );
  MUX2X1 U10852 ( .B(n10013), .A(n9998), .S(n10561), .Y(n10543) );
  MUX2X1 U10853 ( .B(ram[112]), .A(ram[48]), .S(n10721), .Y(n10018) );
  MUX2X1 U10854 ( .B(ram[240]), .A(ram[176]), .S(n10721), .Y(n10017) );
  MUX2X1 U10855 ( .B(ram[368]), .A(ram[304]), .S(n10721), .Y(n10021) );
  MUX2X1 U10856 ( .B(ram[496]), .A(ram[432]), .S(n10721), .Y(n10020) );
  MUX2X1 U10857 ( .B(n10019), .A(n10016), .S(n10583), .Y(n10030) );
  MUX2X1 U10858 ( .B(ram[624]), .A(ram[560]), .S(n10722), .Y(n10024) );
  MUX2X1 U10859 ( .B(ram[752]), .A(ram[688]), .S(n10722), .Y(n10023) );
  MUX2X1 U10860 ( .B(ram[880]), .A(ram[816]), .S(n10722), .Y(n10027) );
  MUX2X1 U10861 ( .B(ram[1008]), .A(ram[944]), .S(n10722), .Y(n10026) );
  MUX2X1 U10862 ( .B(n10025), .A(n10022), .S(n10583), .Y(n10029) );
  MUX2X1 U10863 ( .B(ram[1136]), .A(ram[1072]), .S(n10722), .Y(n10033) );
  MUX2X1 U10864 ( .B(ram[1264]), .A(ram[1200]), .S(n10722), .Y(n10032) );
  MUX2X1 U10865 ( .B(ram[1392]), .A(ram[1328]), .S(n10722), .Y(n10036) );
  MUX2X1 U10866 ( .B(ram[1520]), .A(ram[1456]), .S(n10722), .Y(n10035) );
  MUX2X1 U10867 ( .B(n10034), .A(n10031), .S(n10583), .Y(n10045) );
  MUX2X1 U10868 ( .B(ram[1648]), .A(ram[1584]), .S(n10722), .Y(n10039) );
  MUX2X1 U10869 ( .B(ram[1776]), .A(ram[1712]), .S(n10722), .Y(n10038) );
  MUX2X1 U10870 ( .B(ram[1904]), .A(ram[1840]), .S(n10722), .Y(n10042) );
  MUX2X1 U10871 ( .B(ram[2032]), .A(ram[1968]), .S(n10722), .Y(n10041) );
  MUX2X1 U10872 ( .B(n10040), .A(n10037), .S(n10583), .Y(n10044) );
  MUX2X1 U10873 ( .B(n10043), .A(n10028), .S(n10562), .Y(n10544) );
  MUX2X1 U10874 ( .B(ram[113]), .A(ram[49]), .S(n10723), .Y(n10048) );
  MUX2X1 U10875 ( .B(ram[241]), .A(ram[177]), .S(n10723), .Y(n10047) );
  MUX2X1 U10876 ( .B(ram[369]), .A(ram[305]), .S(n10723), .Y(n10051) );
  MUX2X1 U10877 ( .B(ram[497]), .A(ram[433]), .S(n10723), .Y(n10050) );
  MUX2X1 U10878 ( .B(n10049), .A(n10046), .S(n10569), .Y(n10060) );
  MUX2X1 U10879 ( .B(ram[625]), .A(ram[561]), .S(n10723), .Y(n10054) );
  MUX2X1 U10880 ( .B(ram[753]), .A(ram[689]), .S(n10723), .Y(n10053) );
  MUX2X1 U10881 ( .B(ram[881]), .A(ram[817]), .S(n10723), .Y(n10057) );
  MUX2X1 U10882 ( .B(ram[1009]), .A(ram[945]), .S(n10723), .Y(n10056) );
  MUX2X1 U10883 ( .B(n10055), .A(n10052), .S(n10578), .Y(n10059) );
  MUX2X1 U10884 ( .B(ram[1137]), .A(ram[1073]), .S(n10723), .Y(n10063) );
  MUX2X1 U10885 ( .B(ram[1265]), .A(ram[1201]), .S(n10723), .Y(n10062) );
  MUX2X1 U10886 ( .B(ram[1393]), .A(ram[1329]), .S(n10723), .Y(n10066) );
  MUX2X1 U10887 ( .B(ram[1521]), .A(ram[1457]), .S(n10723), .Y(n10065) );
  MUX2X1 U10888 ( .B(n10064), .A(n10061), .S(n10570), .Y(n10075) );
  MUX2X1 U10889 ( .B(ram[1649]), .A(ram[1585]), .S(n10724), .Y(n10069) );
  MUX2X1 U10890 ( .B(ram[1777]), .A(ram[1713]), .S(n10724), .Y(n10068) );
  MUX2X1 U10891 ( .B(ram[1905]), .A(ram[1841]), .S(n10724), .Y(n10072) );
  MUX2X1 U10892 ( .B(ram[2033]), .A(ram[1969]), .S(n10724), .Y(n10071) );
  MUX2X1 U10893 ( .B(n10070), .A(n10067), .S(n10583), .Y(n10074) );
  MUX2X1 U10894 ( .B(n10073), .A(n10058), .S(n10561), .Y(n10545) );
  MUX2X1 U10895 ( .B(ram[114]), .A(ram[50]), .S(n10724), .Y(n10078) );
  MUX2X1 U10896 ( .B(ram[242]), .A(ram[178]), .S(n10724), .Y(n10077) );
  MUX2X1 U10897 ( .B(ram[370]), .A(ram[306]), .S(n10724), .Y(n10081) );
  MUX2X1 U10898 ( .B(ram[498]), .A(ram[434]), .S(n10724), .Y(n10080) );
  MUX2X1 U10899 ( .B(n10079), .A(n10076), .S(n10575), .Y(n10090) );
  MUX2X1 U10900 ( .B(ram[626]), .A(ram[562]), .S(n10724), .Y(n10084) );
  MUX2X1 U10901 ( .B(ram[754]), .A(ram[690]), .S(n10724), .Y(n10083) );
  MUX2X1 U10902 ( .B(ram[882]), .A(ram[818]), .S(n10724), .Y(n10087) );
  MUX2X1 U10903 ( .B(ram[1010]), .A(ram[946]), .S(n10724), .Y(n10086) );
  MUX2X1 U10904 ( .B(n10085), .A(n10082), .S(n10582), .Y(n10089) );
  MUX2X1 U10905 ( .B(ram[1138]), .A(ram[1074]), .S(n10725), .Y(n10093) );
  MUX2X1 U10906 ( .B(ram[1266]), .A(ram[1202]), .S(n10725), .Y(n10092) );
  MUX2X1 U10907 ( .B(ram[1394]), .A(ram[1330]), .S(n10725), .Y(n10096) );
  MUX2X1 U10908 ( .B(ram[1522]), .A(ram[1458]), .S(n10725), .Y(n10095) );
  MUX2X1 U10909 ( .B(n10094), .A(n10091), .S(n10580), .Y(n10105) );
  MUX2X1 U10910 ( .B(ram[1650]), .A(ram[1586]), .S(n10725), .Y(n10099) );
  MUX2X1 U10911 ( .B(ram[1778]), .A(ram[1714]), .S(n10725), .Y(n10098) );
  MUX2X1 U10912 ( .B(ram[1906]), .A(ram[1842]), .S(n10725), .Y(n10102) );
  MUX2X1 U10913 ( .B(ram[2034]), .A(ram[1970]), .S(n10725), .Y(n10101) );
  MUX2X1 U10914 ( .B(n10100), .A(n10097), .S(n10574), .Y(n10104) );
  MUX2X1 U10915 ( .B(n10103), .A(n10088), .S(read2_addr[0]), .Y(n10546) );
  MUX2X1 U10916 ( .B(ram[115]), .A(ram[51]), .S(n10725), .Y(n10108) );
  MUX2X1 U10917 ( .B(ram[243]), .A(ram[179]), .S(n10725), .Y(n10107) );
  MUX2X1 U10918 ( .B(ram[371]), .A(ram[307]), .S(n10725), .Y(n10111) );
  MUX2X1 U10919 ( .B(ram[499]), .A(ram[435]), .S(n10725), .Y(n10110) );
  MUX2X1 U10920 ( .B(n10109), .A(n10106), .S(n10571), .Y(n10120) );
  MUX2X1 U10921 ( .B(ram[627]), .A(ram[563]), .S(n10726), .Y(n10114) );
  MUX2X1 U10922 ( .B(ram[755]), .A(ram[691]), .S(n10726), .Y(n10113) );
  MUX2X1 U10923 ( .B(ram[883]), .A(ram[819]), .S(n10726), .Y(n10117) );
  MUX2X1 U10924 ( .B(ram[1011]), .A(ram[947]), .S(n10726), .Y(n10116) );
  MUX2X1 U10925 ( .B(n10115), .A(n10112), .S(n10579), .Y(n10119) );
  MUX2X1 U10926 ( .B(ram[1139]), .A(ram[1075]), .S(n10726), .Y(n10123) );
  MUX2X1 U10927 ( .B(ram[1267]), .A(ram[1203]), .S(n10726), .Y(n10122) );
  MUX2X1 U10928 ( .B(ram[1395]), .A(ram[1331]), .S(n10726), .Y(n10126) );
  MUX2X1 U10929 ( .B(ram[1523]), .A(ram[1459]), .S(n10726), .Y(n10125) );
  MUX2X1 U10930 ( .B(n10124), .A(n10121), .S(n10572), .Y(n10135) );
  MUX2X1 U10931 ( .B(ram[1651]), .A(ram[1587]), .S(n10726), .Y(n10129) );
  MUX2X1 U10932 ( .B(ram[1779]), .A(ram[1715]), .S(n10726), .Y(n10128) );
  MUX2X1 U10933 ( .B(ram[1907]), .A(ram[1843]), .S(n10726), .Y(n10132) );
  MUX2X1 U10934 ( .B(ram[2035]), .A(ram[1971]), .S(n10726), .Y(n10131) );
  MUX2X1 U10935 ( .B(n10130), .A(n10127), .S(n10577), .Y(n10134) );
  MUX2X1 U10936 ( .B(n10133), .A(n10118), .S(n10562), .Y(n10547) );
  MUX2X1 U10937 ( .B(ram[116]), .A(ram[52]), .S(n10727), .Y(n10138) );
  MUX2X1 U10938 ( .B(ram[244]), .A(ram[180]), .S(n10727), .Y(n10137) );
  MUX2X1 U10939 ( .B(ram[372]), .A(ram[308]), .S(n10727), .Y(n10141) );
  MUX2X1 U10940 ( .B(ram[500]), .A(ram[436]), .S(n10727), .Y(n10140) );
  MUX2X1 U10941 ( .B(n10139), .A(n10136), .S(n10583), .Y(n10150) );
  MUX2X1 U10942 ( .B(ram[628]), .A(ram[564]), .S(n10727), .Y(n10144) );
  MUX2X1 U10943 ( .B(ram[756]), .A(ram[692]), .S(n10727), .Y(n10143) );
  MUX2X1 U10944 ( .B(ram[884]), .A(ram[820]), .S(n10727), .Y(n10147) );
  MUX2X1 U10945 ( .B(ram[1012]), .A(ram[948]), .S(n10727), .Y(n10146) );
  MUX2X1 U10946 ( .B(n10145), .A(n10142), .S(n10576), .Y(n10149) );
  MUX2X1 U10947 ( .B(ram[1140]), .A(ram[1076]), .S(n10727), .Y(n10153) );
  MUX2X1 U10948 ( .B(ram[1268]), .A(ram[1204]), .S(n10727), .Y(n10152) );
  MUX2X1 U10949 ( .B(ram[1396]), .A(ram[1332]), .S(n10727), .Y(n10156) );
  MUX2X1 U10950 ( .B(ram[1524]), .A(ram[1460]), .S(n10727), .Y(n10155) );
  MUX2X1 U10951 ( .B(n10154), .A(n10151), .S(n10572), .Y(n10165) );
  MUX2X1 U10952 ( .B(ram[1652]), .A(ram[1588]), .S(n10728), .Y(n10159) );
  MUX2X1 U10953 ( .B(ram[1780]), .A(ram[1716]), .S(n10728), .Y(n10158) );
  MUX2X1 U10954 ( .B(ram[1908]), .A(ram[1844]), .S(n10728), .Y(n10162) );
  MUX2X1 U10955 ( .B(ram[2036]), .A(ram[1972]), .S(n10728), .Y(n10161) );
  MUX2X1 U10956 ( .B(n10160), .A(n10157), .S(n10577), .Y(n10164) );
  MUX2X1 U10957 ( .B(n10163), .A(n10148), .S(n10562), .Y(n10548) );
  MUX2X1 U10958 ( .B(ram[117]), .A(ram[53]), .S(n10728), .Y(n10168) );
  MUX2X1 U10959 ( .B(ram[245]), .A(ram[181]), .S(n10728), .Y(n10167) );
  MUX2X1 U10960 ( .B(ram[373]), .A(ram[309]), .S(n10728), .Y(n10171) );
  MUX2X1 U10961 ( .B(ram[501]), .A(ram[437]), .S(n10728), .Y(n10170) );
  MUX2X1 U10962 ( .B(n10169), .A(n10166), .S(n10580), .Y(n10180) );
  MUX2X1 U10963 ( .B(ram[629]), .A(ram[565]), .S(n10728), .Y(n10174) );
  MUX2X1 U10964 ( .B(ram[757]), .A(ram[693]), .S(n10728), .Y(n10173) );
  MUX2X1 U10965 ( .B(ram[885]), .A(ram[821]), .S(n10728), .Y(n10177) );
  MUX2X1 U10966 ( .B(ram[1013]), .A(ram[949]), .S(n10728), .Y(n10176) );
  MUX2X1 U10967 ( .B(n10175), .A(n10172), .S(n10570), .Y(n10179) );
  MUX2X1 U10968 ( .B(ram[1141]), .A(ram[1077]), .S(n10729), .Y(n10183) );
  MUX2X1 U10969 ( .B(ram[1269]), .A(ram[1205]), .S(n10729), .Y(n10182) );
  MUX2X1 U10970 ( .B(ram[1397]), .A(ram[1333]), .S(n10729), .Y(n10186) );
  MUX2X1 U10971 ( .B(ram[1525]), .A(ram[1461]), .S(n10729), .Y(n10185) );
  MUX2X1 U10972 ( .B(n10184), .A(n10181), .S(n10571), .Y(n10195) );
  MUX2X1 U10973 ( .B(ram[1653]), .A(ram[1589]), .S(n10729), .Y(n10189) );
  MUX2X1 U10974 ( .B(ram[1781]), .A(ram[1717]), .S(n10729), .Y(n10188) );
  MUX2X1 U10975 ( .B(ram[1909]), .A(ram[1845]), .S(n10729), .Y(n10192) );
  MUX2X1 U10976 ( .B(ram[2037]), .A(ram[1973]), .S(n10729), .Y(n10191) );
  MUX2X1 U10977 ( .B(n10190), .A(n10187), .S(n10574), .Y(n10194) );
  MUX2X1 U10978 ( .B(n10193), .A(n10178), .S(n10561), .Y(n10549) );
  MUX2X1 U10979 ( .B(ram[118]), .A(ram[54]), .S(n10729), .Y(n10198) );
  MUX2X1 U10980 ( .B(ram[246]), .A(ram[182]), .S(n10729), .Y(n10197) );
  MUX2X1 U10981 ( .B(ram[374]), .A(ram[310]), .S(n10729), .Y(n10201) );
  MUX2X1 U10982 ( .B(ram[502]), .A(ram[438]), .S(n10729), .Y(n10200) );
  MUX2X1 U10983 ( .B(n10199), .A(n10196), .S(n10568), .Y(n10210) );
  MUX2X1 U10984 ( .B(ram[630]), .A(ram[566]), .S(n10730), .Y(n10204) );
  MUX2X1 U10985 ( .B(ram[758]), .A(ram[694]), .S(n10730), .Y(n10203) );
  MUX2X1 U10986 ( .B(ram[886]), .A(ram[822]), .S(n10730), .Y(n10207) );
  MUX2X1 U10987 ( .B(ram[1014]), .A(ram[950]), .S(n10730), .Y(n10206) );
  MUX2X1 U10988 ( .B(n10205), .A(n10202), .S(n10573), .Y(n10209) );
  MUX2X1 U10989 ( .B(ram[1142]), .A(ram[1078]), .S(n10730), .Y(n10213) );
  MUX2X1 U10990 ( .B(ram[1270]), .A(ram[1206]), .S(n10730), .Y(n10212) );
  MUX2X1 U10991 ( .B(ram[1398]), .A(ram[1334]), .S(n10730), .Y(n10216) );
  MUX2X1 U10992 ( .B(ram[1526]), .A(ram[1462]), .S(n10730), .Y(n10215) );
  MUX2X1 U10993 ( .B(n10214), .A(n10211), .S(n10573), .Y(n10225) );
  MUX2X1 U10994 ( .B(ram[1654]), .A(ram[1590]), .S(n10730), .Y(n10219) );
  MUX2X1 U10995 ( .B(ram[1782]), .A(ram[1718]), .S(n10730), .Y(n10218) );
  MUX2X1 U10996 ( .B(ram[1910]), .A(ram[1846]), .S(n10730), .Y(n10222) );
  MUX2X1 U10997 ( .B(ram[2038]), .A(ram[1974]), .S(n10730), .Y(n10221) );
  MUX2X1 U10998 ( .B(n10220), .A(n10217), .S(n10579), .Y(n10224) );
  MUX2X1 U10999 ( .B(n10223), .A(n10208), .S(read2_addr[0]), .Y(n10550) );
  MUX2X1 U11000 ( .B(ram[119]), .A(ram[55]), .S(n10731), .Y(n10228) );
  MUX2X1 U11001 ( .B(ram[247]), .A(ram[183]), .S(n10731), .Y(n10227) );
  MUX2X1 U11002 ( .B(ram[375]), .A(ram[311]), .S(n10731), .Y(n10231) );
  MUX2X1 U11003 ( .B(ram[503]), .A(ram[439]), .S(n10731), .Y(n10230) );
  MUX2X1 U11004 ( .B(n10229), .A(n10226), .S(n10578), .Y(n10240) );
  MUX2X1 U11005 ( .B(ram[631]), .A(ram[567]), .S(n10731), .Y(n10234) );
  MUX2X1 U11006 ( .B(ram[759]), .A(ram[695]), .S(n10731), .Y(n10233) );
  MUX2X1 U11007 ( .B(ram[887]), .A(ram[823]), .S(n10731), .Y(n10237) );
  MUX2X1 U11008 ( .B(ram[1015]), .A(ram[951]), .S(n10731), .Y(n10236) );
  MUX2X1 U11009 ( .B(n10235), .A(n10232), .S(n10581), .Y(n10239) );
  MUX2X1 U11010 ( .B(ram[1143]), .A(ram[1079]), .S(n10731), .Y(n10243) );
  MUX2X1 U11011 ( .B(ram[1271]), .A(ram[1207]), .S(n10731), .Y(n10242) );
  MUX2X1 U11012 ( .B(ram[1399]), .A(ram[1335]), .S(n10731), .Y(n10246) );
  MUX2X1 U11013 ( .B(ram[1527]), .A(ram[1463]), .S(n10731), .Y(n10245) );
  MUX2X1 U11014 ( .B(n10244), .A(n10241), .S(n10568), .Y(n10255) );
  MUX2X1 U11015 ( .B(ram[1655]), .A(ram[1591]), .S(n10732), .Y(n10249) );
  MUX2X1 U11016 ( .B(ram[1783]), .A(ram[1719]), .S(n10732), .Y(n10248) );
  MUX2X1 U11017 ( .B(ram[1911]), .A(ram[1847]), .S(n10732), .Y(n10252) );
  MUX2X1 U11018 ( .B(ram[2039]), .A(ram[1975]), .S(n10732), .Y(n10251) );
  MUX2X1 U11019 ( .B(n10250), .A(n10247), .S(n10578), .Y(n10254) );
  MUX2X1 U11020 ( .B(n10253), .A(n10238), .S(n10561), .Y(n10551) );
  MUX2X1 U11021 ( .B(ram[120]), .A(ram[56]), .S(n10732), .Y(n10258) );
  MUX2X1 U11022 ( .B(ram[248]), .A(ram[184]), .S(n10732), .Y(n10257) );
  MUX2X1 U11023 ( .B(ram[376]), .A(ram[312]), .S(n10732), .Y(n10261) );
  MUX2X1 U11024 ( .B(ram[504]), .A(ram[440]), .S(n10732), .Y(n10260) );
  MUX2X1 U11025 ( .B(n10259), .A(n10256), .S(n10581), .Y(n10270) );
  MUX2X1 U11026 ( .B(ram[632]), .A(ram[568]), .S(n10732), .Y(n10264) );
  MUX2X1 U11027 ( .B(ram[760]), .A(ram[696]), .S(n10732), .Y(n10263) );
  MUX2X1 U11028 ( .B(ram[888]), .A(ram[824]), .S(n10732), .Y(n10267) );
  MUX2X1 U11029 ( .B(ram[1016]), .A(ram[952]), .S(n10732), .Y(n10266) );
  MUX2X1 U11030 ( .B(n10265), .A(n10262), .S(n10581), .Y(n10269) );
  MUX2X1 U11031 ( .B(ram[1144]), .A(ram[1080]), .S(n10733), .Y(n10273) );
  MUX2X1 U11032 ( .B(ram[1272]), .A(ram[1208]), .S(n10733), .Y(n10272) );
  MUX2X1 U11033 ( .B(ram[1400]), .A(ram[1336]), .S(n10733), .Y(n10276) );
  MUX2X1 U11034 ( .B(ram[1528]), .A(ram[1464]), .S(n10733), .Y(n10275) );
  MUX2X1 U11035 ( .B(n10274), .A(n10271), .S(n10568), .Y(n10285) );
  MUX2X1 U11036 ( .B(ram[1656]), .A(ram[1592]), .S(n10733), .Y(n10279) );
  MUX2X1 U11037 ( .B(ram[1784]), .A(ram[1720]), .S(n10733), .Y(n10278) );
  MUX2X1 U11038 ( .B(ram[1912]), .A(ram[1848]), .S(n10733), .Y(n10282) );
  MUX2X1 U11039 ( .B(ram[2040]), .A(ram[1976]), .S(n10733), .Y(n10281) );
  MUX2X1 U11040 ( .B(n10280), .A(n10277), .S(n10577), .Y(n10284) );
  MUX2X1 U11041 ( .B(n10283), .A(n10268), .S(n10562), .Y(n10552) );
  MUX2X1 U11042 ( .B(ram[121]), .A(ram[57]), .S(n10733), .Y(n10288) );
  MUX2X1 U11043 ( .B(ram[249]), .A(ram[185]), .S(n10733), .Y(n10287) );
  MUX2X1 U11044 ( .B(ram[377]), .A(ram[313]), .S(n10733), .Y(n10291) );
  MUX2X1 U11045 ( .B(ram[505]), .A(ram[441]), .S(n10733), .Y(n10290) );
  MUX2X1 U11046 ( .B(n10289), .A(n10286), .S(n10568), .Y(n10300) );
  MUX2X1 U11047 ( .B(ram[633]), .A(ram[569]), .S(n10734), .Y(n10294) );
  MUX2X1 U11048 ( .B(ram[761]), .A(ram[697]), .S(n10734), .Y(n10293) );
  MUX2X1 U11049 ( .B(ram[889]), .A(ram[825]), .S(n10734), .Y(n10297) );
  MUX2X1 U11050 ( .B(ram[1017]), .A(ram[953]), .S(n10734), .Y(n10296) );
  MUX2X1 U11051 ( .B(n10295), .A(n10292), .S(n10583), .Y(n10299) );
  MUX2X1 U11052 ( .B(ram[1145]), .A(ram[1081]), .S(n10734), .Y(n10303) );
  MUX2X1 U11053 ( .B(ram[1273]), .A(ram[1209]), .S(n10734), .Y(n10302) );
  MUX2X1 U11054 ( .B(ram[1401]), .A(ram[1337]), .S(n10734), .Y(n10306) );
  MUX2X1 U11055 ( .B(ram[1529]), .A(ram[1465]), .S(n10734), .Y(n10305) );
  MUX2X1 U11056 ( .B(n10304), .A(n10301), .S(n10583), .Y(n10315) );
  MUX2X1 U11057 ( .B(ram[1657]), .A(ram[1593]), .S(n10734), .Y(n10309) );
  MUX2X1 U11058 ( .B(ram[1785]), .A(ram[1721]), .S(n10734), .Y(n10308) );
  MUX2X1 U11059 ( .B(ram[1913]), .A(ram[1849]), .S(n10734), .Y(n10312) );
  MUX2X1 U11060 ( .B(ram[2041]), .A(ram[1977]), .S(n10734), .Y(n10311) );
  MUX2X1 U11061 ( .B(n10310), .A(n10307), .S(n10575), .Y(n10314) );
  MUX2X1 U11062 ( .B(n10313), .A(n10298), .S(n10561), .Y(n10553) );
  MUX2X1 U11063 ( .B(ram[122]), .A(ram[58]), .S(n10735), .Y(n10318) );
  MUX2X1 U11064 ( .B(ram[250]), .A(ram[186]), .S(n10735), .Y(n10317) );
  MUX2X1 U11065 ( .B(ram[378]), .A(ram[314]), .S(n10735), .Y(n10321) );
  MUX2X1 U11066 ( .B(ram[506]), .A(ram[442]), .S(n10735), .Y(n10320) );
  MUX2X1 U11067 ( .B(n10319), .A(n10316), .S(n10576), .Y(n10330) );
  MUX2X1 U11068 ( .B(ram[634]), .A(ram[570]), .S(n10735), .Y(n10324) );
  MUX2X1 U11069 ( .B(ram[762]), .A(ram[698]), .S(n10735), .Y(n10323) );
  MUX2X1 U11070 ( .B(ram[890]), .A(ram[826]), .S(n10735), .Y(n10327) );
  MUX2X1 U11071 ( .B(ram[1018]), .A(ram[954]), .S(n10735), .Y(n10326) );
  MUX2X1 U11072 ( .B(n10325), .A(n10322), .S(n10582), .Y(n10329) );
  MUX2X1 U11073 ( .B(ram[1146]), .A(ram[1082]), .S(n10735), .Y(n10333) );
  MUX2X1 U11074 ( .B(ram[1274]), .A(ram[1210]), .S(n10735), .Y(n10332) );
  MUX2X1 U11075 ( .B(ram[1402]), .A(ram[1338]), .S(n10735), .Y(n10336) );
  MUX2X1 U11076 ( .B(ram[1530]), .A(ram[1466]), .S(n10735), .Y(n10335) );
  MUX2X1 U11077 ( .B(n10334), .A(n10331), .S(n10569), .Y(n10345) );
  MUX2X1 U11078 ( .B(ram[1658]), .A(ram[1594]), .S(n10736), .Y(n10339) );
  MUX2X1 U11079 ( .B(ram[1786]), .A(ram[1722]), .S(n10736), .Y(n10338) );
  MUX2X1 U11080 ( .B(ram[1914]), .A(ram[1850]), .S(n10736), .Y(n10342) );
  MUX2X1 U11081 ( .B(ram[2042]), .A(ram[1978]), .S(n10736), .Y(n10341) );
  MUX2X1 U11082 ( .B(n10340), .A(n10337), .S(n10577), .Y(n10344) );
  MUX2X1 U11083 ( .B(n10343), .A(n10328), .S(read2_addr[0]), .Y(n10554) );
  MUX2X1 U11084 ( .B(ram[123]), .A(ram[59]), .S(n10736), .Y(n10348) );
  MUX2X1 U11085 ( .B(ram[251]), .A(ram[187]), .S(n10736), .Y(n10347) );
  MUX2X1 U11086 ( .B(ram[379]), .A(ram[315]), .S(n10736), .Y(n10351) );
  MUX2X1 U11087 ( .B(ram[507]), .A(ram[443]), .S(n10736), .Y(n10350) );
  MUX2X1 U11088 ( .B(n10349), .A(n10346), .S(n10575), .Y(n10360) );
  MUX2X1 U11089 ( .B(ram[635]), .A(ram[571]), .S(n10736), .Y(n10354) );
  MUX2X1 U11090 ( .B(ram[763]), .A(ram[699]), .S(n10736), .Y(n10353) );
  MUX2X1 U11091 ( .B(ram[891]), .A(ram[827]), .S(n10736), .Y(n10357) );
  MUX2X1 U11092 ( .B(ram[1019]), .A(ram[955]), .S(n10736), .Y(n10356) );
  MUX2X1 U11093 ( .B(n10355), .A(n10352), .S(n10576), .Y(n10359) );
  MUX2X1 U11094 ( .B(ram[1147]), .A(ram[1083]), .S(n10737), .Y(n10363) );
  MUX2X1 U11095 ( .B(ram[1275]), .A(ram[1211]), .S(n10737), .Y(n10362) );
  MUX2X1 U11096 ( .B(ram[1403]), .A(ram[1339]), .S(n10737), .Y(n10366) );
  MUX2X1 U11097 ( .B(ram[1531]), .A(ram[1467]), .S(n10737), .Y(n10365) );
  MUX2X1 U11098 ( .B(n10364), .A(n10361), .S(n10580), .Y(n10375) );
  MUX2X1 U11099 ( .B(ram[1659]), .A(ram[1595]), .S(n10737), .Y(n10369) );
  MUX2X1 U11100 ( .B(ram[1787]), .A(ram[1723]), .S(n10737), .Y(n10368) );
  MUX2X1 U11101 ( .B(ram[1915]), .A(ram[1851]), .S(n10737), .Y(n10372) );
  MUX2X1 U11102 ( .B(ram[2043]), .A(ram[1979]), .S(n10737), .Y(n10371) );
  MUX2X1 U11103 ( .B(n10370), .A(n10367), .S(n10570), .Y(n10374) );
  MUX2X1 U11104 ( .B(n10373), .A(n10358), .S(read2_addr[0]), .Y(n10555) );
  MUX2X1 U11105 ( .B(ram[124]), .A(ram[60]), .S(n10737), .Y(n10378) );
  MUX2X1 U11106 ( .B(ram[252]), .A(ram[188]), .S(n10737), .Y(n10377) );
  MUX2X1 U11107 ( .B(ram[380]), .A(ram[316]), .S(n10737), .Y(n10381) );
  MUX2X1 U11108 ( .B(ram[508]), .A(ram[444]), .S(n10737), .Y(n10380) );
  MUX2X1 U11109 ( .B(n10379), .A(n10376), .S(n10573), .Y(n10390) );
  MUX2X1 U11110 ( .B(ram[636]), .A(ram[572]), .S(n10738), .Y(n10384) );
  MUX2X1 U11111 ( .B(ram[764]), .A(ram[700]), .S(n10738), .Y(n10383) );
  MUX2X1 U11112 ( .B(ram[892]), .A(ram[828]), .S(n10738), .Y(n10387) );
  MUX2X1 U11113 ( .B(ram[1020]), .A(ram[956]), .S(n10738), .Y(n10386) );
  MUX2X1 U11114 ( .B(n10385), .A(n10382), .S(n10581), .Y(n10389) );
  MUX2X1 U11115 ( .B(ram[1148]), .A(ram[1084]), .S(n10738), .Y(n10393) );
  MUX2X1 U11116 ( .B(ram[1276]), .A(ram[1212]), .S(n10738), .Y(n10392) );
  MUX2X1 U11117 ( .B(ram[1404]), .A(ram[1340]), .S(n10738), .Y(n10396) );
  MUX2X1 U11118 ( .B(ram[1532]), .A(ram[1468]), .S(n10738), .Y(n10395) );
  MUX2X1 U11119 ( .B(n10394), .A(n10391), .S(n10579), .Y(n10405) );
  MUX2X1 U11120 ( .B(ram[1660]), .A(ram[1596]), .S(n10738), .Y(n10399) );
  MUX2X1 U11121 ( .B(ram[1788]), .A(ram[1724]), .S(n10738), .Y(n10398) );
  MUX2X1 U11122 ( .B(ram[1916]), .A(ram[1852]), .S(n10738), .Y(n10402) );
  MUX2X1 U11123 ( .B(ram[2044]), .A(ram[1980]), .S(n10738), .Y(n10401) );
  MUX2X1 U11124 ( .B(n10400), .A(n10397), .S(n10578), .Y(n10404) );
  MUX2X1 U11125 ( .B(n10403), .A(n10388), .S(n10562), .Y(n10556) );
  MUX2X1 U11126 ( .B(ram[125]), .A(ram[61]), .S(n10739), .Y(n10408) );
  MUX2X1 U11127 ( .B(ram[253]), .A(ram[189]), .S(n10739), .Y(n10407) );
  MUX2X1 U11128 ( .B(ram[381]), .A(ram[317]), .S(n10739), .Y(n10411) );
  MUX2X1 U11129 ( .B(ram[509]), .A(ram[445]), .S(n10739), .Y(n10410) );
  MUX2X1 U11130 ( .B(n10409), .A(n10406), .S(n10571), .Y(n10420) );
  MUX2X1 U11131 ( .B(ram[637]), .A(ram[573]), .S(n10739), .Y(n10414) );
  MUX2X1 U11132 ( .B(ram[765]), .A(ram[701]), .S(n10739), .Y(n10413) );
  MUX2X1 U11133 ( .B(ram[893]), .A(ram[829]), .S(n10739), .Y(n10417) );
  MUX2X1 U11134 ( .B(ram[1021]), .A(ram[957]), .S(n10739), .Y(n10416) );
  MUX2X1 U11135 ( .B(n10415), .A(n10412), .S(n10582), .Y(n10419) );
  MUX2X1 U11136 ( .B(ram[1149]), .A(ram[1085]), .S(n10739), .Y(n10423) );
  MUX2X1 U11137 ( .B(ram[1277]), .A(ram[1213]), .S(n10739), .Y(n10422) );
  MUX2X1 U11138 ( .B(ram[1405]), .A(ram[1341]), .S(n10739), .Y(n10426) );
  MUX2X1 U11139 ( .B(ram[1533]), .A(ram[1469]), .S(n10739), .Y(n10425) );
  MUX2X1 U11140 ( .B(n10424), .A(n10421), .S(n10573), .Y(n10435) );
  MUX2X1 U11141 ( .B(ram[1661]), .A(ram[1597]), .S(n10740), .Y(n10429) );
  MUX2X1 U11142 ( .B(ram[1789]), .A(ram[1725]), .S(n10740), .Y(n10428) );
  MUX2X1 U11143 ( .B(ram[1917]), .A(ram[1853]), .S(n10740), .Y(n10432) );
  MUX2X1 U11144 ( .B(ram[2045]), .A(ram[1981]), .S(n10740), .Y(n10431) );
  MUX2X1 U11145 ( .B(n10430), .A(n10427), .S(n10569), .Y(n10434) );
  MUX2X1 U11146 ( .B(n10433), .A(n10418), .S(n10562), .Y(n10557) );
  MUX2X1 U11147 ( .B(ram[126]), .A(ram[62]), .S(n10740), .Y(n10438) );
  MUX2X1 U11148 ( .B(ram[254]), .A(ram[190]), .S(n10740), .Y(n10437) );
  MUX2X1 U11149 ( .B(ram[382]), .A(ram[318]), .S(n10740), .Y(n10441) );
  MUX2X1 U11150 ( .B(ram[510]), .A(ram[446]), .S(n10740), .Y(n10440) );
  MUX2X1 U11151 ( .B(n10439), .A(n10436), .S(n10570), .Y(n10450) );
  MUX2X1 U11152 ( .B(ram[638]), .A(ram[574]), .S(n10740), .Y(n10444) );
  MUX2X1 U11153 ( .B(ram[766]), .A(ram[702]), .S(n10740), .Y(n10443) );
  MUX2X1 U11154 ( .B(ram[894]), .A(ram[830]), .S(n10740), .Y(n10447) );
  MUX2X1 U11155 ( .B(ram[1022]), .A(ram[958]), .S(n10740), .Y(n10446) );
  MUX2X1 U11156 ( .B(n10445), .A(n10442), .S(n10569), .Y(n10449) );
  MUX2X1 U11157 ( .B(ram[1150]), .A(ram[1086]), .S(n10741), .Y(n10453) );
  MUX2X1 U11158 ( .B(ram[1278]), .A(ram[1214]), .S(n10741), .Y(n10452) );
  MUX2X1 U11159 ( .B(ram[1406]), .A(ram[1342]), .S(n10741), .Y(n10456) );
  MUX2X1 U11160 ( .B(ram[1534]), .A(ram[1470]), .S(n10741), .Y(n10455) );
  MUX2X1 U11161 ( .B(n10454), .A(n10451), .S(n10579), .Y(n10465) );
  MUX2X1 U11162 ( .B(ram[1662]), .A(ram[1598]), .S(n10741), .Y(n10459) );
  MUX2X1 U11163 ( .B(ram[1790]), .A(ram[1726]), .S(n10741), .Y(n10458) );
  MUX2X1 U11164 ( .B(ram[1918]), .A(ram[1854]), .S(n10741), .Y(n10462) );
  MUX2X1 U11165 ( .B(ram[2046]), .A(ram[1982]), .S(n10741), .Y(n10461) );
  MUX2X1 U11166 ( .B(n10460), .A(n10457), .S(n10574), .Y(n10464) );
  MUX2X1 U11167 ( .B(n10463), .A(n10448), .S(n10561), .Y(n10558) );
  MUX2X1 U11168 ( .B(ram[127]), .A(ram[63]), .S(n10741), .Y(n10468) );
  MUX2X1 U11169 ( .B(ram[255]), .A(ram[191]), .S(n10741), .Y(n10467) );
  MUX2X1 U11170 ( .B(ram[383]), .A(ram[319]), .S(n10741), .Y(n10471) );
  MUX2X1 U11171 ( .B(ram[511]), .A(ram[447]), .S(n10741), .Y(n10470) );
  MUX2X1 U11172 ( .B(n10469), .A(n10466), .S(n10576), .Y(n10480) );
  MUX2X1 U11173 ( .B(ram[639]), .A(ram[575]), .S(n10742), .Y(n10474) );
  MUX2X1 U11174 ( .B(ram[767]), .A(ram[703]), .S(n10742), .Y(n10473) );
  MUX2X1 U11175 ( .B(ram[895]), .A(ram[831]), .S(n10742), .Y(n10477) );
  MUX2X1 U11176 ( .B(ram[1023]), .A(ram[959]), .S(n10742), .Y(n10476) );
  MUX2X1 U11177 ( .B(n10475), .A(n10472), .S(n10575), .Y(n10479) );
  MUX2X1 U11178 ( .B(ram[1151]), .A(ram[1087]), .S(n10742), .Y(n10483) );
  MUX2X1 U11179 ( .B(ram[1279]), .A(ram[1215]), .S(n10742), .Y(n10482) );
  MUX2X1 U11180 ( .B(ram[1407]), .A(ram[1343]), .S(n10742), .Y(n10486) );
  MUX2X1 U11181 ( .B(ram[1535]), .A(ram[1471]), .S(n10742), .Y(n10485) );
  MUX2X1 U11182 ( .B(n10484), .A(n10481), .S(n10580), .Y(n10495) );
  MUX2X1 U11183 ( .B(ram[1663]), .A(ram[1599]), .S(n10742), .Y(n10489) );
  MUX2X1 U11184 ( .B(ram[1791]), .A(ram[1727]), .S(n10742), .Y(n10488) );
  MUX2X1 U11185 ( .B(ram[1919]), .A(ram[1855]), .S(n10742), .Y(n10492) );
  MUX2X1 U11186 ( .B(ram[2047]), .A(ram[1983]), .S(n10742), .Y(n10491) );
  MUX2X1 U11187 ( .B(n10490), .A(n10487), .S(n10572), .Y(n10494) );
  MUX2X1 U11188 ( .B(n10493), .A(n10478), .S(read2_addr[0]), .Y(n10559) );
  NAND3X1 U11189 ( .A(PPP[1]), .B(n13228), .C(n11016), .Y(n11017) );
  NAND3X1 U11190 ( .A(PPP[2]), .B(PPP[1]), .C(n11016), .Y(n10977) );
  OAI21X1 U11191 ( .A(n4668), .B(n11016), .C(n1677), .Y(n10966) );
  NAND3X1 U11192 ( .A(PPP[2]), .B(n13227), .C(n11016), .Y(n11014) );
  AOI22X1 U11193 ( .A(Din[63]), .B(n10749), .C(current_ram[63]), .D(n10751), 
        .Y(n13099) );
  NAND3X1 U11194 ( .A(n4508), .B(n4577), .C(n4578), .Y(n10968) );
  NAND3X1 U11195 ( .A(n4576), .B(n4579), .C(n4580), .Y(n10967) );
  MUX2X1 U11196 ( .B(n186), .A(n10827), .S(n10761), .Y(n10969) );
  AOI22X1 U11197 ( .A(Din[62]), .B(n10749), .C(current_ram[62]), .D(n10751), 
        .Y(n13101) );
  MUX2X1 U11198 ( .B(n185), .A(n10829), .S(n10761), .Y(n10970) );
  AOI22X1 U11199 ( .A(Din[61]), .B(n10749), .C(current_ram[61]), .D(n10751), 
        .Y(n13103) );
  MUX2X1 U11200 ( .B(n184), .A(n10831), .S(n10761), .Y(n10971) );
  AOI22X1 U11201 ( .A(Din[60]), .B(n10749), .C(current_ram[60]), .D(n10751), 
        .Y(n13105) );
  MUX2X1 U11202 ( .B(n183), .A(n10833), .S(n10761), .Y(n10972) );
  AOI22X1 U11203 ( .A(Din[59]), .B(n10749), .C(current_ram[59]), .D(n10751), 
        .Y(n13107) );
  MUX2X1 U11204 ( .B(n182), .A(n10835), .S(n10761), .Y(n10973) );
  AOI22X1 U11205 ( .A(Din[58]), .B(n10749), .C(current_ram[58]), .D(n10751), 
        .Y(n13109) );
  MUX2X1 U11206 ( .B(n181), .A(n10837), .S(n10761), .Y(n10974) );
  AOI22X1 U11207 ( .A(Din[57]), .B(n10749), .C(current_ram[57]), .D(n10751), 
        .Y(n13111) );
  MUX2X1 U11208 ( .B(n180), .A(n10839), .S(n10761), .Y(n10975) );
  AOI22X1 U11209 ( .A(Din[56]), .B(n10749), .C(current_ram[56]), .D(n10751), 
        .Y(n13113) );
  MUX2X1 U11210 ( .B(n179), .A(n10841), .S(n10761), .Y(n10976) );
  OAI21X1 U11211 ( .A(n1993), .B(PPP[0]), .C(n1677), .Y(n10978) );
  AOI22X1 U11212 ( .A(Din[55]), .B(n10752), .C(current_ram[55]), .D(n10754), 
        .Y(n13115) );
  MUX2X1 U11213 ( .B(n178), .A(n10843), .S(n10761), .Y(n10979) );
  AOI22X1 U11214 ( .A(Din[54]), .B(n10752), .C(current_ram[54]), .D(n10754), 
        .Y(n13117) );
  MUX2X1 U11215 ( .B(n177), .A(n10845), .S(n10761), .Y(n10980) );
  AOI22X1 U11216 ( .A(Din[53]), .B(n10752), .C(current_ram[53]), .D(n10754), 
        .Y(n13119) );
  MUX2X1 U11217 ( .B(n176), .A(n10847), .S(n10761), .Y(n10981) );
  AOI22X1 U11218 ( .A(Din[52]), .B(n10752), .C(current_ram[52]), .D(n10754), 
        .Y(n13121) );
  MUX2X1 U11219 ( .B(n175), .A(n10849), .S(n10761), .Y(n10982) );
  AOI22X1 U11220 ( .A(Din[51]), .B(n10752), .C(current_ram[51]), .D(n10754), 
        .Y(n13123) );
  MUX2X1 U11221 ( .B(n174), .A(n10851), .S(n10762), .Y(n10983) );
  AOI22X1 U11222 ( .A(Din[50]), .B(n10752), .C(current_ram[50]), .D(n10754), 
        .Y(n13125) );
  MUX2X1 U11223 ( .B(n173), .A(n10853), .S(n10762), .Y(n10984) );
  AOI22X1 U11224 ( .A(Din[49]), .B(n10752), .C(current_ram[49]), .D(n10754), 
        .Y(n13127) );
  MUX2X1 U11225 ( .B(n172), .A(n10855), .S(n10762), .Y(n10985) );
  AOI22X1 U11226 ( .A(Din[48]), .B(n10752), .C(current_ram[48]), .D(n10754), 
        .Y(n13129) );
  MUX2X1 U11227 ( .B(n171), .A(n10857), .S(n10762), .Y(n10986) );
  AOI22X1 U11228 ( .A(Din[47]), .B(n10750), .C(current_ram[47]), .D(n10751), 
        .Y(n13131) );
  MUX2X1 U11229 ( .B(n170), .A(n10859), .S(n10762), .Y(n10987) );
  AOI22X1 U11230 ( .A(Din[46]), .B(n10750), .C(current_ram[46]), .D(n10751), 
        .Y(n13133) );
  MUX2X1 U11231 ( .B(n169), .A(n10861), .S(n10762), .Y(n10988) );
  AOI22X1 U11232 ( .A(Din[45]), .B(n10750), .C(current_ram[45]), .D(n10751), 
        .Y(n13135) );
  MUX2X1 U11233 ( .B(n168), .A(n10863), .S(n10762), .Y(n10989) );
  AOI22X1 U11234 ( .A(Din[44]), .B(n10750), .C(current_ram[44]), .D(n10751), 
        .Y(n13137) );
  MUX2X1 U11235 ( .B(n167), .A(n10865), .S(n10762), .Y(n10990) );
  AOI22X1 U11236 ( .A(Din[43]), .B(n10750), .C(current_ram[43]), .D(n10751), 
        .Y(n13139) );
  MUX2X1 U11237 ( .B(n166), .A(n10867), .S(n10762), .Y(n10991) );
  AOI22X1 U11238 ( .A(Din[42]), .B(n10750), .C(current_ram[42]), .D(n10751), 
        .Y(n13141) );
  MUX2X1 U11239 ( .B(n165), .A(n10869), .S(n10762), .Y(n10992) );
  AOI22X1 U11240 ( .A(Din[41]), .B(n10750), .C(current_ram[41]), .D(n10751), 
        .Y(n13143) );
  MUX2X1 U11241 ( .B(n164), .A(n10871), .S(n10762), .Y(n10993) );
  AOI22X1 U11242 ( .A(Din[40]), .B(n10750), .C(current_ram[40]), .D(n10751), 
        .Y(n13145) );
  MUX2X1 U11243 ( .B(n163), .A(n10873), .S(n10762), .Y(n10995) );
  AOI22X1 U11244 ( .A(Din[39]), .B(n10753), .C(current_ram[39]), .D(n10754), 
        .Y(n13147) );
  MUX2X1 U11245 ( .B(n162), .A(n10875), .S(n10761), .Y(n10996) );
  AOI22X1 U11246 ( .A(Din[38]), .B(n10753), .C(current_ram[38]), .D(n10754), 
        .Y(n13149) );
  MUX2X1 U11247 ( .B(n161), .A(n10877), .S(n10762), .Y(n10997) );
  AOI22X1 U11248 ( .A(Din[37]), .B(n10753), .C(current_ram[37]), .D(n10754), 
        .Y(n13151) );
  MUX2X1 U11249 ( .B(n160), .A(n10879), .S(n10761), .Y(n10998) );
  AOI22X1 U11250 ( .A(Din[36]), .B(n10753), .C(current_ram[36]), .D(n10754), 
        .Y(n13153) );
  MUX2X1 U11251 ( .B(n159), .A(n10881), .S(n10762), .Y(n10999) );
  AOI22X1 U11252 ( .A(Din[35]), .B(n10753), .C(current_ram[35]), .D(n10754), 
        .Y(n13155) );
  MUX2X1 U11253 ( .B(n158), .A(n10883), .S(n10761), .Y(n11000) );
  AOI22X1 U11254 ( .A(Din[34]), .B(n10753), .C(current_ram[34]), .D(n10754), 
        .Y(n13157) );
  MUX2X1 U11255 ( .B(n157), .A(n10885), .S(n10762), .Y(n11001) );
  AOI22X1 U11256 ( .A(Din[33]), .B(n10753), .C(current_ram[33]), .D(n10754), 
        .Y(n13159) );
  MUX2X1 U11257 ( .B(n156), .A(n10887), .S(n10761), .Y(n11002) );
  AOI22X1 U11258 ( .A(Din[32]), .B(n10753), .C(current_ram[32]), .D(n10754), 
        .Y(n13161) );
  MUX2X1 U11259 ( .B(n155), .A(n10889), .S(n10762), .Y(n11004) );
  AOI22X1 U11260 ( .A(Din[31]), .B(n10755), .C(current_ram[31]), .D(n10757), 
        .Y(n13163) );
  MUX2X1 U11261 ( .B(n154), .A(n10891), .S(n10761), .Y(n11006) );
  AOI22X1 U11262 ( .A(Din[30]), .B(n10755), .C(current_ram[30]), .D(n10757), 
        .Y(n13165) );
  MUX2X1 U11263 ( .B(n153), .A(n10893), .S(n10762), .Y(n11007) );
  AOI22X1 U11264 ( .A(Din[29]), .B(n10755), .C(current_ram[29]), .D(n10757), 
        .Y(n13167) );
  MUX2X1 U11265 ( .B(n152), .A(n10895), .S(n10761), .Y(n11008) );
  AOI22X1 U11266 ( .A(Din[28]), .B(n10755), .C(current_ram[28]), .D(n10757), 
        .Y(n13169) );
  MUX2X1 U11267 ( .B(n151), .A(n10897), .S(n10761), .Y(n11009) );
  AOI22X1 U11268 ( .A(Din[27]), .B(n10755), .C(current_ram[27]), .D(n10757), 
        .Y(n13171) );
  MUX2X1 U11269 ( .B(n150), .A(n10899), .S(n10762), .Y(n11010) );
  AOI22X1 U11270 ( .A(Din[26]), .B(n10755), .C(current_ram[26]), .D(n10757), 
        .Y(n13173) );
  MUX2X1 U11271 ( .B(n149), .A(n10901), .S(n10762), .Y(n11011) );
  AOI22X1 U11272 ( .A(Din[25]), .B(n10755), .C(current_ram[25]), .D(n10757), 
        .Y(n13175) );
  MUX2X1 U11273 ( .B(n148), .A(n10903), .S(n10761), .Y(n11012) );
  AOI22X1 U11274 ( .A(Din[24]), .B(n10755), .C(current_ram[24]), .D(n10757), 
        .Y(n13177) );
  MUX2X1 U11275 ( .B(n147), .A(n10905), .S(n10761), .Y(n11013) );
  AOI22X1 U11276 ( .A(n1), .B(n10758), .C(current_ram[23]), .D(n10760), .Y(
        n13179) );
  MUX2X1 U11277 ( .B(n146), .A(n10907), .S(n10761), .Y(n11018) );
  AOI22X1 U11278 ( .A(Din[22]), .B(n10758), .C(current_ram[22]), .D(n10760), 
        .Y(n13181) );
  MUX2X1 U11279 ( .B(n145), .A(n10909), .S(n10762), .Y(n11019) );
  AOI22X1 U11280 ( .A(Din[21]), .B(n10758), .C(current_ram[21]), .D(n10760), 
        .Y(n13183) );
  MUX2X1 U11281 ( .B(n144), .A(n10911), .S(n10762), .Y(n11020) );
  AOI22X1 U11282 ( .A(Din[20]), .B(n10758), .C(current_ram[20]), .D(n10760), 
        .Y(n13185) );
  MUX2X1 U11283 ( .B(n143), .A(n10913), .S(n10762), .Y(n11021) );
  AOI22X1 U11284 ( .A(Din[19]), .B(n10758), .C(current_ram[19]), .D(n10760), 
        .Y(n13187) );
  MUX2X1 U11285 ( .B(n142), .A(n10915), .S(n10761), .Y(n11022) );
  AOI22X1 U11286 ( .A(Din[18]), .B(n10758), .C(current_ram[18]), .D(n10760), 
        .Y(n13189) );
  MUX2X1 U11287 ( .B(n141), .A(n10917), .S(n10762), .Y(n11023) );
  AOI22X1 U11288 ( .A(Din[17]), .B(n10758), .C(current_ram[17]), .D(n10760), 
        .Y(n13191) );
  MUX2X1 U11289 ( .B(n140), .A(n10919), .S(n10761), .Y(n11024) );
  AOI22X1 U11290 ( .A(Din[16]), .B(n10758), .C(current_ram[16]), .D(n10760), 
        .Y(n13193) );
  MUX2X1 U11291 ( .B(n139), .A(n10921), .S(n10761), .Y(n11025) );
  AOI22X1 U11292 ( .A(Din[15]), .B(n10756), .C(current_ram[15]), .D(n10757), 
        .Y(n13195) );
  MUX2X1 U11293 ( .B(n138), .A(n10923), .S(n10762), .Y(n11026) );
  AOI22X1 U11294 ( .A(Din[14]), .B(n10756), .C(current_ram[14]), .D(n10757), 
        .Y(n13197) );
  MUX2X1 U11295 ( .B(n137), .A(n10925), .S(n10761), .Y(n11027) );
  AOI22X1 U11296 ( .A(Din[13]), .B(n10756), .C(current_ram[13]), .D(n10757), 
        .Y(n13199) );
  MUX2X1 U11297 ( .B(n136), .A(n10927), .S(n10762), .Y(n11028) );
  AOI22X1 U11298 ( .A(Din[12]), .B(n10756), .C(current_ram[12]), .D(n10757), 
        .Y(n13201) );
  MUX2X1 U11299 ( .B(n135), .A(n10929), .S(n10762), .Y(n11029) );
  AOI22X1 U11300 ( .A(Din[11]), .B(n10756), .C(current_ram[11]), .D(n10757), 
        .Y(n13203) );
  MUX2X1 U11301 ( .B(n134), .A(n10931), .S(n10762), .Y(n11030) );
  AOI22X1 U11302 ( .A(Din[10]), .B(n10756), .C(current_ram[10]), .D(n10757), 
        .Y(n13205) );
  MUX2X1 U11303 ( .B(n133), .A(n10933), .S(n10761), .Y(n11031) );
  AOI22X1 U11304 ( .A(Din[9]), .B(n10756), .C(current_ram[9]), .D(n10757), .Y(
        n13207) );
  MUX2X1 U11305 ( .B(n132), .A(n10935), .S(n10762), .Y(n11032) );
  AOI22X1 U11306 ( .A(Din[8]), .B(n10756), .C(current_ram[8]), .D(n10757), .Y(
        n13209) );
  MUX2X1 U11307 ( .B(n131), .A(n10937), .S(n10761), .Y(n11034) );
  AOI22X1 U11308 ( .A(Din[7]), .B(n10759), .C(current_ram[7]), .D(n10760), .Y(
        n13211) );
  MUX2X1 U11309 ( .B(n130), .A(n10939), .S(n10761), .Y(n11035) );
  AOI22X1 U11310 ( .A(Din[6]), .B(n10759), .C(current_ram[6]), .D(n10760), .Y(
        n13213) );
  MUX2X1 U11311 ( .B(n129), .A(n10941), .S(n10761), .Y(n11036) );
  AOI22X1 U11312 ( .A(Din[5]), .B(n10759), .C(current_ram[5]), .D(n10760), .Y(
        n13215) );
  MUX2X1 U11313 ( .B(n128), .A(n10943), .S(n10762), .Y(n11037) );
  AOI22X1 U11314 ( .A(Din[4]), .B(n10759), .C(current_ram[4]), .D(n10760), .Y(
        n13217) );
  MUX2X1 U11315 ( .B(n127), .A(n10945), .S(n10762), .Y(n11038) );
  AOI22X1 U11316 ( .A(Din[3]), .B(n10759), .C(current_ram[3]), .D(n10760), .Y(
        n13219) );
  MUX2X1 U11317 ( .B(n126), .A(n10947), .S(n10762), .Y(n11039) );
  AOI22X1 U11318 ( .A(Din[2]), .B(n10759), .C(current_ram[2]), .D(n10760), .Y(
        n13221) );
  MUX2X1 U11319 ( .B(n125), .A(n10949), .S(n10762), .Y(n11040) );
  AOI22X1 U11320 ( .A(Din[1]), .B(n10759), .C(current_ram[1]), .D(n10760), .Y(
        n13223) );
  MUX2X1 U11321 ( .B(n124), .A(n10951), .S(n10761), .Y(n11041) );
  AOI22X1 U11322 ( .A(Din[0]), .B(n10759), .C(current_ram[0]), .D(n10760), .Y(
        n13226) );
  MUX2X1 U11323 ( .B(n123), .A(n10955), .S(n10761), .Y(n11044) );
  NAND3X1 U11324 ( .A(n4508), .B(n4663), .C(n4664), .Y(n11046) );
  NAND3X1 U11325 ( .A(n4662), .B(n4665), .C(n4666), .Y(n11045) );
  MUX2X1 U11326 ( .B(n119), .A(n10827), .S(n10763), .Y(n11047) );
  MUX2X1 U11327 ( .B(n118), .A(n10829), .S(n10764), .Y(n11048) );
  MUX2X1 U11328 ( .B(n117), .A(n10831), .S(n10763), .Y(n11049) );
  MUX2X1 U11329 ( .B(n116), .A(n10833), .S(n10765), .Y(n11050) );
  MUX2X1 U11330 ( .B(n115), .A(n10835), .S(n10765), .Y(n11051) );
  MUX2X1 U11331 ( .B(n114), .A(n10837), .S(n10765), .Y(n11052) );
  MUX2X1 U11332 ( .B(n113), .A(n10839), .S(n10764), .Y(n11053) );
  MUX2X1 U11333 ( .B(n112), .A(n10841), .S(n10764), .Y(n11054) );
  MUX2X1 U11334 ( .B(n111), .A(n10843), .S(n10765), .Y(n11055) );
  MUX2X1 U11335 ( .B(n110), .A(n10845), .S(n10763), .Y(n11056) );
  MUX2X1 U11336 ( .B(n109), .A(n10847), .S(n10764), .Y(n11057) );
  MUX2X1 U11337 ( .B(n108), .A(n10849), .S(n10763), .Y(n11058) );
  MUX2X1 U11338 ( .B(n107), .A(n10851), .S(n10763), .Y(n11059) );
  MUX2X1 U11339 ( .B(n106), .A(n10853), .S(n10763), .Y(n11060) );
  MUX2X1 U11340 ( .B(n105), .A(n10855), .S(n10763), .Y(n11061) );
  MUX2X1 U11341 ( .B(n104), .A(n10857), .S(n10763), .Y(n11062) );
  MUX2X1 U11342 ( .B(n103), .A(n10859), .S(n10763), .Y(n11063) );
  MUX2X1 U11343 ( .B(n102), .A(n10861), .S(n10763), .Y(n11064) );
  MUX2X1 U11344 ( .B(n101), .A(n10863), .S(n10763), .Y(n11065) );
  MUX2X1 U11345 ( .B(n100), .A(n10865), .S(n10763), .Y(n11066) );
  MUX2X1 U11346 ( .B(n99), .A(n10867), .S(n10763), .Y(n11067) );
  MUX2X1 U11347 ( .B(n98), .A(n10869), .S(n10763), .Y(n11068) );
  MUX2X1 U11348 ( .B(n97), .A(n10871), .S(n10763), .Y(n11069) );
  MUX2X1 U11349 ( .B(n96), .A(n10873), .S(n10763), .Y(n11070) );
  MUX2X1 U11350 ( .B(n95), .A(n10875), .S(n10765), .Y(n11071) );
  MUX2X1 U11351 ( .B(n94), .A(n10877), .S(n10763), .Y(n11072) );
  MUX2X1 U11352 ( .B(n93), .A(n10879), .S(n10764), .Y(n11073) );
  MUX2X1 U11353 ( .B(n92), .A(n10881), .S(n10763), .Y(n11074) );
  MUX2X1 U11354 ( .B(n91), .A(n10883), .S(n10765), .Y(n11075) );
  MUX2X1 U11355 ( .B(n90), .A(n10885), .S(n10765), .Y(n11076) );
  MUX2X1 U11356 ( .B(n89), .A(n10887), .S(n10763), .Y(n11077) );
  MUX2X1 U11357 ( .B(n88), .A(n10889), .S(n10763), .Y(n11078) );
  MUX2X1 U11358 ( .B(n87), .A(n10891), .S(n10764), .Y(n11079) );
  MUX2X1 U11359 ( .B(n86), .A(n10893), .S(n10763), .Y(n11080) );
  MUX2X1 U11360 ( .B(n85), .A(n10895), .S(n10765), .Y(n11081) );
  MUX2X1 U11361 ( .B(n84), .A(n10897), .S(n10764), .Y(n11082) );
  MUX2X1 U11362 ( .B(n83), .A(n10899), .S(n10764), .Y(n11083) );
  MUX2X1 U11363 ( .B(n82), .A(n10901), .S(n10764), .Y(n11084) );
  MUX2X1 U11364 ( .B(n81), .A(n10903), .S(n10764), .Y(n11085) );
  MUX2X1 U11365 ( .B(n80), .A(n10905), .S(n10764), .Y(n11086) );
  MUX2X1 U11366 ( .B(n79), .A(n10907), .S(n10764), .Y(n11087) );
  MUX2X1 U11367 ( .B(n78), .A(n10909), .S(n10764), .Y(n11088) );
  MUX2X1 U11368 ( .B(n77), .A(n10911), .S(n10764), .Y(n11089) );
  MUX2X1 U11369 ( .B(n76), .A(n10913), .S(n10764), .Y(n11090) );
  MUX2X1 U11370 ( .B(n75), .A(n10915), .S(n10764), .Y(n11091) );
  MUX2X1 U11371 ( .B(n74), .A(n10917), .S(n10764), .Y(n11092) );
  MUX2X1 U11372 ( .B(n73), .A(n10919), .S(n10764), .Y(n11093) );
  MUX2X1 U11373 ( .B(n72), .A(n10921), .S(n10764), .Y(n11094) );
  MUX2X1 U11374 ( .B(n71), .A(n10923), .S(n10765), .Y(n11095) );
  MUX2X1 U11375 ( .B(n70), .A(n10925), .S(n10765), .Y(n11096) );
  MUX2X1 U11376 ( .B(n69), .A(n10927), .S(n10765), .Y(n11097) );
  MUX2X1 U11377 ( .B(n68), .A(n10929), .S(n10765), .Y(n11098) );
  MUX2X1 U11378 ( .B(n67), .A(n10931), .S(n10765), .Y(n11099) );
  MUX2X1 U11379 ( .B(n66), .A(n10933), .S(n10765), .Y(n11100) );
  MUX2X1 U11380 ( .B(n65), .A(n10935), .S(n10765), .Y(n11101) );
  MUX2X1 U11381 ( .B(n64), .A(n10937), .S(n10765), .Y(n11102) );
  MUX2X1 U11382 ( .B(n63), .A(n10939), .S(n10765), .Y(n11103) );
  MUX2X1 U11383 ( .B(n62), .A(n10941), .S(n10765), .Y(n11104) );
  MUX2X1 U11384 ( .B(n61), .A(n10943), .S(n10765), .Y(n11105) );
  MUX2X1 U11385 ( .B(n60), .A(n10945), .S(n10765), .Y(n11106) );
  MUX2X1 U11386 ( .B(n59), .A(n10947), .S(n10764), .Y(n11107) );
  MUX2X1 U11387 ( .B(n58), .A(n10949), .S(n10764), .Y(n11108) );
  MUX2X1 U11388 ( .B(n57), .A(n10951), .S(n10765), .Y(n11109) );
  MUX2X1 U11389 ( .B(n56), .A(n10955), .S(n10764), .Y(n11111) );
  NAND3X1 U11390 ( .A(n4152), .B(n10963), .C(n11112), .Y(n11575) );
  OAI21X1 U11391 ( .A(n1520), .B(n2153), .C(n10956), .Y(n11113) );
  OAI21X1 U11392 ( .A(n10826), .B(n10767), .C(n2149), .Y(n4669) );
  OAI21X1 U11393 ( .A(n10828), .B(n10767), .C(n1992), .Y(n4670) );
  OAI21X1 U11394 ( .A(n10830), .B(n10767), .C(n1834), .Y(n4671) );
  OAI21X1 U11395 ( .A(n10832), .B(n10767), .C(n1675), .Y(n4672) );
  OAI21X1 U11396 ( .A(n10834), .B(n10767), .C(n1518), .Y(n4673) );
  OAI21X1 U11397 ( .A(n10836), .B(n10767), .C(n1392), .Y(n4674) );
  OAI21X1 U11398 ( .A(n10838), .B(n10767), .C(n1267), .Y(n4675) );
  OAI21X1 U11399 ( .A(n10840), .B(n10767), .C(n1142), .Y(n4676) );
  OAI21X1 U11400 ( .A(n10842), .B(n10767), .C(n1019), .Y(n4677) );
  OAI21X1 U11401 ( .A(n10844), .B(n10767), .C(n907), .Y(n4678) );
  OAI21X1 U11402 ( .A(n10846), .B(n10767), .C(n795), .Y(n4679) );
  OAI21X1 U11403 ( .A(n10848), .B(n10767), .C(n683), .Y(n4680) );
  OAI21X1 U11404 ( .A(n10850), .B(n10767), .C(n2148), .Y(n4681) );
  OAI21X1 U11405 ( .A(n10852), .B(n10767), .C(n1991), .Y(n4682) );
  OAI21X1 U11406 ( .A(n10854), .B(n10767), .C(n1833), .Y(n4683) );
  OAI21X1 U11407 ( .A(n10856), .B(n10767), .C(n1674), .Y(n4684) );
  OAI21X1 U11408 ( .A(n10858), .B(n10767), .C(n1517), .Y(n4685) );
  OAI21X1 U11409 ( .A(n10860), .B(n10767), .C(n1391), .Y(n4686) );
  OAI21X1 U11410 ( .A(n10862), .B(n10767), .C(n1266), .Y(n4687) );
  OAI21X1 U11411 ( .A(n10864), .B(n10767), .C(n1141), .Y(n4688) );
  OAI21X1 U11412 ( .A(n10866), .B(n10767), .C(n1018), .Y(n4689) );
  OAI21X1 U11413 ( .A(n10868), .B(n10767), .C(n906), .Y(n4690) );
  OAI21X1 U11414 ( .A(n10870), .B(n10767), .C(n794), .Y(n4691) );
  OAI21X1 U11415 ( .A(n10872), .B(n10767), .C(n682), .Y(n4692) );
  OAI21X1 U11416 ( .A(n10874), .B(n10767), .C(n575), .Y(n4693) );
  OAI21X1 U11417 ( .A(n10876), .B(n10767), .C(n2147), .Y(n4694) );
  OAI21X1 U11418 ( .A(n10878), .B(n10767), .C(n1990), .Y(n4695) );
  OAI21X1 U11419 ( .A(n10880), .B(n10767), .C(n1832), .Y(n4696) );
  OAI21X1 U11420 ( .A(n10882), .B(n10767), .C(n1673), .Y(n4697) );
  OAI21X1 U11421 ( .A(n10884), .B(n10767), .C(n1516), .Y(n4698) );
  OAI21X1 U11422 ( .A(n10886), .B(n10767), .C(n1390), .Y(n4699) );
  OAI21X1 U11423 ( .A(n10888), .B(n10767), .C(n1265), .Y(n4700) );
  OAI21X1 U11424 ( .A(n10890), .B(n10767), .C(n1140), .Y(n4701) );
  OAI21X1 U11425 ( .A(n10892), .B(n10767), .C(n1017), .Y(n4702) );
  OAI21X1 U11426 ( .A(n10894), .B(n10767), .C(n905), .Y(n4703) );
  OAI21X1 U11427 ( .A(n10896), .B(n10767), .C(n793), .Y(n4704) );
  OAI21X1 U11428 ( .A(n10898), .B(n10767), .C(n681), .Y(n4705) );
  OAI21X1 U11429 ( .A(n10900), .B(n10767), .C(n574), .Y(n4706) );
  OAI21X1 U11430 ( .A(n10902), .B(n10767), .C(n2146), .Y(n4707) );
  OAI21X1 U11431 ( .A(n10904), .B(n10767), .C(n1989), .Y(n4708) );
  OAI21X1 U11432 ( .A(n10906), .B(n10767), .C(n1831), .Y(n4709) );
  OAI21X1 U11433 ( .A(n10908), .B(n10767), .C(n1672), .Y(n4710) );
  OAI21X1 U11434 ( .A(n10910), .B(n10767), .C(n1515), .Y(n4711) );
  OAI21X1 U11435 ( .A(n10912), .B(n10767), .C(n1389), .Y(n4712) );
  OAI21X1 U11436 ( .A(n10914), .B(n10767), .C(n1264), .Y(n4713) );
  OAI21X1 U11437 ( .A(n10916), .B(n10767), .C(n1139), .Y(n4714) );
  OAI21X1 U11438 ( .A(n10918), .B(n10767), .C(n1016), .Y(n4715) );
  OAI21X1 U11439 ( .A(n10920), .B(n10767), .C(n904), .Y(n4716) );
  OAI21X1 U11440 ( .A(n10922), .B(n10767), .C(n792), .Y(n4717) );
  OAI21X1 U11441 ( .A(n10924), .B(n10767), .C(n680), .Y(n4718) );
  OAI21X1 U11442 ( .A(n10926), .B(n10767), .C(n573), .Y(n4719) );
  OAI21X1 U11443 ( .A(n10928), .B(n10767), .C(n2145), .Y(n4720) );
  OAI21X1 U11444 ( .A(n10930), .B(n10767), .C(n1988), .Y(n4721) );
  OAI21X1 U11445 ( .A(n10932), .B(n10767), .C(n1830), .Y(n4722) );
  OAI21X1 U11446 ( .A(n10934), .B(n10767), .C(n1671), .Y(n4723) );
  OAI21X1 U11447 ( .A(n10936), .B(n10767), .C(n1514), .Y(n4724) );
  OAI21X1 U11448 ( .A(n10938), .B(n10767), .C(n1388), .Y(n4725) );
  OAI21X1 U11449 ( .A(n10940), .B(n10767), .C(n1263), .Y(n4726) );
  OAI21X1 U11450 ( .A(n10942), .B(n10767), .C(n1138), .Y(n4727) );
  OAI21X1 U11451 ( .A(n10944), .B(n10767), .C(n1015), .Y(n4728) );
  OAI21X1 U11452 ( .A(n10946), .B(n10767), .C(n903), .Y(n4729) );
  OAI21X1 U11453 ( .A(n10948), .B(n10767), .C(n791), .Y(n4730) );
  OAI21X1 U11454 ( .A(n10950), .B(n10767), .C(n679), .Y(n4731) );
  OAI21X1 U11455 ( .A(n10954), .B(n10767), .C(n572), .Y(n4732) );
  OAI21X1 U11456 ( .A(n1395), .B(n2153), .C(n10956), .Y(n11179) );
  OAI21X1 U11457 ( .A(n10826), .B(n10769), .C(n1987), .Y(n4733) );
  OAI21X1 U11458 ( .A(n10828), .B(n10769), .C(n2144), .Y(n4734) );
  OAI21X1 U11459 ( .A(n10830), .B(n10769), .C(n1670), .Y(n4735) );
  OAI21X1 U11460 ( .A(n10832), .B(n10769), .C(n1829), .Y(n4736) );
  OAI21X1 U11461 ( .A(n10834), .B(n10769), .C(n1387), .Y(n4737) );
  OAI21X1 U11462 ( .A(n10836), .B(n10769), .C(n1513), .Y(n4738) );
  OAI21X1 U11463 ( .A(n10838), .B(n10769), .C(n1137), .Y(n4739) );
  OAI21X1 U11464 ( .A(n10840), .B(n10769), .C(n1262), .Y(n4740) );
  OAI21X1 U11465 ( .A(n10842), .B(n10769), .C(n902), .Y(n4741) );
  OAI21X1 U11466 ( .A(n10844), .B(n10769), .C(n1014), .Y(n4742) );
  OAI21X1 U11467 ( .A(n10846), .B(n10769), .C(n678), .Y(n4743) );
  OAI21X1 U11468 ( .A(n10848), .B(n10769), .C(n790), .Y(n4744) );
  OAI21X1 U11469 ( .A(n10850), .B(n10769), .C(n1986), .Y(n4745) );
  OAI21X1 U11470 ( .A(n10852), .B(n10769), .C(n2143), .Y(n4746) );
  OAI21X1 U11471 ( .A(n10854), .B(n10769), .C(n1669), .Y(n4747) );
  OAI21X1 U11472 ( .A(n10856), .B(n10769), .C(n1828), .Y(n4748) );
  OAI21X1 U11473 ( .A(n10858), .B(n10769), .C(n1386), .Y(n4749) );
  OAI21X1 U11474 ( .A(n10860), .B(n10769), .C(n1512), .Y(n4750) );
  OAI21X1 U11475 ( .A(n10862), .B(n10769), .C(n1136), .Y(n4751) );
  OAI21X1 U11476 ( .A(n10864), .B(n10769), .C(n1261), .Y(n4752) );
  OAI21X1 U11477 ( .A(n10866), .B(n10769), .C(n901), .Y(n4753) );
  OAI21X1 U11478 ( .A(n10868), .B(n10769), .C(n1013), .Y(n4754) );
  OAI21X1 U11479 ( .A(n10870), .B(n10769), .C(n677), .Y(n4755) );
  OAI21X1 U11480 ( .A(n10872), .B(n10769), .C(n789), .Y(n4756) );
  OAI21X1 U11481 ( .A(n10874), .B(n10769), .C(n468), .Y(n4757) );
  OAI21X1 U11482 ( .A(n10876), .B(n10769), .C(n1985), .Y(n4758) );
  OAI21X1 U11483 ( .A(n10878), .B(n10769), .C(n2142), .Y(n4759) );
  OAI21X1 U11484 ( .A(n10880), .B(n10769), .C(n1668), .Y(n4760) );
  OAI21X1 U11485 ( .A(n10882), .B(n10769), .C(n1827), .Y(n4761) );
  OAI21X1 U11486 ( .A(n10884), .B(n10769), .C(n1385), .Y(n4762) );
  OAI21X1 U11487 ( .A(n10886), .B(n10769), .C(n1511), .Y(n4763) );
  OAI21X1 U11488 ( .A(n10888), .B(n10769), .C(n1135), .Y(n4764) );
  OAI21X1 U11489 ( .A(n10890), .B(n10769), .C(n1260), .Y(n4765) );
  OAI21X1 U11490 ( .A(n10892), .B(n10769), .C(n900), .Y(n4766) );
  OAI21X1 U11491 ( .A(n10894), .B(n10769), .C(n1012), .Y(n4767) );
  OAI21X1 U11492 ( .A(n10896), .B(n10769), .C(n676), .Y(n4768) );
  OAI21X1 U11493 ( .A(n10898), .B(n10769), .C(n788), .Y(n4769) );
  OAI21X1 U11494 ( .A(n10900), .B(n10769), .C(n467), .Y(n4770) );
  OAI21X1 U11495 ( .A(n10902), .B(n10769), .C(n1984), .Y(n4771) );
  OAI21X1 U11496 ( .A(n10904), .B(n10769), .C(n2141), .Y(n4772) );
  OAI21X1 U11497 ( .A(n10906), .B(n10769), .C(n1667), .Y(n4773) );
  OAI21X1 U11498 ( .A(n10908), .B(n10769), .C(n1826), .Y(n4774) );
  OAI21X1 U11499 ( .A(n10910), .B(n10769), .C(n1384), .Y(n4775) );
  OAI21X1 U11500 ( .A(n10912), .B(n10769), .C(n1510), .Y(n4776) );
  OAI21X1 U11501 ( .A(n10914), .B(n10769), .C(n1134), .Y(n4777) );
  OAI21X1 U11502 ( .A(n10916), .B(n10769), .C(n1259), .Y(n4778) );
  OAI21X1 U11503 ( .A(n10918), .B(n10769), .C(n899), .Y(n4779) );
  OAI21X1 U11504 ( .A(n10920), .B(n10769), .C(n1011), .Y(n4780) );
  OAI21X1 U11505 ( .A(n10922), .B(n10769), .C(n675), .Y(n4781) );
  OAI21X1 U11506 ( .A(n10924), .B(n10769), .C(n787), .Y(n4782) );
  OAI21X1 U11507 ( .A(n10926), .B(n10769), .C(n466), .Y(n4783) );
  OAI21X1 U11508 ( .A(n10928), .B(n10769), .C(n1983), .Y(n4784) );
  OAI21X1 U11509 ( .A(n10930), .B(n10769), .C(n2140), .Y(n4785) );
  OAI21X1 U11510 ( .A(n10932), .B(n10769), .C(n1666), .Y(n4786) );
  OAI21X1 U11511 ( .A(n10934), .B(n10769), .C(n1825), .Y(n4787) );
  OAI21X1 U11512 ( .A(n10936), .B(n10769), .C(n1383), .Y(n4788) );
  OAI21X1 U11513 ( .A(n10938), .B(n10769), .C(n1509), .Y(n4789) );
  OAI21X1 U11514 ( .A(n10940), .B(n10769), .C(n1133), .Y(n4790) );
  OAI21X1 U11515 ( .A(n10942), .B(n10769), .C(n1258), .Y(n4791) );
  OAI21X1 U11516 ( .A(n10944), .B(n10769), .C(n898), .Y(n4792) );
  OAI21X1 U11517 ( .A(n10946), .B(n10769), .C(n1010), .Y(n4793) );
  OAI21X1 U11518 ( .A(n10948), .B(n10769), .C(n674), .Y(n4794) );
  OAI21X1 U11519 ( .A(n10950), .B(n10769), .C(n786), .Y(n4795) );
  OAI21X1 U11520 ( .A(n10954), .B(n10769), .C(n465), .Y(n4796) );
  OAI21X1 U11521 ( .A(n1269), .B(n2153), .C(n10956), .Y(n11245) );
  OAI21X1 U11522 ( .A(n10826), .B(n10771), .C(n1824), .Y(n4797) );
  OAI21X1 U11523 ( .A(n10828), .B(n10771), .C(n1665), .Y(n4798) );
  OAI21X1 U11524 ( .A(n10830), .B(n10771), .C(n2139), .Y(n4799) );
  OAI21X1 U11525 ( .A(n10832), .B(n10771), .C(n1982), .Y(n4800) );
  OAI21X1 U11526 ( .A(n10834), .B(n10771), .C(n1257), .Y(n4801) );
  OAI21X1 U11527 ( .A(n10836), .B(n10771), .C(n1132), .Y(n4802) );
  OAI21X1 U11528 ( .A(n10838), .B(n10771), .C(n1508), .Y(n4803) );
  OAI21X1 U11529 ( .A(n10840), .B(n10771), .C(n1382), .Y(n4804) );
  OAI21X1 U11530 ( .A(n10842), .B(n10771), .C(n785), .Y(n4805) );
  OAI21X1 U11531 ( .A(n10844), .B(n10771), .C(n673), .Y(n4806) );
  OAI21X1 U11532 ( .A(n10846), .B(n10771), .C(n1009), .Y(n4807) );
  OAI21X1 U11533 ( .A(n10848), .B(n10771), .C(n897), .Y(n4808) );
  OAI21X1 U11534 ( .A(n10850), .B(n10771), .C(n1823), .Y(n4809) );
  OAI21X1 U11535 ( .A(n10852), .B(n10771), .C(n1664), .Y(n4810) );
  OAI21X1 U11536 ( .A(n10854), .B(n10771), .C(n2138), .Y(n4811) );
  OAI21X1 U11537 ( .A(n10856), .B(n10771), .C(n1981), .Y(n4812) );
  OAI21X1 U11538 ( .A(n10858), .B(n10771), .C(n1256), .Y(n4813) );
  OAI21X1 U11539 ( .A(n10860), .B(n10771), .C(n1131), .Y(n4814) );
  OAI21X1 U11540 ( .A(n10862), .B(n10771), .C(n1507), .Y(n4815) );
  OAI21X1 U11541 ( .A(n10864), .B(n10771), .C(n1381), .Y(n4816) );
  OAI21X1 U11542 ( .A(n10866), .B(n10771), .C(n784), .Y(n4817) );
  OAI21X1 U11543 ( .A(n10868), .B(n10771), .C(n672), .Y(n4818) );
  OAI21X1 U11544 ( .A(n10870), .B(n10771), .C(n1008), .Y(n4819) );
  OAI21X1 U11545 ( .A(n10872), .B(n10771), .C(n896), .Y(n4820) );
  OAI21X1 U11546 ( .A(n10874), .B(n10771), .C(n361), .Y(n4821) );
  OAI21X1 U11547 ( .A(n10876), .B(n10771), .C(n1822), .Y(n4822) );
  OAI21X1 U11548 ( .A(n10878), .B(n10771), .C(n1663), .Y(n4823) );
  OAI21X1 U11549 ( .A(n10880), .B(n10771), .C(n2137), .Y(n4824) );
  OAI21X1 U11550 ( .A(n10882), .B(n10771), .C(n1980), .Y(n4825) );
  OAI21X1 U11551 ( .A(n10884), .B(n10771), .C(n1255), .Y(n4826) );
  OAI21X1 U11552 ( .A(n10886), .B(n10771), .C(n1130), .Y(n4827) );
  OAI21X1 U11553 ( .A(n10888), .B(n10771), .C(n1506), .Y(n4828) );
  OAI21X1 U11554 ( .A(n10890), .B(n10771), .C(n1380), .Y(n4829) );
  OAI21X1 U11555 ( .A(n10892), .B(n10771), .C(n783), .Y(n4830) );
  OAI21X1 U11556 ( .A(n10894), .B(n10771), .C(n671), .Y(n4831) );
  OAI21X1 U11557 ( .A(n10896), .B(n10771), .C(n1007), .Y(n4832) );
  OAI21X1 U11558 ( .A(n10898), .B(n10771), .C(n895), .Y(n4833) );
  OAI21X1 U11559 ( .A(n10900), .B(n10771), .C(n360), .Y(n4834) );
  OAI21X1 U11560 ( .A(n10902), .B(n10771), .C(n1821), .Y(n4835) );
  OAI21X1 U11561 ( .A(n10904), .B(n10771), .C(n1662), .Y(n4836) );
  OAI21X1 U11562 ( .A(n10906), .B(n10771), .C(n2136), .Y(n4837) );
  OAI21X1 U11563 ( .A(n10908), .B(n10771), .C(n1979), .Y(n4838) );
  OAI21X1 U11564 ( .A(n10910), .B(n10771), .C(n1254), .Y(n4839) );
  OAI21X1 U11565 ( .A(n10912), .B(n10771), .C(n1129), .Y(n4840) );
  OAI21X1 U11566 ( .A(n10914), .B(n10771), .C(n1505), .Y(n4841) );
  OAI21X1 U11567 ( .A(n10916), .B(n10771), .C(n1379), .Y(n4842) );
  OAI21X1 U11568 ( .A(n10918), .B(n10771), .C(n782), .Y(n4843) );
  OAI21X1 U11569 ( .A(n10920), .B(n10771), .C(n670), .Y(n4844) );
  OAI21X1 U11570 ( .A(n10922), .B(n10771), .C(n1006), .Y(n4845) );
  OAI21X1 U11571 ( .A(n10924), .B(n10771), .C(n894), .Y(n4846) );
  OAI21X1 U11572 ( .A(n10926), .B(n10771), .C(n359), .Y(n4847) );
  OAI21X1 U11573 ( .A(n10928), .B(n10771), .C(n1820), .Y(n4848) );
  OAI21X1 U11574 ( .A(n10930), .B(n10771), .C(n1661), .Y(n4849) );
  OAI21X1 U11575 ( .A(n10932), .B(n10771), .C(n2135), .Y(n4850) );
  OAI21X1 U11576 ( .A(n10934), .B(n10771), .C(n1978), .Y(n4851) );
  OAI21X1 U11577 ( .A(n10936), .B(n10771), .C(n1253), .Y(n4852) );
  OAI21X1 U11578 ( .A(n10938), .B(n10771), .C(n1128), .Y(n4853) );
  OAI21X1 U11579 ( .A(n10940), .B(n10771), .C(n1504), .Y(n4854) );
  OAI21X1 U11580 ( .A(n10942), .B(n10771), .C(n1378), .Y(n4855) );
  OAI21X1 U11581 ( .A(n10944), .B(n10771), .C(n781), .Y(n4856) );
  OAI21X1 U11582 ( .A(n10946), .B(n10771), .C(n669), .Y(n4857) );
  OAI21X1 U11583 ( .A(n10948), .B(n10771), .C(n1005), .Y(n4858) );
  OAI21X1 U11584 ( .A(n10950), .B(n10771), .C(n893), .Y(n4859) );
  OAI21X1 U11585 ( .A(n10954), .B(n10771), .C(n358), .Y(n4860) );
  OAI21X1 U11586 ( .A(n1144), .B(n2153), .C(n10956), .Y(n11311) );
  OAI21X1 U11587 ( .A(n10826), .B(n10773), .C(n1660), .Y(n4861) );
  OAI21X1 U11588 ( .A(n10828), .B(n10773), .C(n1819), .Y(n4862) );
  OAI21X1 U11589 ( .A(n10830), .B(n10773), .C(n1977), .Y(n4863) );
  OAI21X1 U11590 ( .A(n10832), .B(n10773), .C(n2134), .Y(n4864) );
  OAI21X1 U11591 ( .A(n10834), .B(n10773), .C(n1127), .Y(n4865) );
  OAI21X1 U11592 ( .A(n10836), .B(n10773), .C(n1252), .Y(n4866) );
  OAI21X1 U11593 ( .A(n10838), .B(n10773), .C(n1377), .Y(n4867) );
  OAI21X1 U11594 ( .A(n10840), .B(n10773), .C(n1503), .Y(n4868) );
  OAI21X1 U11595 ( .A(n10842), .B(n10773), .C(n668), .Y(n4869) );
  OAI21X1 U11596 ( .A(n10844), .B(n10773), .C(n780), .Y(n4870) );
  OAI21X1 U11597 ( .A(n10846), .B(n10773), .C(n892), .Y(n4871) );
  OAI21X1 U11598 ( .A(n10848), .B(n10773), .C(n1004), .Y(n4872) );
  OAI21X1 U11599 ( .A(n10850), .B(n10773), .C(n1659), .Y(n4873) );
  OAI21X1 U11600 ( .A(n10852), .B(n10773), .C(n1818), .Y(n4874) );
  OAI21X1 U11601 ( .A(n10854), .B(n10773), .C(n1976), .Y(n4875) );
  OAI21X1 U11602 ( .A(n10856), .B(n10773), .C(n2133), .Y(n4876) );
  OAI21X1 U11603 ( .A(n10858), .B(n10773), .C(n1126), .Y(n4877) );
  OAI21X1 U11604 ( .A(n10860), .B(n10773), .C(n1251), .Y(n4878) );
  OAI21X1 U11605 ( .A(n10862), .B(n10773), .C(n1376), .Y(n4879) );
  OAI21X1 U11606 ( .A(n10864), .B(n10773), .C(n1502), .Y(n4880) );
  OAI21X1 U11607 ( .A(n10866), .B(n10773), .C(n667), .Y(n4881) );
  OAI21X1 U11608 ( .A(n10868), .B(n10773), .C(n779), .Y(n4882) );
  OAI21X1 U11609 ( .A(n10870), .B(n10773), .C(n891), .Y(n4883) );
  OAI21X1 U11610 ( .A(n10872), .B(n10773), .C(n1003), .Y(n4884) );
  OAI21X1 U11611 ( .A(n10874), .B(n10773), .C(n254), .Y(n4885) );
  OAI21X1 U11612 ( .A(n10876), .B(n10773), .C(n1658), .Y(n4886) );
  OAI21X1 U11613 ( .A(n10878), .B(n10773), .C(n1817), .Y(n4887) );
  OAI21X1 U11614 ( .A(n10880), .B(n10773), .C(n1975), .Y(n4888) );
  OAI21X1 U11615 ( .A(n10882), .B(n10773), .C(n2132), .Y(n4889) );
  OAI21X1 U11616 ( .A(n10884), .B(n10773), .C(n1125), .Y(n4890) );
  OAI21X1 U11617 ( .A(n10886), .B(n10773), .C(n1250), .Y(n4891) );
  OAI21X1 U11618 ( .A(n10888), .B(n10773), .C(n1375), .Y(n4892) );
  OAI21X1 U11619 ( .A(n10890), .B(n10773), .C(n1501), .Y(n4893) );
  OAI21X1 U11620 ( .A(n10892), .B(n10773), .C(n666), .Y(n4894) );
  OAI21X1 U11621 ( .A(n10894), .B(n10773), .C(n778), .Y(n4895) );
  OAI21X1 U11622 ( .A(n10896), .B(n10773), .C(n890), .Y(n4896) );
  OAI21X1 U11623 ( .A(n10898), .B(n10773), .C(n1002), .Y(n4897) );
  OAI21X1 U11624 ( .A(n10900), .B(n10773), .C(n253), .Y(n4898) );
  OAI21X1 U11625 ( .A(n10902), .B(n10773), .C(n1657), .Y(n4899) );
  OAI21X1 U11626 ( .A(n10904), .B(n10773), .C(n1816), .Y(n4900) );
  OAI21X1 U11627 ( .A(n10906), .B(n10773), .C(n1974), .Y(n4901) );
  OAI21X1 U11628 ( .A(n10908), .B(n10773), .C(n2131), .Y(n4902) );
  OAI21X1 U11629 ( .A(n10910), .B(n10773), .C(n1124), .Y(n4903) );
  OAI21X1 U11630 ( .A(n10912), .B(n10773), .C(n1249), .Y(n4904) );
  OAI21X1 U11631 ( .A(n10914), .B(n10773), .C(n1374), .Y(n4905) );
  OAI21X1 U11632 ( .A(n10916), .B(n10773), .C(n1500), .Y(n4906) );
  OAI21X1 U11633 ( .A(n10918), .B(n10773), .C(n665), .Y(n4907) );
  OAI21X1 U11634 ( .A(n10920), .B(n10773), .C(n777), .Y(n4908) );
  OAI21X1 U11635 ( .A(n10922), .B(n10773), .C(n889), .Y(n4909) );
  OAI21X1 U11636 ( .A(n10924), .B(n10773), .C(n1001), .Y(n4910) );
  OAI21X1 U11637 ( .A(n10926), .B(n10773), .C(n252), .Y(n4911) );
  OAI21X1 U11638 ( .A(n10928), .B(n10773), .C(n1656), .Y(n4912) );
  OAI21X1 U11639 ( .A(n10930), .B(n10773), .C(n1815), .Y(n4913) );
  OAI21X1 U11640 ( .A(n10932), .B(n10773), .C(n1973), .Y(n4914) );
  OAI21X1 U11641 ( .A(n10934), .B(n10773), .C(n2130), .Y(n4915) );
  OAI21X1 U11642 ( .A(n10936), .B(n10773), .C(n1123), .Y(n4916) );
  OAI21X1 U11643 ( .A(n10938), .B(n10773), .C(n1248), .Y(n4917) );
  OAI21X1 U11644 ( .A(n10940), .B(n10773), .C(n1373), .Y(n4918) );
  OAI21X1 U11645 ( .A(n10942), .B(n10773), .C(n1499), .Y(n4919) );
  OAI21X1 U11646 ( .A(n10944), .B(n10773), .C(n664), .Y(n4920) );
  OAI21X1 U11647 ( .A(n10946), .B(n10773), .C(n776), .Y(n4921) );
  OAI21X1 U11648 ( .A(n10948), .B(n10773), .C(n888), .Y(n4922) );
  OAI21X1 U11649 ( .A(n10950), .B(n10773), .C(n1000), .Y(n4923) );
  OAI21X1 U11650 ( .A(n10954), .B(n10773), .C(n251), .Y(n4924) );
  OAI21X1 U11651 ( .A(n1143), .B(n2153), .C(n10956), .Y(n11377) );
  OAI21X1 U11652 ( .A(n10826), .B(n10775), .C(n1498), .Y(n4925) );
  OAI21X1 U11653 ( .A(n10828), .B(n10775), .C(n1372), .Y(n4926) );
  OAI21X1 U11654 ( .A(n10830), .B(n10775), .C(n1247), .Y(n4927) );
  OAI21X1 U11655 ( .A(n10832), .B(n10775), .C(n1122), .Y(n4928) );
  OAI21X1 U11656 ( .A(n10834), .B(n10775), .C(n2129), .Y(n4929) );
  OAI21X1 U11657 ( .A(n10836), .B(n10775), .C(n1972), .Y(n4930) );
  OAI21X1 U11658 ( .A(n10838), .B(n10775), .C(n1814), .Y(n4931) );
  OAI21X1 U11659 ( .A(n10840), .B(n10775), .C(n1655), .Y(n4932) );
  OAI21X1 U11660 ( .A(n10842), .B(n10775), .C(n571), .Y(n4933) );
  OAI21X1 U11661 ( .A(n10844), .B(n10775), .C(n464), .Y(n4934) );
  OAI21X1 U11662 ( .A(n10846), .B(n10775), .C(n357), .Y(n4935) );
  OAI21X1 U11663 ( .A(n10848), .B(n10775), .C(n250), .Y(n4936) );
  OAI21X1 U11664 ( .A(n10850), .B(n10775), .C(n1497), .Y(n4937) );
  OAI21X1 U11665 ( .A(n10852), .B(n10775), .C(n1371), .Y(n4938) );
  OAI21X1 U11666 ( .A(n10854), .B(n10775), .C(n1246), .Y(n4939) );
  OAI21X1 U11667 ( .A(n10856), .B(n10775), .C(n1121), .Y(n4940) );
  OAI21X1 U11668 ( .A(n10858), .B(n10775), .C(n2128), .Y(n4941) );
  OAI21X1 U11669 ( .A(n10860), .B(n10775), .C(n1971), .Y(n4942) );
  OAI21X1 U11670 ( .A(n10862), .B(n10775), .C(n1813), .Y(n4943) );
  OAI21X1 U11671 ( .A(n10864), .B(n10775), .C(n1654), .Y(n4944) );
  OAI21X1 U11672 ( .A(n10866), .B(n10775), .C(n570), .Y(n4945) );
  OAI21X1 U11673 ( .A(n10868), .B(n10775), .C(n463), .Y(n4946) );
  OAI21X1 U11674 ( .A(n10870), .B(n10775), .C(n356), .Y(n4947) );
  OAI21X1 U11675 ( .A(n10872), .B(n10775), .C(n249), .Y(n4948) );
  OAI21X1 U11676 ( .A(n10874), .B(n10775), .C(n999), .Y(n4949) );
  OAI21X1 U11677 ( .A(n10876), .B(n10775), .C(n1496), .Y(n4950) );
  OAI21X1 U11678 ( .A(n10878), .B(n10775), .C(n1370), .Y(n4951) );
  OAI21X1 U11679 ( .A(n10880), .B(n10775), .C(n1245), .Y(n4952) );
  OAI21X1 U11680 ( .A(n10882), .B(n10775), .C(n1120), .Y(n4953) );
  OAI21X1 U11681 ( .A(n10884), .B(n10775), .C(n2127), .Y(n4954) );
  OAI21X1 U11682 ( .A(n10886), .B(n10775), .C(n1970), .Y(n4955) );
  OAI21X1 U11683 ( .A(n10888), .B(n10775), .C(n1812), .Y(n4956) );
  OAI21X1 U11684 ( .A(n10890), .B(n10775), .C(n1653), .Y(n4957) );
  OAI21X1 U11685 ( .A(n10892), .B(n10775), .C(n569), .Y(n4958) );
  OAI21X1 U11686 ( .A(n10894), .B(n10775), .C(n462), .Y(n4959) );
  OAI21X1 U11687 ( .A(n10896), .B(n10775), .C(n355), .Y(n4960) );
  OAI21X1 U11688 ( .A(n10898), .B(n10775), .C(n248), .Y(n4961) );
  OAI21X1 U11689 ( .A(n10900), .B(n10775), .C(n998), .Y(n4962) );
  OAI21X1 U11690 ( .A(n10902), .B(n10775), .C(n1495), .Y(n4963) );
  OAI21X1 U11691 ( .A(n10904), .B(n10775), .C(n1369), .Y(n4964) );
  OAI21X1 U11692 ( .A(n10906), .B(n10775), .C(n1244), .Y(n4965) );
  OAI21X1 U11693 ( .A(n10908), .B(n10775), .C(n1119), .Y(n4966) );
  OAI21X1 U11694 ( .A(n10910), .B(n10775), .C(n2126), .Y(n4967) );
  OAI21X1 U11695 ( .A(n10912), .B(n10775), .C(n1969), .Y(n4968) );
  OAI21X1 U11696 ( .A(n10914), .B(n10775), .C(n1811), .Y(n4969) );
  OAI21X1 U11697 ( .A(n10916), .B(n10775), .C(n1652), .Y(n4970) );
  OAI21X1 U11698 ( .A(n10918), .B(n10775), .C(n568), .Y(n4971) );
  OAI21X1 U11699 ( .A(n10920), .B(n10775), .C(n461), .Y(n4972) );
  OAI21X1 U11700 ( .A(n10922), .B(n10775), .C(n354), .Y(n4973) );
  OAI21X1 U11701 ( .A(n10924), .B(n10775), .C(n247), .Y(n4974) );
  OAI21X1 U11702 ( .A(n10926), .B(n10775), .C(n997), .Y(n4975) );
  OAI21X1 U11703 ( .A(n10928), .B(n10775), .C(n1494), .Y(n4976) );
  OAI21X1 U11704 ( .A(n10930), .B(n10775), .C(n1368), .Y(n4977) );
  OAI21X1 U11705 ( .A(n10932), .B(n10775), .C(n1243), .Y(n4978) );
  OAI21X1 U11706 ( .A(n10934), .B(n10775), .C(n1118), .Y(n4979) );
  OAI21X1 U11707 ( .A(n10936), .B(n10775), .C(n2125), .Y(n4980) );
  OAI21X1 U11708 ( .A(n10938), .B(n10775), .C(n1968), .Y(n4981) );
  OAI21X1 U11709 ( .A(n10940), .B(n10775), .C(n1810), .Y(n4982) );
  OAI21X1 U11710 ( .A(n10942), .B(n10775), .C(n1651), .Y(n4983) );
  OAI21X1 U11711 ( .A(n10944), .B(n10775), .C(n567), .Y(n4984) );
  OAI21X1 U11712 ( .A(n10946), .B(n10775), .C(n460), .Y(n4985) );
  OAI21X1 U11713 ( .A(n10948), .B(n10775), .C(n353), .Y(n4986) );
  OAI21X1 U11714 ( .A(n10950), .B(n10775), .C(n246), .Y(n4987) );
  OAI21X1 U11715 ( .A(n10954), .B(n10775), .C(n996), .Y(n4988) );
  OAI21X1 U11716 ( .A(n1268), .B(n2153), .C(n10956), .Y(n11443) );
  OAI21X1 U11717 ( .A(n10826), .B(n10777), .C(n1367), .Y(n4989) );
  OAI21X1 U11718 ( .A(n10828), .B(n10777), .C(n1493), .Y(n4990) );
  OAI21X1 U11719 ( .A(n10830), .B(n10777), .C(n1117), .Y(n4991) );
  OAI21X1 U11720 ( .A(n10832), .B(n10777), .C(n1242), .Y(n4992) );
  OAI21X1 U11721 ( .A(n10834), .B(n10777), .C(n1967), .Y(n4993) );
  OAI21X1 U11722 ( .A(n10836), .B(n10777), .C(n2124), .Y(n4994) );
  OAI21X1 U11723 ( .A(n10838), .B(n10777), .C(n1650), .Y(n4995) );
  OAI21X1 U11724 ( .A(n10840), .B(n10777), .C(n1809), .Y(n4996) );
  OAI21X1 U11725 ( .A(n10842), .B(n10777), .C(n459), .Y(n4997) );
  OAI21X1 U11726 ( .A(n10844), .B(n10777), .C(n566), .Y(n4998) );
  OAI21X1 U11727 ( .A(n10846), .B(n10777), .C(n245), .Y(n4999) );
  OAI21X1 U11728 ( .A(n10848), .B(n10777), .C(n352), .Y(n5000) );
  OAI21X1 U11729 ( .A(n10850), .B(n10777), .C(n1366), .Y(n5001) );
  OAI21X1 U11730 ( .A(n10852), .B(n10777), .C(n1492), .Y(n5002) );
  OAI21X1 U11731 ( .A(n10854), .B(n10777), .C(n1116), .Y(n5003) );
  OAI21X1 U11732 ( .A(n10856), .B(n10777), .C(n1241), .Y(n5004) );
  OAI21X1 U11733 ( .A(n10858), .B(n10777), .C(n1966), .Y(n5005) );
  OAI21X1 U11734 ( .A(n10860), .B(n10777), .C(n2123), .Y(n5006) );
  OAI21X1 U11735 ( .A(n10862), .B(n10777), .C(n1649), .Y(n5007) );
  OAI21X1 U11736 ( .A(n10864), .B(n10777), .C(n1808), .Y(n5008) );
  OAI21X1 U11737 ( .A(n10866), .B(n10777), .C(n458), .Y(n5009) );
  OAI21X1 U11738 ( .A(n10868), .B(n10777), .C(n565), .Y(n5010) );
  OAI21X1 U11739 ( .A(n10870), .B(n10777), .C(n244), .Y(n5011) );
  OAI21X1 U11740 ( .A(n10872), .B(n10777), .C(n351), .Y(n5012) );
  OAI21X1 U11741 ( .A(n10874), .B(n10777), .C(n887), .Y(n5013) );
  OAI21X1 U11742 ( .A(n10876), .B(n10777), .C(n1365), .Y(n5014) );
  OAI21X1 U11743 ( .A(n10878), .B(n10777), .C(n1491), .Y(n5015) );
  OAI21X1 U11744 ( .A(n10880), .B(n10777), .C(n1115), .Y(n5016) );
  OAI21X1 U11745 ( .A(n10882), .B(n10777), .C(n1240), .Y(n5017) );
  OAI21X1 U11746 ( .A(n10884), .B(n10777), .C(n1965), .Y(n5018) );
  OAI21X1 U11747 ( .A(n10886), .B(n10777), .C(n2122), .Y(n5019) );
  OAI21X1 U11748 ( .A(n10888), .B(n10777), .C(n1648), .Y(n5020) );
  OAI21X1 U11749 ( .A(n10890), .B(n10777), .C(n1807), .Y(n5021) );
  OAI21X1 U11750 ( .A(n10892), .B(n10777), .C(n457), .Y(n5022) );
  OAI21X1 U11751 ( .A(n10894), .B(n10777), .C(n564), .Y(n5023) );
  OAI21X1 U11752 ( .A(n10896), .B(n10777), .C(n243), .Y(n5024) );
  OAI21X1 U11753 ( .A(n10898), .B(n10777), .C(n350), .Y(n5025) );
  OAI21X1 U11754 ( .A(n10900), .B(n10777), .C(n886), .Y(n5026) );
  OAI21X1 U11755 ( .A(n10902), .B(n10777), .C(n1364), .Y(n5027) );
  OAI21X1 U11756 ( .A(n10904), .B(n10777), .C(n1490), .Y(n5028) );
  OAI21X1 U11757 ( .A(n10906), .B(n10777), .C(n1114), .Y(n5029) );
  OAI21X1 U11758 ( .A(n10908), .B(n10777), .C(n1239), .Y(n5030) );
  OAI21X1 U11759 ( .A(n10910), .B(n10777), .C(n1964), .Y(n5031) );
  OAI21X1 U11760 ( .A(n10912), .B(n10777), .C(n2121), .Y(n5032) );
  OAI21X1 U11761 ( .A(n10914), .B(n10777), .C(n1647), .Y(n5033) );
  OAI21X1 U11762 ( .A(n10916), .B(n10777), .C(n1806), .Y(n5034) );
  OAI21X1 U11763 ( .A(n10918), .B(n10777), .C(n456), .Y(n5035) );
  OAI21X1 U11764 ( .A(n10920), .B(n10777), .C(n563), .Y(n5036) );
  OAI21X1 U11765 ( .A(n10922), .B(n10777), .C(n242), .Y(n5037) );
  OAI21X1 U11766 ( .A(n10924), .B(n10777), .C(n349), .Y(n5038) );
  OAI21X1 U11767 ( .A(n10926), .B(n10777), .C(n885), .Y(n5039) );
  OAI21X1 U11768 ( .A(n10928), .B(n10777), .C(n1363), .Y(n5040) );
  OAI21X1 U11769 ( .A(n10930), .B(n10777), .C(n1489), .Y(n5041) );
  OAI21X1 U11770 ( .A(n10932), .B(n10777), .C(n1113), .Y(n5042) );
  OAI21X1 U11771 ( .A(n10934), .B(n10777), .C(n1238), .Y(n5043) );
  OAI21X1 U11772 ( .A(n10936), .B(n10777), .C(n1963), .Y(n5044) );
  OAI21X1 U11773 ( .A(n10938), .B(n10777), .C(n2120), .Y(n5045) );
  OAI21X1 U11774 ( .A(n10940), .B(n10777), .C(n1646), .Y(n5046) );
  OAI21X1 U11775 ( .A(n10942), .B(n10777), .C(n1805), .Y(n5047) );
  OAI21X1 U11776 ( .A(n10944), .B(n10777), .C(n455), .Y(n5048) );
  OAI21X1 U11777 ( .A(n10946), .B(n10777), .C(n562), .Y(n5049) );
  OAI21X1 U11778 ( .A(n10948), .B(n10777), .C(n241), .Y(n5050) );
  OAI21X1 U11779 ( .A(n10950), .B(n10777), .C(n348), .Y(n5051) );
  OAI21X1 U11780 ( .A(n10954), .B(n10777), .C(n884), .Y(n5052) );
  OAI21X1 U11781 ( .A(n1394), .B(n2153), .C(n10956), .Y(n11509) );
  OAI21X1 U11782 ( .A(n10826), .B(n10779), .C(n1237), .Y(n5053) );
  OAI21X1 U11783 ( .A(n10828), .B(n10779), .C(n1112), .Y(n5054) );
  OAI21X1 U11784 ( .A(n10830), .B(n10779), .C(n1488), .Y(n5055) );
  OAI21X1 U11785 ( .A(n10832), .B(n10779), .C(n1362), .Y(n5056) );
  OAI21X1 U11786 ( .A(n10834), .B(n10779), .C(n1804), .Y(n5057) );
  OAI21X1 U11787 ( .A(n10836), .B(n10779), .C(n1645), .Y(n5058) );
  OAI21X1 U11788 ( .A(n10838), .B(n10779), .C(n2119), .Y(n5059) );
  OAI21X1 U11789 ( .A(n10840), .B(n10779), .C(n1962), .Y(n5060) );
  OAI21X1 U11790 ( .A(n10842), .B(n10779), .C(n347), .Y(n5061) );
  OAI21X1 U11791 ( .A(n10844), .B(n10779), .C(n240), .Y(n5062) );
  OAI21X1 U11792 ( .A(n10846), .B(n10779), .C(n561), .Y(n5063) );
  OAI21X1 U11793 ( .A(n10848), .B(n10779), .C(n454), .Y(n5064) );
  OAI21X1 U11794 ( .A(n10850), .B(n10779), .C(n1236), .Y(n5065) );
  OAI21X1 U11795 ( .A(n10852), .B(n10779), .C(n1111), .Y(n5066) );
  OAI21X1 U11796 ( .A(n10854), .B(n10779), .C(n1487), .Y(n5067) );
  OAI21X1 U11797 ( .A(n10856), .B(n10779), .C(n1361), .Y(n5068) );
  OAI21X1 U11798 ( .A(n10858), .B(n10779), .C(n1803), .Y(n5069) );
  OAI21X1 U11799 ( .A(n10860), .B(n10779), .C(n1644), .Y(n5070) );
  OAI21X1 U11800 ( .A(n10862), .B(n10779), .C(n2118), .Y(n5071) );
  OAI21X1 U11801 ( .A(n10864), .B(n10779), .C(n1961), .Y(n5072) );
  OAI21X1 U11802 ( .A(n10866), .B(n10779), .C(n346), .Y(n5073) );
  OAI21X1 U11803 ( .A(n10868), .B(n10779), .C(n239), .Y(n5074) );
  OAI21X1 U11804 ( .A(n10870), .B(n10779), .C(n560), .Y(n5075) );
  OAI21X1 U11805 ( .A(n10872), .B(n10779), .C(n453), .Y(n5076) );
  OAI21X1 U11806 ( .A(n10874), .B(n10779), .C(n775), .Y(n5077) );
  OAI21X1 U11807 ( .A(n10876), .B(n10779), .C(n1235), .Y(n5078) );
  OAI21X1 U11808 ( .A(n10878), .B(n10779), .C(n1110), .Y(n5079) );
  OAI21X1 U11809 ( .A(n10880), .B(n10779), .C(n1486), .Y(n5080) );
  OAI21X1 U11810 ( .A(n10882), .B(n10779), .C(n1360), .Y(n5081) );
  OAI21X1 U11811 ( .A(n10884), .B(n10779), .C(n1802), .Y(n5082) );
  OAI21X1 U11812 ( .A(n10886), .B(n10779), .C(n1643), .Y(n5083) );
  OAI21X1 U11813 ( .A(n10888), .B(n10779), .C(n2117), .Y(n5084) );
  OAI21X1 U11814 ( .A(n10890), .B(n10779), .C(n1960), .Y(n5085) );
  OAI21X1 U11815 ( .A(n10892), .B(n10779), .C(n345), .Y(n5086) );
  OAI21X1 U11816 ( .A(n10894), .B(n10779), .C(n238), .Y(n5087) );
  OAI21X1 U11817 ( .A(n10896), .B(n10779), .C(n559), .Y(n5088) );
  OAI21X1 U11818 ( .A(n10898), .B(n10779), .C(n452), .Y(n5089) );
  OAI21X1 U11819 ( .A(n10900), .B(n10779), .C(n774), .Y(n5090) );
  OAI21X1 U11820 ( .A(n10902), .B(n10779), .C(n1234), .Y(n5091) );
  OAI21X1 U11821 ( .A(n10904), .B(n10779), .C(n1109), .Y(n5092) );
  OAI21X1 U11822 ( .A(n10906), .B(n10779), .C(n1485), .Y(n5093) );
  OAI21X1 U11823 ( .A(n10908), .B(n10779), .C(n1359), .Y(n5094) );
  OAI21X1 U11824 ( .A(n10910), .B(n10779), .C(n1801), .Y(n5095) );
  OAI21X1 U11825 ( .A(n10912), .B(n10779), .C(n1642), .Y(n5096) );
  OAI21X1 U11826 ( .A(n10914), .B(n10779), .C(n2116), .Y(n5097) );
  OAI21X1 U11827 ( .A(n10916), .B(n10779), .C(n1959), .Y(n5098) );
  OAI21X1 U11828 ( .A(n10918), .B(n10779), .C(n344), .Y(n5099) );
  OAI21X1 U11829 ( .A(n10920), .B(n10779), .C(n237), .Y(n5100) );
  OAI21X1 U11830 ( .A(n10922), .B(n10779), .C(n558), .Y(n5101) );
  OAI21X1 U11831 ( .A(n10924), .B(n10779), .C(n451), .Y(n5102) );
  OAI21X1 U11832 ( .A(n10926), .B(n10779), .C(n773), .Y(n5103) );
  OAI21X1 U11833 ( .A(n10928), .B(n10779), .C(n1233), .Y(n5104) );
  OAI21X1 U11834 ( .A(n10930), .B(n10779), .C(n1108), .Y(n5105) );
  OAI21X1 U11835 ( .A(n10932), .B(n10779), .C(n1484), .Y(n5106) );
  OAI21X1 U11836 ( .A(n10934), .B(n10779), .C(n1358), .Y(n5107) );
  OAI21X1 U11837 ( .A(n10936), .B(n10779), .C(n1800), .Y(n5108) );
  OAI21X1 U11838 ( .A(n10938), .B(n10779), .C(n1641), .Y(n5109) );
  OAI21X1 U11839 ( .A(n10940), .B(n10779), .C(n2115), .Y(n5110) );
  OAI21X1 U11840 ( .A(n10942), .B(n10779), .C(n1958), .Y(n5111) );
  OAI21X1 U11841 ( .A(n10944), .B(n10779), .C(n343), .Y(n5112) );
  OAI21X1 U11842 ( .A(n10946), .B(n10779), .C(n236), .Y(n5113) );
  OAI21X1 U11843 ( .A(n10948), .B(n10779), .C(n557), .Y(n5114) );
  OAI21X1 U11844 ( .A(n10950), .B(n10779), .C(n450), .Y(n5115) );
  OAI21X1 U11845 ( .A(n10954), .B(n10779), .C(n772), .Y(n5116) );
  OAI21X1 U11846 ( .A(n1678), .B(n2153), .C(n10956), .Y(n11576) );
  OAI21X1 U11847 ( .A(n10826), .B(n10781), .C(n1107), .Y(n5117) );
  OAI21X1 U11848 ( .A(n10828), .B(n10781), .C(n1232), .Y(n5118) );
  OAI21X1 U11849 ( .A(n10830), .B(n10781), .C(n1357), .Y(n5119) );
  OAI21X1 U11850 ( .A(n10832), .B(n10781), .C(n1483), .Y(n5120) );
  OAI21X1 U11851 ( .A(n10834), .B(n10781), .C(n1640), .Y(n5121) );
  OAI21X1 U11852 ( .A(n10836), .B(n10781), .C(n1799), .Y(n5122) );
  OAI21X1 U11853 ( .A(n10838), .B(n10781), .C(n1957), .Y(n5123) );
  OAI21X1 U11854 ( .A(n10840), .B(n10781), .C(n2114), .Y(n5124) );
  OAI21X1 U11855 ( .A(n10842), .B(n10781), .C(n235), .Y(n5125) );
  OAI21X1 U11856 ( .A(n10844), .B(n10781), .C(n342), .Y(n5126) );
  OAI21X1 U11857 ( .A(n10846), .B(n10781), .C(n449), .Y(n5127) );
  OAI21X1 U11858 ( .A(n10848), .B(n10781), .C(n556), .Y(n5128) );
  OAI21X1 U11859 ( .A(n10850), .B(n10781), .C(n1106), .Y(n5129) );
  OAI21X1 U11860 ( .A(n10852), .B(n10781), .C(n1231), .Y(n5130) );
  OAI21X1 U11861 ( .A(n10854), .B(n10781), .C(n1356), .Y(n5131) );
  OAI21X1 U11862 ( .A(n10856), .B(n10781), .C(n1482), .Y(n5132) );
  OAI21X1 U11863 ( .A(n10858), .B(n10781), .C(n1639), .Y(n5133) );
  OAI21X1 U11864 ( .A(n10860), .B(n10781), .C(n1798), .Y(n5134) );
  OAI21X1 U11865 ( .A(n10862), .B(n10781), .C(n1956), .Y(n5135) );
  OAI21X1 U11866 ( .A(n10864), .B(n10781), .C(n2113), .Y(n5136) );
  OAI21X1 U11867 ( .A(n10866), .B(n10781), .C(n234), .Y(n5137) );
  OAI21X1 U11868 ( .A(n10868), .B(n10781), .C(n341), .Y(n5138) );
  OAI21X1 U11869 ( .A(n10870), .B(n10781), .C(n448), .Y(n5139) );
  OAI21X1 U11870 ( .A(n10872), .B(n10781), .C(n555), .Y(n5140) );
  OAI21X1 U11871 ( .A(n10874), .B(n10781), .C(n663), .Y(n5141) );
  OAI21X1 U11872 ( .A(n10876), .B(n10781), .C(n1105), .Y(n5142) );
  OAI21X1 U11873 ( .A(n10878), .B(n10781), .C(n1230), .Y(n5143) );
  OAI21X1 U11874 ( .A(n10880), .B(n10781), .C(n1355), .Y(n5144) );
  OAI21X1 U11875 ( .A(n10882), .B(n10781), .C(n1481), .Y(n5145) );
  OAI21X1 U11876 ( .A(n10884), .B(n10781), .C(n1638), .Y(n5146) );
  OAI21X1 U11877 ( .A(n10886), .B(n10781), .C(n1797), .Y(n5147) );
  OAI21X1 U11878 ( .A(n10888), .B(n10781), .C(n1955), .Y(n5148) );
  OAI21X1 U11879 ( .A(n10890), .B(n10781), .C(n2112), .Y(n5149) );
  OAI21X1 U11880 ( .A(n10892), .B(n10781), .C(n233), .Y(n5150) );
  OAI21X1 U11881 ( .A(n10894), .B(n10781), .C(n340), .Y(n5151) );
  OAI21X1 U11882 ( .A(n10896), .B(n10781), .C(n447), .Y(n5152) );
  OAI21X1 U11883 ( .A(n10898), .B(n10781), .C(n554), .Y(n5153) );
  OAI21X1 U11884 ( .A(n10900), .B(n10781), .C(n662), .Y(n5154) );
  OAI21X1 U11885 ( .A(n10902), .B(n10781), .C(n1104), .Y(n5155) );
  OAI21X1 U11886 ( .A(n10904), .B(n10781), .C(n1229), .Y(n5156) );
  OAI21X1 U11887 ( .A(n10906), .B(n10781), .C(n1354), .Y(n5157) );
  OAI21X1 U11888 ( .A(n10908), .B(n10781), .C(n1480), .Y(n5158) );
  OAI21X1 U11889 ( .A(n10910), .B(n10781), .C(n1637), .Y(n5159) );
  OAI21X1 U11890 ( .A(n10912), .B(n10781), .C(n1796), .Y(n5160) );
  OAI21X1 U11891 ( .A(n10914), .B(n10781), .C(n1954), .Y(n5161) );
  OAI21X1 U11892 ( .A(n10916), .B(n10781), .C(n2111), .Y(n5162) );
  OAI21X1 U11893 ( .A(n10918), .B(n10781), .C(n232), .Y(n5163) );
  OAI21X1 U11894 ( .A(n10920), .B(n10781), .C(n339), .Y(n5164) );
  OAI21X1 U11895 ( .A(n10922), .B(n10781), .C(n446), .Y(n5165) );
  OAI21X1 U11896 ( .A(n10924), .B(n10781), .C(n553), .Y(n5166) );
  OAI21X1 U11897 ( .A(n10926), .B(n10781), .C(n661), .Y(n5167) );
  OAI21X1 U11898 ( .A(n10928), .B(n10781), .C(n1103), .Y(n5168) );
  OAI21X1 U11899 ( .A(n10930), .B(n10781), .C(n1228), .Y(n5169) );
  OAI21X1 U11900 ( .A(n10932), .B(n10781), .C(n1353), .Y(n5170) );
  OAI21X1 U11901 ( .A(n10934), .B(n10781), .C(n1479), .Y(n5171) );
  OAI21X1 U11902 ( .A(n10936), .B(n10781), .C(n1636), .Y(n5172) );
  OAI21X1 U11903 ( .A(n10938), .B(n10781), .C(n1795), .Y(n5173) );
  OAI21X1 U11904 ( .A(n10940), .B(n10781), .C(n1953), .Y(n5174) );
  OAI21X1 U11905 ( .A(n10942), .B(n10781), .C(n2110), .Y(n5175) );
  OAI21X1 U11906 ( .A(n10944), .B(n10781), .C(n231), .Y(n5176) );
  OAI21X1 U11907 ( .A(n10946), .B(n10781), .C(n338), .Y(n5177) );
  OAI21X1 U11908 ( .A(n10948), .B(n10781), .C(n445), .Y(n5178) );
  OAI21X1 U11909 ( .A(n10950), .B(n10781), .C(n552), .Y(n5179) );
  OAI21X1 U11910 ( .A(n10954), .B(n10781), .C(n660), .Y(n5180) );
  NAND3X1 U11911 ( .A(n4152), .B(n10964), .C(n11112), .Y(n12104) );
  OAI21X1 U11912 ( .A(n1520), .B(n1994), .C(n10956), .Y(n11642) );
  OAI21X1 U11913 ( .A(n10826), .B(n10783), .C(n995), .Y(n5181) );
  OAI21X1 U11914 ( .A(n10828), .B(n10783), .C(n883), .Y(n5182) );
  OAI21X1 U11915 ( .A(n10830), .B(n10783), .C(n771), .Y(n5183) );
  OAI21X1 U11916 ( .A(n10832), .B(n10783), .C(n659), .Y(n5184) );
  OAI21X1 U11917 ( .A(n10834), .B(n10783), .C(n551), .Y(n5185) );
  OAI21X1 U11918 ( .A(n10836), .B(n10783), .C(n444), .Y(n5186) );
  OAI21X1 U11919 ( .A(n10838), .B(n10783), .C(n337), .Y(n5187) );
  OAI21X1 U11920 ( .A(n10840), .B(n10783), .C(n230), .Y(n5188) );
  OAI21X1 U11921 ( .A(n10842), .B(n10783), .C(n2109), .Y(n5189) );
  OAI21X1 U11922 ( .A(n10844), .B(n10783), .C(n1952), .Y(n5190) );
  OAI21X1 U11923 ( .A(n10846), .B(n10783), .C(n1794), .Y(n5191) );
  OAI21X1 U11924 ( .A(n10848), .B(n10783), .C(n1635), .Y(n5192) );
  OAI21X1 U11925 ( .A(n10850), .B(n10783), .C(n994), .Y(n5193) );
  OAI21X1 U11926 ( .A(n10852), .B(n10783), .C(n882), .Y(n5194) );
  OAI21X1 U11927 ( .A(n10854), .B(n10783), .C(n770), .Y(n5195) );
  OAI21X1 U11928 ( .A(n10856), .B(n10783), .C(n658), .Y(n5196) );
  OAI21X1 U11929 ( .A(n10858), .B(n10783), .C(n550), .Y(n5197) );
  OAI21X1 U11930 ( .A(n10860), .B(n10783), .C(n443), .Y(n5198) );
  OAI21X1 U11931 ( .A(n10862), .B(n10783), .C(n336), .Y(n5199) );
  OAI21X1 U11932 ( .A(n10864), .B(n10783), .C(n229), .Y(n5200) );
  OAI21X1 U11933 ( .A(n10866), .B(n10783), .C(n2108), .Y(n5201) );
  OAI21X1 U11934 ( .A(n10868), .B(n10783), .C(n1951), .Y(n5202) );
  OAI21X1 U11935 ( .A(n10870), .B(n10783), .C(n1793), .Y(n5203) );
  OAI21X1 U11936 ( .A(n10872), .B(n10783), .C(n1634), .Y(n5204) );
  OAI21X1 U11937 ( .A(n10874), .B(n10783), .C(n1478), .Y(n5205) );
  OAI21X1 U11938 ( .A(n10876), .B(n10783), .C(n993), .Y(n5206) );
  OAI21X1 U11939 ( .A(n10878), .B(n10783), .C(n881), .Y(n5207) );
  OAI21X1 U11940 ( .A(n10880), .B(n10783), .C(n769), .Y(n5208) );
  OAI21X1 U11941 ( .A(n10882), .B(n10783), .C(n657), .Y(n5209) );
  OAI21X1 U11942 ( .A(n10884), .B(n10783), .C(n549), .Y(n5210) );
  OAI21X1 U11943 ( .A(n10886), .B(n10783), .C(n442), .Y(n5211) );
  OAI21X1 U11944 ( .A(n10888), .B(n10783), .C(n335), .Y(n5212) );
  OAI21X1 U11945 ( .A(n10890), .B(n10783), .C(n228), .Y(n5213) );
  OAI21X1 U11946 ( .A(n10892), .B(n10783), .C(n2107), .Y(n5214) );
  OAI21X1 U11947 ( .A(n10894), .B(n10783), .C(n1950), .Y(n5215) );
  OAI21X1 U11948 ( .A(n10896), .B(n10783), .C(n1792), .Y(n5216) );
  OAI21X1 U11949 ( .A(n10898), .B(n10783), .C(n1633), .Y(n5217) );
  OAI21X1 U11950 ( .A(n10900), .B(n10783), .C(n1477), .Y(n5218) );
  OAI21X1 U11951 ( .A(n10902), .B(n10783), .C(n992), .Y(n5219) );
  OAI21X1 U11952 ( .A(n10904), .B(n10783), .C(n880), .Y(n5220) );
  OAI21X1 U11953 ( .A(n10906), .B(n10783), .C(n768), .Y(n5221) );
  OAI21X1 U11954 ( .A(n10908), .B(n10783), .C(n656), .Y(n5222) );
  OAI21X1 U11955 ( .A(n10910), .B(n10783), .C(n548), .Y(n5223) );
  OAI21X1 U11956 ( .A(n10912), .B(n10783), .C(n441), .Y(n5224) );
  OAI21X1 U11957 ( .A(n10914), .B(n10783), .C(n334), .Y(n5225) );
  OAI21X1 U11958 ( .A(n10916), .B(n10783), .C(n227), .Y(n5226) );
  OAI21X1 U11959 ( .A(n10918), .B(n10783), .C(n2106), .Y(n5227) );
  OAI21X1 U11960 ( .A(n10920), .B(n10783), .C(n1949), .Y(n5228) );
  OAI21X1 U11961 ( .A(n10922), .B(n10783), .C(n1791), .Y(n5229) );
  OAI21X1 U11962 ( .A(n10924), .B(n10783), .C(n1632), .Y(n5230) );
  OAI21X1 U11963 ( .A(n10926), .B(n10783), .C(n1476), .Y(n5231) );
  OAI21X1 U11964 ( .A(n10928), .B(n10783), .C(n991), .Y(n5232) );
  OAI21X1 U11965 ( .A(n10930), .B(n10783), .C(n879), .Y(n5233) );
  OAI21X1 U11966 ( .A(n10932), .B(n10783), .C(n767), .Y(n5234) );
  OAI21X1 U11967 ( .A(n10934), .B(n10783), .C(n655), .Y(n5235) );
  OAI21X1 U11968 ( .A(n10936), .B(n10783), .C(n547), .Y(n5236) );
  OAI21X1 U11969 ( .A(n10938), .B(n10783), .C(n440), .Y(n5237) );
  OAI21X1 U11970 ( .A(n10940), .B(n10783), .C(n333), .Y(n5238) );
  OAI21X1 U11971 ( .A(n10942), .B(n10783), .C(n226), .Y(n5239) );
  OAI21X1 U11972 ( .A(n10944), .B(n10783), .C(n2105), .Y(n5240) );
  OAI21X1 U11973 ( .A(n10946), .B(n10783), .C(n1948), .Y(n5241) );
  OAI21X1 U11974 ( .A(n10948), .B(n10783), .C(n1790), .Y(n5242) );
  OAI21X1 U11975 ( .A(n10950), .B(n10783), .C(n1631), .Y(n5243) );
  OAI21X1 U11976 ( .A(n10954), .B(n10783), .C(n1475), .Y(n5244) );
  OAI21X1 U11977 ( .A(n1395), .B(n1994), .C(n10956), .Y(n11708) );
  OAI21X1 U11978 ( .A(n10826), .B(n10785), .C(n878), .Y(n5245) );
  OAI21X1 U11979 ( .A(n10828), .B(n10785), .C(n990), .Y(n5246) );
  OAI21X1 U11980 ( .A(n10830), .B(n10785), .C(n654), .Y(n5247) );
  OAI21X1 U11981 ( .A(n10832), .B(n10785), .C(n766), .Y(n5248) );
  OAI21X1 U11982 ( .A(n10834), .B(n10785), .C(n439), .Y(n5249) );
  OAI21X1 U11983 ( .A(n10836), .B(n10785), .C(n546), .Y(n5250) );
  OAI21X1 U11984 ( .A(n10838), .B(n10785), .C(n225), .Y(n5251) );
  OAI21X1 U11985 ( .A(n10840), .B(n10785), .C(n332), .Y(n5252) );
  OAI21X1 U11986 ( .A(n10842), .B(n10785), .C(n1947), .Y(n5253) );
  OAI21X1 U11987 ( .A(n10844), .B(n10785), .C(n2104), .Y(n5254) );
  OAI21X1 U11988 ( .A(n10846), .B(n10785), .C(n1630), .Y(n5255) );
  OAI21X1 U11989 ( .A(n10848), .B(n10785), .C(n1789), .Y(n5256) );
  OAI21X1 U11990 ( .A(n10850), .B(n10785), .C(n877), .Y(n5257) );
  OAI21X1 U11991 ( .A(n10852), .B(n10785), .C(n989), .Y(n5258) );
  OAI21X1 U11992 ( .A(n10854), .B(n10785), .C(n653), .Y(n5259) );
  OAI21X1 U11993 ( .A(n10856), .B(n10785), .C(n765), .Y(n5260) );
  OAI21X1 U11994 ( .A(n10858), .B(n10785), .C(n438), .Y(n5261) );
  OAI21X1 U11995 ( .A(n10860), .B(n10785), .C(n545), .Y(n5262) );
  OAI21X1 U11996 ( .A(n10862), .B(n10785), .C(n224), .Y(n5263) );
  OAI21X1 U11997 ( .A(n10864), .B(n10785), .C(n331), .Y(n5264) );
  OAI21X1 U11998 ( .A(n10866), .B(n10785), .C(n1946), .Y(n5265) );
  OAI21X1 U11999 ( .A(n10868), .B(n10785), .C(n2103), .Y(n5266) );
  OAI21X1 U12000 ( .A(n10870), .B(n10785), .C(n1629), .Y(n5267) );
  OAI21X1 U12001 ( .A(n10872), .B(n10785), .C(n1788), .Y(n5268) );
  OAI21X1 U12002 ( .A(n10874), .B(n10785), .C(n1352), .Y(n5269) );
  OAI21X1 U12003 ( .A(n10876), .B(n10785), .C(n876), .Y(n5270) );
  OAI21X1 U12004 ( .A(n10878), .B(n10785), .C(n988), .Y(n5271) );
  OAI21X1 U12005 ( .A(n10880), .B(n10785), .C(n652), .Y(n5272) );
  OAI21X1 U12006 ( .A(n10882), .B(n10785), .C(n764), .Y(n5273) );
  OAI21X1 U12007 ( .A(n10884), .B(n10785), .C(n437), .Y(n5274) );
  OAI21X1 U12008 ( .A(n10886), .B(n10785), .C(n544), .Y(n5275) );
  OAI21X1 U12009 ( .A(n10888), .B(n10785), .C(n223), .Y(n5276) );
  OAI21X1 U12010 ( .A(n10890), .B(n10785), .C(n330), .Y(n5277) );
  OAI21X1 U12011 ( .A(n10892), .B(n10785), .C(n1945), .Y(n5278) );
  OAI21X1 U12012 ( .A(n10894), .B(n10785), .C(n2102), .Y(n5279) );
  OAI21X1 U12013 ( .A(n10896), .B(n10785), .C(n1628), .Y(n5280) );
  OAI21X1 U12014 ( .A(n10898), .B(n10785), .C(n1787), .Y(n5281) );
  OAI21X1 U12015 ( .A(n10900), .B(n10785), .C(n1351), .Y(n5282) );
  OAI21X1 U12016 ( .A(n10902), .B(n10785), .C(n875), .Y(n5283) );
  OAI21X1 U12017 ( .A(n10904), .B(n10785), .C(n987), .Y(n5284) );
  OAI21X1 U12018 ( .A(n10906), .B(n10785), .C(n651), .Y(n5285) );
  OAI21X1 U12019 ( .A(n10908), .B(n10785), .C(n763), .Y(n5286) );
  OAI21X1 U12020 ( .A(n10910), .B(n10785), .C(n436), .Y(n5287) );
  OAI21X1 U12021 ( .A(n10912), .B(n10785), .C(n543), .Y(n5288) );
  OAI21X1 U12022 ( .A(n10914), .B(n10785), .C(n222), .Y(n5289) );
  OAI21X1 U12023 ( .A(n10916), .B(n10785), .C(n329), .Y(n5290) );
  OAI21X1 U12024 ( .A(n10918), .B(n10785), .C(n1944), .Y(n5291) );
  OAI21X1 U12025 ( .A(n10920), .B(n10785), .C(n2101), .Y(n5292) );
  OAI21X1 U12026 ( .A(n10922), .B(n10785), .C(n1627), .Y(n5293) );
  OAI21X1 U12027 ( .A(n10924), .B(n10785), .C(n1786), .Y(n5294) );
  OAI21X1 U12028 ( .A(n10926), .B(n10785), .C(n1350), .Y(n5295) );
  OAI21X1 U12029 ( .A(n10928), .B(n10785), .C(n874), .Y(n5296) );
  OAI21X1 U12030 ( .A(n10930), .B(n10785), .C(n986), .Y(n5297) );
  OAI21X1 U12031 ( .A(n10932), .B(n10785), .C(n650), .Y(n5298) );
  OAI21X1 U12032 ( .A(n10934), .B(n10785), .C(n762), .Y(n5299) );
  OAI21X1 U12033 ( .A(n10936), .B(n10785), .C(n435), .Y(n5300) );
  OAI21X1 U12034 ( .A(n10938), .B(n10785), .C(n542), .Y(n5301) );
  OAI21X1 U12035 ( .A(n10940), .B(n10785), .C(n221), .Y(n5302) );
  OAI21X1 U12036 ( .A(n10942), .B(n10785), .C(n328), .Y(n5303) );
  OAI21X1 U12037 ( .A(n10944), .B(n10785), .C(n1943), .Y(n5304) );
  OAI21X1 U12038 ( .A(n10946), .B(n10785), .C(n2100), .Y(n5305) );
  OAI21X1 U12039 ( .A(n10948), .B(n10785), .C(n1626), .Y(n5306) );
  OAI21X1 U12040 ( .A(n10950), .B(n10785), .C(n1785), .Y(n5307) );
  OAI21X1 U12041 ( .A(n10954), .B(n10785), .C(n1349), .Y(n5308) );
  OAI21X1 U12042 ( .A(n1269), .B(n1994), .C(n10956), .Y(n11774) );
  OAI21X1 U12043 ( .A(n10826), .B(n10787), .C(n761), .Y(n5309) );
  OAI21X1 U12044 ( .A(n10828), .B(n10787), .C(n649), .Y(n5310) );
  OAI21X1 U12045 ( .A(n10830), .B(n10787), .C(n985), .Y(n5311) );
  OAI21X1 U12046 ( .A(n10832), .B(n10787), .C(n873), .Y(n5312) );
  OAI21X1 U12047 ( .A(n10834), .B(n10787), .C(n327), .Y(n5313) );
  OAI21X1 U12048 ( .A(n10836), .B(n10787), .C(n220), .Y(n5314) );
  OAI21X1 U12049 ( .A(n10838), .B(n10787), .C(n541), .Y(n5315) );
  OAI21X1 U12050 ( .A(n10840), .B(n10787), .C(n434), .Y(n5316) );
  OAI21X1 U12051 ( .A(n10842), .B(n10787), .C(n1784), .Y(n5317) );
  OAI21X1 U12052 ( .A(n10844), .B(n10787), .C(n1625), .Y(n5318) );
  OAI21X1 U12053 ( .A(n10846), .B(n10787), .C(n2099), .Y(n5319) );
  OAI21X1 U12054 ( .A(n10848), .B(n10787), .C(n1942), .Y(n5320) );
  OAI21X1 U12055 ( .A(n10850), .B(n10787), .C(n760), .Y(n5321) );
  OAI21X1 U12056 ( .A(n10852), .B(n10787), .C(n648), .Y(n5322) );
  OAI21X1 U12057 ( .A(n10854), .B(n10787), .C(n984), .Y(n5323) );
  OAI21X1 U12058 ( .A(n10856), .B(n10787), .C(n872), .Y(n5324) );
  OAI21X1 U12059 ( .A(n10858), .B(n10787), .C(n326), .Y(n5325) );
  OAI21X1 U12060 ( .A(n10860), .B(n10787), .C(n219), .Y(n5326) );
  OAI21X1 U12061 ( .A(n10862), .B(n10787), .C(n540), .Y(n5327) );
  OAI21X1 U12062 ( .A(n10864), .B(n10787), .C(n433), .Y(n5328) );
  OAI21X1 U12063 ( .A(n10866), .B(n10787), .C(n1783), .Y(n5329) );
  OAI21X1 U12064 ( .A(n10868), .B(n10787), .C(n1624), .Y(n5330) );
  OAI21X1 U12065 ( .A(n10870), .B(n10787), .C(n2098), .Y(n5331) );
  OAI21X1 U12066 ( .A(n10872), .B(n10787), .C(n1941), .Y(n5332) );
  OAI21X1 U12067 ( .A(n10874), .B(n10787), .C(n1227), .Y(n5333) );
  OAI21X1 U12068 ( .A(n10876), .B(n10787), .C(n759), .Y(n5334) );
  OAI21X1 U12069 ( .A(n10878), .B(n10787), .C(n647), .Y(n5335) );
  OAI21X1 U12070 ( .A(n10880), .B(n10787), .C(n983), .Y(n5336) );
  OAI21X1 U12071 ( .A(n10882), .B(n10787), .C(n871), .Y(n5337) );
  OAI21X1 U12072 ( .A(n10884), .B(n10787), .C(n325), .Y(n5338) );
  OAI21X1 U12073 ( .A(n10886), .B(n10787), .C(n218), .Y(n5339) );
  OAI21X1 U12074 ( .A(n10888), .B(n10787), .C(n539), .Y(n5340) );
  OAI21X1 U12075 ( .A(n10890), .B(n10787), .C(n432), .Y(n5341) );
  OAI21X1 U12076 ( .A(n10892), .B(n10787), .C(n1782), .Y(n5342) );
  OAI21X1 U12077 ( .A(n10894), .B(n10787), .C(n1623), .Y(n5343) );
  OAI21X1 U12078 ( .A(n10896), .B(n10787), .C(n2097), .Y(n5344) );
  OAI21X1 U12079 ( .A(n10898), .B(n10787), .C(n1940), .Y(n5345) );
  OAI21X1 U12080 ( .A(n10900), .B(n10787), .C(n1226), .Y(n5346) );
  OAI21X1 U12081 ( .A(n10902), .B(n10787), .C(n758), .Y(n5347) );
  OAI21X1 U12082 ( .A(n10904), .B(n10787), .C(n646), .Y(n5348) );
  OAI21X1 U12083 ( .A(n10906), .B(n10787), .C(n982), .Y(n5349) );
  OAI21X1 U12084 ( .A(n10908), .B(n10787), .C(n870), .Y(n5350) );
  OAI21X1 U12085 ( .A(n10910), .B(n10787), .C(n324), .Y(n5351) );
  OAI21X1 U12086 ( .A(n10912), .B(n10787), .C(n217), .Y(n5352) );
  OAI21X1 U12087 ( .A(n10914), .B(n10787), .C(n538), .Y(n5353) );
  OAI21X1 U12088 ( .A(n10916), .B(n10787), .C(n431), .Y(n5354) );
  OAI21X1 U12089 ( .A(n10918), .B(n10787), .C(n1781), .Y(n5355) );
  OAI21X1 U12090 ( .A(n10920), .B(n10787), .C(n1622), .Y(n5356) );
  OAI21X1 U12091 ( .A(n10922), .B(n10787), .C(n2096), .Y(n5357) );
  OAI21X1 U12092 ( .A(n10924), .B(n10787), .C(n1939), .Y(n5358) );
  OAI21X1 U12093 ( .A(n10926), .B(n10787), .C(n1225), .Y(n5359) );
  OAI21X1 U12094 ( .A(n10928), .B(n10787), .C(n757), .Y(n5360) );
  OAI21X1 U12095 ( .A(n10930), .B(n10787), .C(n645), .Y(n5361) );
  OAI21X1 U12096 ( .A(n10932), .B(n10787), .C(n981), .Y(n5362) );
  OAI21X1 U12097 ( .A(n10934), .B(n10787), .C(n869), .Y(n5363) );
  OAI21X1 U12098 ( .A(n10936), .B(n10787), .C(n323), .Y(n5364) );
  OAI21X1 U12099 ( .A(n10938), .B(n10787), .C(n216), .Y(n5365) );
  OAI21X1 U12100 ( .A(n10940), .B(n10787), .C(n537), .Y(n5366) );
  OAI21X1 U12101 ( .A(n10942), .B(n10787), .C(n430), .Y(n5367) );
  OAI21X1 U12102 ( .A(n10944), .B(n10787), .C(n1780), .Y(n5368) );
  OAI21X1 U12103 ( .A(n10946), .B(n10787), .C(n1621), .Y(n5369) );
  OAI21X1 U12104 ( .A(n10948), .B(n10787), .C(n2095), .Y(n5370) );
  OAI21X1 U12105 ( .A(n10950), .B(n10787), .C(n1938), .Y(n5371) );
  OAI21X1 U12106 ( .A(n10954), .B(n10787), .C(n1224), .Y(n5372) );
  OAI21X1 U12107 ( .A(n1144), .B(n1994), .C(n10956), .Y(n11840) );
  OAI21X1 U12108 ( .A(n10826), .B(n10789), .C(n644), .Y(n5373) );
  OAI21X1 U12109 ( .A(n10828), .B(n10789), .C(n756), .Y(n5374) );
  OAI21X1 U12110 ( .A(n10830), .B(n10789), .C(n868), .Y(n5375) );
  OAI21X1 U12111 ( .A(n10832), .B(n10789), .C(n980), .Y(n5376) );
  OAI21X1 U12112 ( .A(n10834), .B(n10789), .C(n215), .Y(n5377) );
  OAI21X1 U12113 ( .A(n10836), .B(n10789), .C(n322), .Y(n5378) );
  OAI21X1 U12114 ( .A(n10838), .B(n10789), .C(n429), .Y(n5379) );
  OAI21X1 U12115 ( .A(n10840), .B(n10789), .C(n536), .Y(n5380) );
  OAI21X1 U12116 ( .A(n10842), .B(n10789), .C(n1620), .Y(n5381) );
  OAI21X1 U12117 ( .A(n10844), .B(n10789), .C(n1779), .Y(n5382) );
  OAI21X1 U12118 ( .A(n10846), .B(n10789), .C(n1937), .Y(n5383) );
  OAI21X1 U12119 ( .A(n10848), .B(n10789), .C(n2094), .Y(n5384) );
  OAI21X1 U12120 ( .A(n10850), .B(n10789), .C(n643), .Y(n5385) );
  OAI21X1 U12121 ( .A(n10852), .B(n10789), .C(n755), .Y(n5386) );
  OAI21X1 U12122 ( .A(n10854), .B(n10789), .C(n867), .Y(n5387) );
  OAI21X1 U12123 ( .A(n10856), .B(n10789), .C(n979), .Y(n5388) );
  OAI21X1 U12124 ( .A(n10858), .B(n10789), .C(n214), .Y(n5389) );
  OAI21X1 U12125 ( .A(n10860), .B(n10789), .C(n321), .Y(n5390) );
  OAI21X1 U12126 ( .A(n10862), .B(n10789), .C(n428), .Y(n5391) );
  OAI21X1 U12127 ( .A(n10864), .B(n10789), .C(n535), .Y(n5392) );
  OAI21X1 U12128 ( .A(n10866), .B(n10789), .C(n1619), .Y(n5393) );
  OAI21X1 U12129 ( .A(n10868), .B(n10789), .C(n1778), .Y(n5394) );
  OAI21X1 U12130 ( .A(n10870), .B(n10789), .C(n1936), .Y(n5395) );
  OAI21X1 U12131 ( .A(n10872), .B(n10789), .C(n2093), .Y(n5396) );
  OAI21X1 U12132 ( .A(n10874), .B(n10789), .C(n1102), .Y(n5397) );
  OAI21X1 U12133 ( .A(n10876), .B(n10789), .C(n642), .Y(n5398) );
  OAI21X1 U12134 ( .A(n10878), .B(n10789), .C(n754), .Y(n5399) );
  OAI21X1 U12135 ( .A(n10880), .B(n10789), .C(n866), .Y(n5400) );
  OAI21X1 U12136 ( .A(n10882), .B(n10789), .C(n978), .Y(n5401) );
  OAI21X1 U12137 ( .A(n10884), .B(n10789), .C(n213), .Y(n5402) );
  OAI21X1 U12138 ( .A(n10886), .B(n10789), .C(n320), .Y(n5403) );
  OAI21X1 U12139 ( .A(n10888), .B(n10789), .C(n427), .Y(n5404) );
  OAI21X1 U12140 ( .A(n10890), .B(n10789), .C(n534), .Y(n5405) );
  OAI21X1 U12141 ( .A(n10892), .B(n10789), .C(n1618), .Y(n5406) );
  OAI21X1 U12142 ( .A(n10894), .B(n10789), .C(n1777), .Y(n5407) );
  OAI21X1 U12143 ( .A(n10896), .B(n10789), .C(n1935), .Y(n5408) );
  OAI21X1 U12144 ( .A(n10898), .B(n10789), .C(n2092), .Y(n5409) );
  OAI21X1 U12145 ( .A(n10900), .B(n10789), .C(n1101), .Y(n5410) );
  OAI21X1 U12146 ( .A(n10902), .B(n10789), .C(n641), .Y(n5411) );
  OAI21X1 U12147 ( .A(n10904), .B(n10789), .C(n753), .Y(n5412) );
  OAI21X1 U12148 ( .A(n10906), .B(n10789), .C(n865), .Y(n5413) );
  OAI21X1 U12149 ( .A(n10908), .B(n10789), .C(n977), .Y(n5414) );
  OAI21X1 U12150 ( .A(n10910), .B(n10789), .C(n212), .Y(n5415) );
  OAI21X1 U12151 ( .A(n10912), .B(n10789), .C(n319), .Y(n5416) );
  OAI21X1 U12152 ( .A(n10914), .B(n10789), .C(n426), .Y(n5417) );
  OAI21X1 U12153 ( .A(n10916), .B(n10789), .C(n533), .Y(n5418) );
  OAI21X1 U12154 ( .A(n10918), .B(n10789), .C(n1617), .Y(n5419) );
  OAI21X1 U12155 ( .A(n10920), .B(n10789), .C(n1776), .Y(n5420) );
  OAI21X1 U12156 ( .A(n10922), .B(n10789), .C(n1934), .Y(n5421) );
  OAI21X1 U12157 ( .A(n10924), .B(n10789), .C(n2091), .Y(n5422) );
  OAI21X1 U12158 ( .A(n10926), .B(n10789), .C(n1100), .Y(n5423) );
  OAI21X1 U12159 ( .A(n10928), .B(n10789), .C(n640), .Y(n5424) );
  OAI21X1 U12160 ( .A(n10930), .B(n10789), .C(n752), .Y(n5425) );
  OAI21X1 U12161 ( .A(n10932), .B(n10789), .C(n864), .Y(n5426) );
  OAI21X1 U12162 ( .A(n10934), .B(n10789), .C(n976), .Y(n5427) );
  OAI21X1 U12163 ( .A(n10936), .B(n10789), .C(n211), .Y(n5428) );
  OAI21X1 U12164 ( .A(n10938), .B(n10789), .C(n318), .Y(n5429) );
  OAI21X1 U12165 ( .A(n10940), .B(n10789), .C(n425), .Y(n5430) );
  OAI21X1 U12166 ( .A(n10942), .B(n10789), .C(n532), .Y(n5431) );
  OAI21X1 U12167 ( .A(n10944), .B(n10789), .C(n1616), .Y(n5432) );
  OAI21X1 U12168 ( .A(n10946), .B(n10789), .C(n1775), .Y(n5433) );
  OAI21X1 U12169 ( .A(n10948), .B(n10789), .C(n1933), .Y(n5434) );
  OAI21X1 U12170 ( .A(n10950), .B(n10789), .C(n2090), .Y(n5435) );
  OAI21X1 U12171 ( .A(n10954), .B(n10789), .C(n1099), .Y(n5436) );
  OAI21X1 U12172 ( .A(n1143), .B(n1994), .C(n10956), .Y(n11906) );
  OAI21X1 U12173 ( .A(n10826), .B(n10791), .C(n2089), .Y(n5437) );
  OAI21X1 U12174 ( .A(n10828), .B(n10791), .C(n1932), .Y(n5438) );
  OAI21X1 U12175 ( .A(n10830), .B(n10791), .C(n1774), .Y(n5439) );
  OAI21X1 U12176 ( .A(n10832), .B(n10791), .C(n1615), .Y(n5440) );
  OAI21X1 U12177 ( .A(n10834), .B(n10791), .C(n1474), .Y(n5441) );
  OAI21X1 U12178 ( .A(n10836), .B(n10791), .C(n1348), .Y(n5442) );
  OAI21X1 U12179 ( .A(n10838), .B(n10791), .C(n1223), .Y(n5443) );
  OAI21X1 U12180 ( .A(n10840), .B(n10791), .C(n1098), .Y(n5444) );
  OAI21X1 U12181 ( .A(n10842), .B(n10791), .C(n975), .Y(n5445) );
  OAI21X1 U12182 ( .A(n10844), .B(n10791), .C(n863), .Y(n5446) );
  OAI21X1 U12183 ( .A(n10846), .B(n10791), .C(n751), .Y(n5447) );
  OAI21X1 U12184 ( .A(n10848), .B(n10791), .C(n639), .Y(n5448) );
  OAI21X1 U12185 ( .A(n10850), .B(n10791), .C(n2088), .Y(n5449) );
  OAI21X1 U12186 ( .A(n10852), .B(n10791), .C(n1931), .Y(n5450) );
  OAI21X1 U12187 ( .A(n10854), .B(n10791), .C(n1773), .Y(n5451) );
  OAI21X1 U12188 ( .A(n10856), .B(n10791), .C(n1614), .Y(n5452) );
  OAI21X1 U12189 ( .A(n10858), .B(n10791), .C(n1473), .Y(n5453) );
  OAI21X1 U12190 ( .A(n10860), .B(n10791), .C(n1347), .Y(n5454) );
  OAI21X1 U12191 ( .A(n10862), .B(n10791), .C(n1222), .Y(n5455) );
  OAI21X1 U12192 ( .A(n10864), .B(n10791), .C(n1097), .Y(n5456) );
  OAI21X1 U12193 ( .A(n10866), .B(n10791), .C(n974), .Y(n5457) );
  OAI21X1 U12194 ( .A(n10868), .B(n10791), .C(n862), .Y(n5458) );
  OAI21X1 U12195 ( .A(n10870), .B(n10791), .C(n750), .Y(n5459) );
  OAI21X1 U12196 ( .A(n10872), .B(n10791), .C(n638), .Y(n5460) );
  OAI21X1 U12197 ( .A(n10874), .B(n10791), .C(n531), .Y(n5461) );
  OAI21X1 U12198 ( .A(n10876), .B(n10791), .C(n2087), .Y(n5462) );
  OAI21X1 U12199 ( .A(n10878), .B(n10791), .C(n1930), .Y(n5463) );
  OAI21X1 U12200 ( .A(n10880), .B(n10791), .C(n1772), .Y(n5464) );
  OAI21X1 U12201 ( .A(n10882), .B(n10791), .C(n1613), .Y(n5465) );
  OAI21X1 U12202 ( .A(n10884), .B(n10791), .C(n1472), .Y(n5466) );
  OAI21X1 U12203 ( .A(n10886), .B(n10791), .C(n1346), .Y(n5467) );
  OAI21X1 U12204 ( .A(n10888), .B(n10791), .C(n1221), .Y(n5468) );
  OAI21X1 U12205 ( .A(n10890), .B(n10791), .C(n1096), .Y(n5469) );
  OAI21X1 U12206 ( .A(n10892), .B(n10791), .C(n973), .Y(n5470) );
  OAI21X1 U12207 ( .A(n10894), .B(n10791), .C(n861), .Y(n5471) );
  OAI21X1 U12208 ( .A(n10896), .B(n10791), .C(n749), .Y(n5472) );
  OAI21X1 U12209 ( .A(n10898), .B(n10791), .C(n637), .Y(n5473) );
  OAI21X1 U12210 ( .A(n10900), .B(n10791), .C(n530), .Y(n5474) );
  OAI21X1 U12211 ( .A(n10902), .B(n10791), .C(n2086), .Y(n5475) );
  OAI21X1 U12212 ( .A(n10904), .B(n10791), .C(n1929), .Y(n5476) );
  OAI21X1 U12213 ( .A(n10906), .B(n10791), .C(n1771), .Y(n5477) );
  OAI21X1 U12214 ( .A(n10908), .B(n10791), .C(n1612), .Y(n5478) );
  OAI21X1 U12215 ( .A(n10910), .B(n10791), .C(n1471), .Y(n5479) );
  OAI21X1 U12216 ( .A(n10912), .B(n10791), .C(n1345), .Y(n5480) );
  OAI21X1 U12217 ( .A(n10914), .B(n10791), .C(n1220), .Y(n5481) );
  OAI21X1 U12218 ( .A(n10916), .B(n10791), .C(n1095), .Y(n5482) );
  OAI21X1 U12219 ( .A(n10918), .B(n10791), .C(n972), .Y(n5483) );
  OAI21X1 U12220 ( .A(n10920), .B(n10791), .C(n860), .Y(n5484) );
  OAI21X1 U12221 ( .A(n10922), .B(n10791), .C(n748), .Y(n5485) );
  OAI21X1 U12222 ( .A(n10924), .B(n10791), .C(n636), .Y(n5486) );
  OAI21X1 U12223 ( .A(n10926), .B(n10791), .C(n529), .Y(n5487) );
  OAI21X1 U12224 ( .A(n10928), .B(n10791), .C(n2085), .Y(n5488) );
  OAI21X1 U12225 ( .A(n10930), .B(n10791), .C(n1928), .Y(n5489) );
  OAI21X1 U12226 ( .A(n10932), .B(n10791), .C(n1770), .Y(n5490) );
  OAI21X1 U12227 ( .A(n10934), .B(n10791), .C(n1611), .Y(n5491) );
  OAI21X1 U12228 ( .A(n10936), .B(n10791), .C(n1470), .Y(n5492) );
  OAI21X1 U12229 ( .A(n10938), .B(n10791), .C(n1344), .Y(n5493) );
  OAI21X1 U12230 ( .A(n10940), .B(n10791), .C(n1219), .Y(n5494) );
  OAI21X1 U12231 ( .A(n10942), .B(n10791), .C(n1094), .Y(n5495) );
  OAI21X1 U12232 ( .A(n10944), .B(n10791), .C(n971), .Y(n5496) );
  OAI21X1 U12233 ( .A(n10946), .B(n10791), .C(n859), .Y(n5497) );
  OAI21X1 U12234 ( .A(n10948), .B(n10791), .C(n747), .Y(n5498) );
  OAI21X1 U12235 ( .A(n10950), .B(n10791), .C(n635), .Y(n5499) );
  OAI21X1 U12236 ( .A(n10954), .B(n10791), .C(n528), .Y(n5500) );
  OAI21X1 U12237 ( .A(n1268), .B(n1994), .C(n10956), .Y(n11972) );
  OAI21X1 U12238 ( .A(n10826), .B(n10793), .C(n1927), .Y(n5501) );
  OAI21X1 U12239 ( .A(n10828), .B(n10793), .C(n2084), .Y(n5502) );
  OAI21X1 U12240 ( .A(n10830), .B(n10793), .C(n1610), .Y(n5503) );
  OAI21X1 U12241 ( .A(n10832), .B(n10793), .C(n1769), .Y(n5504) );
  OAI21X1 U12242 ( .A(n10834), .B(n10793), .C(n1343), .Y(n5505) );
  OAI21X1 U12243 ( .A(n10836), .B(n10793), .C(n1469), .Y(n5506) );
  OAI21X1 U12244 ( .A(n10838), .B(n10793), .C(n1093), .Y(n5507) );
  OAI21X1 U12245 ( .A(n10840), .B(n10793), .C(n1218), .Y(n5508) );
  OAI21X1 U12246 ( .A(n10842), .B(n10793), .C(n858), .Y(n5509) );
  OAI21X1 U12247 ( .A(n10844), .B(n10793), .C(n970), .Y(n5510) );
  OAI21X1 U12248 ( .A(n10846), .B(n10793), .C(n634), .Y(n5511) );
  OAI21X1 U12249 ( .A(n10848), .B(n10793), .C(n746), .Y(n5512) );
  OAI21X1 U12250 ( .A(n10850), .B(n10793), .C(n1926), .Y(n5513) );
  OAI21X1 U12251 ( .A(n10852), .B(n10793), .C(n2083), .Y(n5514) );
  OAI21X1 U12252 ( .A(n10854), .B(n10793), .C(n1609), .Y(n5515) );
  OAI21X1 U12253 ( .A(n10856), .B(n10793), .C(n1768), .Y(n5516) );
  OAI21X1 U12254 ( .A(n10858), .B(n10793), .C(n1342), .Y(n5517) );
  OAI21X1 U12255 ( .A(n10860), .B(n10793), .C(n1468), .Y(n5518) );
  OAI21X1 U12256 ( .A(n10862), .B(n10793), .C(n1092), .Y(n5519) );
  OAI21X1 U12257 ( .A(n10864), .B(n10793), .C(n1217), .Y(n5520) );
  OAI21X1 U12258 ( .A(n10866), .B(n10793), .C(n857), .Y(n5521) );
  OAI21X1 U12259 ( .A(n10868), .B(n10793), .C(n969), .Y(n5522) );
  OAI21X1 U12260 ( .A(n10870), .B(n10793), .C(n633), .Y(n5523) );
  OAI21X1 U12261 ( .A(n10872), .B(n10793), .C(n745), .Y(n5524) );
  OAI21X1 U12262 ( .A(n10874), .B(n10793), .C(n424), .Y(n5525) );
  OAI21X1 U12263 ( .A(n10876), .B(n10793), .C(n1925), .Y(n5526) );
  OAI21X1 U12264 ( .A(n10878), .B(n10793), .C(n2082), .Y(n5527) );
  OAI21X1 U12265 ( .A(n10880), .B(n10793), .C(n1608), .Y(n5528) );
  OAI21X1 U12266 ( .A(n10882), .B(n10793), .C(n1767), .Y(n5529) );
  OAI21X1 U12267 ( .A(n10884), .B(n10793), .C(n1341), .Y(n5530) );
  OAI21X1 U12268 ( .A(n10886), .B(n10793), .C(n1467), .Y(n5531) );
  OAI21X1 U12269 ( .A(n10888), .B(n10793), .C(n1091), .Y(n5532) );
  OAI21X1 U12270 ( .A(n10890), .B(n10793), .C(n1216), .Y(n5533) );
  OAI21X1 U12271 ( .A(n10892), .B(n10793), .C(n856), .Y(n5534) );
  OAI21X1 U12272 ( .A(n10894), .B(n10793), .C(n968), .Y(n5535) );
  OAI21X1 U12273 ( .A(n10896), .B(n10793), .C(n632), .Y(n5536) );
  OAI21X1 U12274 ( .A(n10898), .B(n10793), .C(n744), .Y(n5537) );
  OAI21X1 U12275 ( .A(n10900), .B(n10793), .C(n423), .Y(n5538) );
  OAI21X1 U12276 ( .A(n10902), .B(n10793), .C(n1924), .Y(n5539) );
  OAI21X1 U12277 ( .A(n10904), .B(n10793), .C(n2081), .Y(n5540) );
  OAI21X1 U12278 ( .A(n10906), .B(n10793), .C(n1607), .Y(n5541) );
  OAI21X1 U12279 ( .A(n10908), .B(n10793), .C(n1766), .Y(n5542) );
  OAI21X1 U12280 ( .A(n10910), .B(n10793), .C(n1340), .Y(n5543) );
  OAI21X1 U12281 ( .A(n10912), .B(n10793), .C(n1466), .Y(n5544) );
  OAI21X1 U12282 ( .A(n10914), .B(n10793), .C(n1090), .Y(n5545) );
  OAI21X1 U12283 ( .A(n10916), .B(n10793), .C(n1215), .Y(n5546) );
  OAI21X1 U12284 ( .A(n10918), .B(n10793), .C(n855), .Y(n5547) );
  OAI21X1 U12285 ( .A(n10920), .B(n10793), .C(n967), .Y(n5548) );
  OAI21X1 U12286 ( .A(n10922), .B(n10793), .C(n631), .Y(n5549) );
  OAI21X1 U12287 ( .A(n10924), .B(n10793), .C(n743), .Y(n5550) );
  OAI21X1 U12288 ( .A(n10926), .B(n10793), .C(n422), .Y(n5551) );
  OAI21X1 U12289 ( .A(n10928), .B(n10793), .C(n1923), .Y(n5552) );
  OAI21X1 U12290 ( .A(n10930), .B(n10793), .C(n2080), .Y(n5553) );
  OAI21X1 U12291 ( .A(n10932), .B(n10793), .C(n1606), .Y(n5554) );
  OAI21X1 U12292 ( .A(n10934), .B(n10793), .C(n1765), .Y(n5555) );
  OAI21X1 U12293 ( .A(n10936), .B(n10793), .C(n1339), .Y(n5556) );
  OAI21X1 U12294 ( .A(n10938), .B(n10793), .C(n1465), .Y(n5557) );
  OAI21X1 U12295 ( .A(n10940), .B(n10793), .C(n1089), .Y(n5558) );
  OAI21X1 U12296 ( .A(n10942), .B(n10793), .C(n1214), .Y(n5559) );
  OAI21X1 U12297 ( .A(n10944), .B(n10793), .C(n854), .Y(n5560) );
  OAI21X1 U12298 ( .A(n10946), .B(n10793), .C(n966), .Y(n5561) );
  OAI21X1 U12299 ( .A(n10948), .B(n10793), .C(n630), .Y(n5562) );
  OAI21X1 U12300 ( .A(n10950), .B(n10793), .C(n742), .Y(n5563) );
  OAI21X1 U12301 ( .A(n10954), .B(n10793), .C(n421), .Y(n5564) );
  OAI21X1 U12302 ( .A(n1394), .B(n1994), .C(n10956), .Y(n12038) );
  OAI21X1 U12303 ( .A(n10826), .B(n10795), .C(n1764), .Y(n5565) );
  OAI21X1 U12304 ( .A(n10828), .B(n10795), .C(n1605), .Y(n5566) );
  OAI21X1 U12305 ( .A(n10830), .B(n10795), .C(n2079), .Y(n5567) );
  OAI21X1 U12306 ( .A(n10832), .B(n10795), .C(n1922), .Y(n5568) );
  OAI21X1 U12307 ( .A(n10834), .B(n10795), .C(n1213), .Y(n5569) );
  OAI21X1 U12308 ( .A(n10836), .B(n10795), .C(n1088), .Y(n5570) );
  OAI21X1 U12309 ( .A(n10838), .B(n10795), .C(n1464), .Y(n5571) );
  OAI21X1 U12310 ( .A(n10840), .B(n10795), .C(n1338), .Y(n5572) );
  OAI21X1 U12311 ( .A(n10842), .B(n10795), .C(n741), .Y(n5573) );
  OAI21X1 U12312 ( .A(n10844), .B(n10795), .C(n629), .Y(n5574) );
  OAI21X1 U12313 ( .A(n10846), .B(n10795), .C(n965), .Y(n5575) );
  OAI21X1 U12314 ( .A(n10848), .B(n10795), .C(n853), .Y(n5576) );
  OAI21X1 U12315 ( .A(n10850), .B(n10795), .C(n1763), .Y(n5577) );
  OAI21X1 U12316 ( .A(n10852), .B(n10795), .C(n1604), .Y(n5578) );
  OAI21X1 U12317 ( .A(n10854), .B(n10795), .C(n2078), .Y(n5579) );
  OAI21X1 U12318 ( .A(n10856), .B(n10795), .C(n1921), .Y(n5580) );
  OAI21X1 U12319 ( .A(n10858), .B(n10795), .C(n1212), .Y(n5581) );
  OAI21X1 U12320 ( .A(n10860), .B(n10795), .C(n1087), .Y(n5582) );
  OAI21X1 U12321 ( .A(n10862), .B(n10795), .C(n1463), .Y(n5583) );
  OAI21X1 U12322 ( .A(n10864), .B(n10795), .C(n1337), .Y(n5584) );
  OAI21X1 U12323 ( .A(n10866), .B(n10795), .C(n740), .Y(n5585) );
  OAI21X1 U12324 ( .A(n10868), .B(n10795), .C(n628), .Y(n5586) );
  OAI21X1 U12325 ( .A(n10870), .B(n10795), .C(n964), .Y(n5587) );
  OAI21X1 U12326 ( .A(n10872), .B(n10795), .C(n852), .Y(n5588) );
  OAI21X1 U12327 ( .A(n10874), .B(n10795), .C(n317), .Y(n5589) );
  OAI21X1 U12328 ( .A(n10876), .B(n10795), .C(n1762), .Y(n5590) );
  OAI21X1 U12329 ( .A(n10878), .B(n10795), .C(n1603), .Y(n5591) );
  OAI21X1 U12330 ( .A(n10880), .B(n10795), .C(n2077), .Y(n5592) );
  OAI21X1 U12331 ( .A(n10882), .B(n10795), .C(n1920), .Y(n5593) );
  OAI21X1 U12332 ( .A(n10884), .B(n10795), .C(n1211), .Y(n5594) );
  OAI21X1 U12333 ( .A(n10886), .B(n10795), .C(n1086), .Y(n5595) );
  OAI21X1 U12334 ( .A(n10888), .B(n10795), .C(n1462), .Y(n5596) );
  OAI21X1 U12335 ( .A(n10890), .B(n10795), .C(n1336), .Y(n5597) );
  OAI21X1 U12336 ( .A(n10892), .B(n10795), .C(n739), .Y(n5598) );
  OAI21X1 U12337 ( .A(n10894), .B(n10795), .C(n627), .Y(n5599) );
  OAI21X1 U12338 ( .A(n10896), .B(n10795), .C(n963), .Y(n5600) );
  OAI21X1 U12339 ( .A(n10898), .B(n10795), .C(n851), .Y(n5601) );
  OAI21X1 U12340 ( .A(n10900), .B(n10795), .C(n316), .Y(n5602) );
  OAI21X1 U12341 ( .A(n10902), .B(n10795), .C(n1761), .Y(n5603) );
  OAI21X1 U12342 ( .A(n10904), .B(n10795), .C(n1602), .Y(n5604) );
  OAI21X1 U12343 ( .A(n10906), .B(n10795), .C(n2076), .Y(n5605) );
  OAI21X1 U12344 ( .A(n10908), .B(n10795), .C(n1919), .Y(n5606) );
  OAI21X1 U12345 ( .A(n10910), .B(n10795), .C(n1210), .Y(n5607) );
  OAI21X1 U12346 ( .A(n10912), .B(n10795), .C(n1085), .Y(n5608) );
  OAI21X1 U12347 ( .A(n10914), .B(n10795), .C(n1461), .Y(n5609) );
  OAI21X1 U12348 ( .A(n10916), .B(n10795), .C(n1335), .Y(n5610) );
  OAI21X1 U12349 ( .A(n10918), .B(n10795), .C(n738), .Y(n5611) );
  OAI21X1 U12350 ( .A(n10920), .B(n10795), .C(n626), .Y(n5612) );
  OAI21X1 U12351 ( .A(n10922), .B(n10795), .C(n962), .Y(n5613) );
  OAI21X1 U12352 ( .A(n10924), .B(n10795), .C(n850), .Y(n5614) );
  OAI21X1 U12353 ( .A(n10926), .B(n10795), .C(n315), .Y(n5615) );
  OAI21X1 U12354 ( .A(n10928), .B(n10795), .C(n1760), .Y(n5616) );
  OAI21X1 U12355 ( .A(n10930), .B(n10795), .C(n1601), .Y(n5617) );
  OAI21X1 U12356 ( .A(n10932), .B(n10795), .C(n2075), .Y(n5618) );
  OAI21X1 U12357 ( .A(n10934), .B(n10795), .C(n1918), .Y(n5619) );
  OAI21X1 U12358 ( .A(n10936), .B(n10795), .C(n1209), .Y(n5620) );
  OAI21X1 U12359 ( .A(n10938), .B(n10795), .C(n1084), .Y(n5621) );
  OAI21X1 U12360 ( .A(n10940), .B(n10795), .C(n1460), .Y(n5622) );
  OAI21X1 U12361 ( .A(n10942), .B(n10795), .C(n1334), .Y(n5623) );
  OAI21X1 U12362 ( .A(n10944), .B(n10795), .C(n737), .Y(n5624) );
  OAI21X1 U12363 ( .A(n10946), .B(n10795), .C(n625), .Y(n5625) );
  OAI21X1 U12364 ( .A(n10948), .B(n10795), .C(n961), .Y(n5626) );
  OAI21X1 U12365 ( .A(n10950), .B(n10795), .C(n849), .Y(n5627) );
  OAI21X1 U12366 ( .A(n10954), .B(n10795), .C(n314), .Y(n5628) );
  OAI21X1 U12367 ( .A(n1678), .B(n1994), .C(n10956), .Y(n12105) );
  OAI21X1 U12368 ( .A(n10826), .B(n10797), .C(n1600), .Y(n5629) );
  OAI21X1 U12369 ( .A(n10828), .B(n10797), .C(n1759), .Y(n5630) );
  OAI21X1 U12370 ( .A(n10830), .B(n10797), .C(n1917), .Y(n5631) );
  OAI21X1 U12371 ( .A(n10832), .B(n10797), .C(n2074), .Y(n5632) );
  OAI21X1 U12372 ( .A(n10834), .B(n10797), .C(n1083), .Y(n5633) );
  OAI21X1 U12373 ( .A(n10836), .B(n10797), .C(n1208), .Y(n5634) );
  OAI21X1 U12374 ( .A(n10838), .B(n10797), .C(n1333), .Y(n5635) );
  OAI21X1 U12375 ( .A(n10840), .B(n10797), .C(n1459), .Y(n5636) );
  OAI21X1 U12376 ( .A(n10842), .B(n10797), .C(n624), .Y(n5637) );
  OAI21X1 U12377 ( .A(n10844), .B(n10797), .C(n736), .Y(n5638) );
  OAI21X1 U12378 ( .A(n10846), .B(n10797), .C(n848), .Y(n5639) );
  OAI21X1 U12379 ( .A(n10848), .B(n10797), .C(n960), .Y(n5640) );
  OAI21X1 U12380 ( .A(n10850), .B(n10797), .C(n1599), .Y(n5641) );
  OAI21X1 U12381 ( .A(n10852), .B(n10797), .C(n1758), .Y(n5642) );
  OAI21X1 U12382 ( .A(n10854), .B(n10797), .C(n1916), .Y(n5643) );
  OAI21X1 U12383 ( .A(n10856), .B(n10797), .C(n2073), .Y(n5644) );
  OAI21X1 U12384 ( .A(n10858), .B(n10797), .C(n1082), .Y(n5645) );
  OAI21X1 U12385 ( .A(n10860), .B(n10797), .C(n1207), .Y(n5646) );
  OAI21X1 U12386 ( .A(n10862), .B(n10797), .C(n1332), .Y(n5647) );
  OAI21X1 U12387 ( .A(n10864), .B(n10797), .C(n1458), .Y(n5648) );
  OAI21X1 U12388 ( .A(n10866), .B(n10797), .C(n623), .Y(n5649) );
  OAI21X1 U12389 ( .A(n10868), .B(n10797), .C(n735), .Y(n5650) );
  OAI21X1 U12390 ( .A(n10870), .B(n10797), .C(n847), .Y(n5651) );
  OAI21X1 U12391 ( .A(n10872), .B(n10797), .C(n959), .Y(n5652) );
  OAI21X1 U12392 ( .A(n10874), .B(n10797), .C(n210), .Y(n5653) );
  OAI21X1 U12393 ( .A(n10876), .B(n10797), .C(n1598), .Y(n5654) );
  OAI21X1 U12394 ( .A(n10878), .B(n10797), .C(n1757), .Y(n5655) );
  OAI21X1 U12395 ( .A(n10880), .B(n10797), .C(n1915), .Y(n5656) );
  OAI21X1 U12396 ( .A(n10882), .B(n10797), .C(n2072), .Y(n5657) );
  OAI21X1 U12397 ( .A(n10884), .B(n10797), .C(n1081), .Y(n5658) );
  OAI21X1 U12398 ( .A(n10886), .B(n10797), .C(n1206), .Y(n5659) );
  OAI21X1 U12399 ( .A(n10888), .B(n10797), .C(n1331), .Y(n5660) );
  OAI21X1 U12400 ( .A(n10890), .B(n10797), .C(n1457), .Y(n5661) );
  OAI21X1 U12401 ( .A(n10892), .B(n10797), .C(n622), .Y(n5662) );
  OAI21X1 U12402 ( .A(n10894), .B(n10797), .C(n734), .Y(n5663) );
  OAI21X1 U12403 ( .A(n10896), .B(n10797), .C(n846), .Y(n5664) );
  OAI21X1 U12404 ( .A(n10898), .B(n10797), .C(n958), .Y(n5665) );
  OAI21X1 U12405 ( .A(n10900), .B(n10797), .C(n209), .Y(n5666) );
  OAI21X1 U12406 ( .A(n10902), .B(n10797), .C(n1597), .Y(n5667) );
  OAI21X1 U12407 ( .A(n10904), .B(n10797), .C(n1756), .Y(n5668) );
  OAI21X1 U12408 ( .A(n10906), .B(n10797), .C(n1914), .Y(n5669) );
  OAI21X1 U12409 ( .A(n10908), .B(n10797), .C(n2071), .Y(n5670) );
  OAI21X1 U12410 ( .A(n10910), .B(n10797), .C(n1080), .Y(n5671) );
  OAI21X1 U12411 ( .A(n10912), .B(n10797), .C(n1205), .Y(n5672) );
  OAI21X1 U12412 ( .A(n10914), .B(n10797), .C(n1330), .Y(n5673) );
  OAI21X1 U12413 ( .A(n10916), .B(n10797), .C(n1456), .Y(n5674) );
  OAI21X1 U12414 ( .A(n10918), .B(n10797), .C(n621), .Y(n5675) );
  OAI21X1 U12415 ( .A(n10920), .B(n10797), .C(n733), .Y(n5676) );
  OAI21X1 U12416 ( .A(n10922), .B(n10797), .C(n845), .Y(n5677) );
  OAI21X1 U12417 ( .A(n10924), .B(n10797), .C(n957), .Y(n5678) );
  OAI21X1 U12418 ( .A(n10926), .B(n10797), .C(n208), .Y(n5679) );
  OAI21X1 U12419 ( .A(n10928), .B(n10797), .C(n1596), .Y(n5680) );
  OAI21X1 U12420 ( .A(n10930), .B(n10797), .C(n1755), .Y(n5681) );
  OAI21X1 U12421 ( .A(n10932), .B(n10797), .C(n1913), .Y(n5682) );
  OAI21X1 U12422 ( .A(n10934), .B(n10797), .C(n2070), .Y(n5683) );
  OAI21X1 U12423 ( .A(n10936), .B(n10797), .C(n1079), .Y(n5684) );
  OAI21X1 U12424 ( .A(n10938), .B(n10797), .C(n1204), .Y(n5685) );
  OAI21X1 U12425 ( .A(n10940), .B(n10797), .C(n1329), .Y(n5686) );
  OAI21X1 U12426 ( .A(n10942), .B(n10797), .C(n1455), .Y(n5687) );
  OAI21X1 U12427 ( .A(n10944), .B(n10797), .C(n620), .Y(n5688) );
  OAI21X1 U12428 ( .A(n10946), .B(n10797), .C(n732), .Y(n5689) );
  OAI21X1 U12429 ( .A(n10948), .B(n10797), .C(n844), .Y(n5690) );
  OAI21X1 U12430 ( .A(n10950), .B(n10797), .C(n956), .Y(n5691) );
  OAI21X1 U12431 ( .A(n10954), .B(n10797), .C(n207), .Y(n5692) );
  NAND3X1 U12432 ( .A(n10963), .B(n10965), .C(n11112), .Y(n12633) );
  OAI21X1 U12433 ( .A(n1520), .B(n1837), .C(n10956), .Y(n12171) );
  OAI21X1 U12434 ( .A(n10826), .B(n10799), .C(n1454), .Y(n5693) );
  OAI21X1 U12435 ( .A(n10828), .B(n10799), .C(n1328), .Y(n5694) );
  OAI21X1 U12436 ( .A(n10830), .B(n10799), .C(n1203), .Y(n5695) );
  OAI21X1 U12437 ( .A(n10832), .B(n10799), .C(n1078), .Y(n5696) );
  OAI21X1 U12438 ( .A(n10834), .B(n10799), .C(n2069), .Y(n5697) );
  OAI21X1 U12439 ( .A(n10836), .B(n10799), .C(n1912), .Y(n5698) );
  OAI21X1 U12440 ( .A(n10838), .B(n10799), .C(n1754), .Y(n5699) );
  OAI21X1 U12441 ( .A(n10840), .B(n10799), .C(n1595), .Y(n5700) );
  OAI21X1 U12442 ( .A(n10842), .B(n10799), .C(n527), .Y(n5701) );
  OAI21X1 U12443 ( .A(n10844), .B(n10799), .C(n420), .Y(n5702) );
  OAI21X1 U12444 ( .A(n10846), .B(n10799), .C(n313), .Y(n5703) );
  OAI21X1 U12445 ( .A(n10848), .B(n10799), .C(n206), .Y(n5704) );
  OAI21X1 U12446 ( .A(n10850), .B(n10799), .C(n1453), .Y(n5705) );
  OAI21X1 U12447 ( .A(n10852), .B(n10799), .C(n1327), .Y(n5706) );
  OAI21X1 U12448 ( .A(n10854), .B(n10799), .C(n1202), .Y(n5707) );
  OAI21X1 U12449 ( .A(n10856), .B(n10799), .C(n1077), .Y(n5708) );
  OAI21X1 U12450 ( .A(n10858), .B(n10799), .C(n2068), .Y(n5709) );
  OAI21X1 U12451 ( .A(n10860), .B(n10799), .C(n1911), .Y(n5710) );
  OAI21X1 U12452 ( .A(n10862), .B(n10799), .C(n1753), .Y(n5711) );
  OAI21X1 U12453 ( .A(n10864), .B(n10799), .C(n1594), .Y(n5712) );
  OAI21X1 U12454 ( .A(n10866), .B(n10799), .C(n526), .Y(n5713) );
  OAI21X1 U12455 ( .A(n10868), .B(n10799), .C(n419), .Y(n5714) );
  OAI21X1 U12456 ( .A(n10870), .B(n10799), .C(n312), .Y(n5715) );
  OAI21X1 U12457 ( .A(n10872), .B(n10799), .C(n205), .Y(n5716) );
  OAI21X1 U12458 ( .A(n10874), .B(n10799), .C(n955), .Y(n5717) );
  OAI21X1 U12459 ( .A(n10876), .B(n10799), .C(n1452), .Y(n5718) );
  OAI21X1 U12460 ( .A(n10878), .B(n10799), .C(n1326), .Y(n5719) );
  OAI21X1 U12461 ( .A(n10880), .B(n10799), .C(n1201), .Y(n5720) );
  OAI21X1 U12462 ( .A(n10882), .B(n10799), .C(n1076), .Y(n5721) );
  OAI21X1 U12463 ( .A(n10884), .B(n10799), .C(n2067), .Y(n5722) );
  OAI21X1 U12464 ( .A(n10886), .B(n10799), .C(n1910), .Y(n5723) );
  OAI21X1 U12465 ( .A(n10888), .B(n10799), .C(n1752), .Y(n5724) );
  OAI21X1 U12466 ( .A(n10890), .B(n10799), .C(n1593), .Y(n5725) );
  OAI21X1 U12467 ( .A(n10892), .B(n10799), .C(n525), .Y(n5726) );
  OAI21X1 U12468 ( .A(n10894), .B(n10799), .C(n418), .Y(n5727) );
  OAI21X1 U12469 ( .A(n10896), .B(n10799), .C(n311), .Y(n5728) );
  OAI21X1 U12470 ( .A(n10898), .B(n10799), .C(n204), .Y(n5729) );
  OAI21X1 U12471 ( .A(n10900), .B(n10799), .C(n954), .Y(n5730) );
  OAI21X1 U12472 ( .A(n10902), .B(n10799), .C(n1451), .Y(n5731) );
  OAI21X1 U12473 ( .A(n10904), .B(n10799), .C(n1325), .Y(n5732) );
  OAI21X1 U12474 ( .A(n10906), .B(n10799), .C(n1200), .Y(n5733) );
  OAI21X1 U12475 ( .A(n10908), .B(n10799), .C(n1075), .Y(n5734) );
  OAI21X1 U12476 ( .A(n10910), .B(n10799), .C(n2066), .Y(n5735) );
  OAI21X1 U12477 ( .A(n10912), .B(n10799), .C(n1909), .Y(n5736) );
  OAI21X1 U12478 ( .A(n10914), .B(n10799), .C(n1751), .Y(n5737) );
  OAI21X1 U12479 ( .A(n10916), .B(n10799), .C(n1592), .Y(n5738) );
  OAI21X1 U12480 ( .A(n10918), .B(n10799), .C(n524), .Y(n5739) );
  OAI21X1 U12481 ( .A(n10920), .B(n10799), .C(n417), .Y(n5740) );
  OAI21X1 U12482 ( .A(n10922), .B(n10799), .C(n310), .Y(n5741) );
  OAI21X1 U12483 ( .A(n10924), .B(n10799), .C(n203), .Y(n5742) );
  OAI21X1 U12484 ( .A(n10926), .B(n10799), .C(n953), .Y(n5743) );
  OAI21X1 U12485 ( .A(n10928), .B(n10799), .C(n1450), .Y(n5744) );
  OAI21X1 U12486 ( .A(n10930), .B(n10799), .C(n1324), .Y(n5745) );
  OAI21X1 U12487 ( .A(n10932), .B(n10799), .C(n1199), .Y(n5746) );
  OAI21X1 U12488 ( .A(n10934), .B(n10799), .C(n1074), .Y(n5747) );
  OAI21X1 U12489 ( .A(n10936), .B(n10799), .C(n2065), .Y(n5748) );
  OAI21X1 U12490 ( .A(n10938), .B(n10799), .C(n1908), .Y(n5749) );
  OAI21X1 U12491 ( .A(n10940), .B(n10799), .C(n1750), .Y(n5750) );
  OAI21X1 U12492 ( .A(n10942), .B(n10799), .C(n1591), .Y(n5751) );
  OAI21X1 U12493 ( .A(n10944), .B(n10799), .C(n523), .Y(n5752) );
  OAI21X1 U12494 ( .A(n10946), .B(n10799), .C(n416), .Y(n5753) );
  OAI21X1 U12495 ( .A(n10948), .B(n10799), .C(n309), .Y(n5754) );
  OAI21X1 U12496 ( .A(n10950), .B(n10799), .C(n202), .Y(n5755) );
  OAI21X1 U12497 ( .A(n10954), .B(n10799), .C(n952), .Y(n5756) );
  OAI21X1 U12498 ( .A(n1395), .B(n1837), .C(n10956), .Y(n12237) );
  OAI21X1 U12499 ( .A(n10826), .B(n10801), .C(n1323), .Y(n5757) );
  OAI21X1 U12500 ( .A(n10828), .B(n10801), .C(n1449), .Y(n5758) );
  OAI21X1 U12501 ( .A(n10830), .B(n10801), .C(n1073), .Y(n5759) );
  OAI21X1 U12502 ( .A(n10832), .B(n10801), .C(n1198), .Y(n5760) );
  OAI21X1 U12503 ( .A(n10834), .B(n10801), .C(n1907), .Y(n5761) );
  OAI21X1 U12504 ( .A(n10836), .B(n10801), .C(n2064), .Y(n5762) );
  OAI21X1 U12505 ( .A(n10838), .B(n10801), .C(n1590), .Y(n5763) );
  OAI21X1 U12506 ( .A(n10840), .B(n10801), .C(n1749), .Y(n5764) );
  OAI21X1 U12507 ( .A(n10842), .B(n10801), .C(n415), .Y(n5765) );
  OAI21X1 U12508 ( .A(n10844), .B(n10801), .C(n522), .Y(n5766) );
  OAI21X1 U12509 ( .A(n10846), .B(n10801), .C(n201), .Y(n5767) );
  OAI21X1 U12510 ( .A(n10848), .B(n10801), .C(n308), .Y(n5768) );
  OAI21X1 U12511 ( .A(n10850), .B(n10801), .C(n1322), .Y(n5769) );
  OAI21X1 U12512 ( .A(n10852), .B(n10801), .C(n1448), .Y(n5770) );
  OAI21X1 U12513 ( .A(n10854), .B(n10801), .C(n1072), .Y(n5771) );
  OAI21X1 U12514 ( .A(n10856), .B(n10801), .C(n1197), .Y(n5772) );
  OAI21X1 U12515 ( .A(n10858), .B(n10801), .C(n1906), .Y(n5773) );
  OAI21X1 U12516 ( .A(n10860), .B(n10801), .C(n2063), .Y(n5774) );
  OAI21X1 U12517 ( .A(n10862), .B(n10801), .C(n1589), .Y(n5775) );
  OAI21X1 U12518 ( .A(n10864), .B(n10801), .C(n1748), .Y(n5776) );
  OAI21X1 U12519 ( .A(n10866), .B(n10801), .C(n414), .Y(n5777) );
  OAI21X1 U12520 ( .A(n10868), .B(n10801), .C(n521), .Y(n5778) );
  OAI21X1 U12521 ( .A(n10870), .B(n10801), .C(n200), .Y(n5779) );
  OAI21X1 U12522 ( .A(n10872), .B(n10801), .C(n307), .Y(n5780) );
  OAI21X1 U12523 ( .A(n10874), .B(n10801), .C(n843), .Y(n5781) );
  OAI21X1 U12524 ( .A(n10876), .B(n10801), .C(n1321), .Y(n5782) );
  OAI21X1 U12525 ( .A(n10878), .B(n10801), .C(n1447), .Y(n5783) );
  OAI21X1 U12526 ( .A(n10880), .B(n10801), .C(n1071), .Y(n5784) );
  OAI21X1 U12527 ( .A(n10882), .B(n10801), .C(n1196), .Y(n5785) );
  OAI21X1 U12528 ( .A(n10884), .B(n10801), .C(n1905), .Y(n5786) );
  OAI21X1 U12529 ( .A(n10886), .B(n10801), .C(n2062), .Y(n5787) );
  OAI21X1 U12530 ( .A(n10888), .B(n10801), .C(n1588), .Y(n5788) );
  OAI21X1 U12531 ( .A(n10890), .B(n10801), .C(n1747), .Y(n5789) );
  OAI21X1 U12532 ( .A(n10892), .B(n10801), .C(n413), .Y(n5790) );
  OAI21X1 U12533 ( .A(n10894), .B(n10801), .C(n520), .Y(n5791) );
  OAI21X1 U12534 ( .A(n10896), .B(n10801), .C(n199), .Y(n5792) );
  OAI21X1 U12535 ( .A(n10898), .B(n10801), .C(n306), .Y(n5793) );
  OAI21X1 U12536 ( .A(n10900), .B(n10801), .C(n842), .Y(n5794) );
  OAI21X1 U12537 ( .A(n10902), .B(n10801), .C(n1320), .Y(n5795) );
  OAI21X1 U12538 ( .A(n10904), .B(n10801), .C(n1446), .Y(n5796) );
  OAI21X1 U12539 ( .A(n10906), .B(n10801), .C(n1070), .Y(n5797) );
  OAI21X1 U12540 ( .A(n10908), .B(n10801), .C(n1195), .Y(n5798) );
  OAI21X1 U12541 ( .A(n10910), .B(n10801), .C(n1904), .Y(n5799) );
  OAI21X1 U12542 ( .A(n10912), .B(n10801), .C(n2061), .Y(n5800) );
  OAI21X1 U12543 ( .A(n10914), .B(n10801), .C(n1587), .Y(n5801) );
  OAI21X1 U12544 ( .A(n10916), .B(n10801), .C(n1746), .Y(n5802) );
  OAI21X1 U12545 ( .A(n10918), .B(n10801), .C(n412), .Y(n5803) );
  OAI21X1 U12546 ( .A(n10920), .B(n10801), .C(n519), .Y(n5804) );
  OAI21X1 U12547 ( .A(n10922), .B(n10801), .C(n198), .Y(n5805) );
  OAI21X1 U12548 ( .A(n10924), .B(n10801), .C(n305), .Y(n5806) );
  OAI21X1 U12549 ( .A(n10926), .B(n10801), .C(n841), .Y(n5807) );
  OAI21X1 U12550 ( .A(n10928), .B(n10801), .C(n1319), .Y(n5808) );
  OAI21X1 U12551 ( .A(n10930), .B(n10801), .C(n1445), .Y(n5809) );
  OAI21X1 U12552 ( .A(n10932), .B(n10801), .C(n1069), .Y(n5810) );
  OAI21X1 U12553 ( .A(n10934), .B(n10801), .C(n1194), .Y(n5811) );
  OAI21X1 U12554 ( .A(n10936), .B(n10801), .C(n1903), .Y(n5812) );
  OAI21X1 U12555 ( .A(n10938), .B(n10801), .C(n2060), .Y(n5813) );
  OAI21X1 U12556 ( .A(n10940), .B(n10801), .C(n1586), .Y(n5814) );
  OAI21X1 U12557 ( .A(n10942), .B(n10801), .C(n1745), .Y(n5815) );
  OAI21X1 U12558 ( .A(n10944), .B(n10801), .C(n411), .Y(n5816) );
  OAI21X1 U12559 ( .A(n10946), .B(n10801), .C(n518), .Y(n5817) );
  OAI21X1 U12560 ( .A(n10948), .B(n10801), .C(n197), .Y(n5818) );
  OAI21X1 U12561 ( .A(n10950), .B(n10801), .C(n304), .Y(n5819) );
  OAI21X1 U12562 ( .A(n10954), .B(n10801), .C(n840), .Y(n5820) );
  OAI21X1 U12563 ( .A(n1269), .B(n1837), .C(n10956), .Y(n12303) );
  OAI21X1 U12564 ( .A(n10826), .B(n10803), .C(n1193), .Y(n5821) );
  OAI21X1 U12565 ( .A(n10828), .B(n10803), .C(n1068), .Y(n5822) );
  OAI21X1 U12566 ( .A(n10830), .B(n10803), .C(n1444), .Y(n5823) );
  OAI21X1 U12567 ( .A(n10832), .B(n10803), .C(n1318), .Y(n5824) );
  OAI21X1 U12568 ( .A(n10834), .B(n10803), .C(n1744), .Y(n5825) );
  OAI21X1 U12569 ( .A(n10836), .B(n10803), .C(n1585), .Y(n5826) );
  OAI21X1 U12570 ( .A(n10838), .B(n10803), .C(n2059), .Y(n5827) );
  OAI21X1 U12571 ( .A(n10840), .B(n10803), .C(n1902), .Y(n5828) );
  OAI21X1 U12572 ( .A(n10842), .B(n10803), .C(n303), .Y(n5829) );
  OAI21X1 U12573 ( .A(n10844), .B(n10803), .C(n196), .Y(n5830) );
  OAI21X1 U12574 ( .A(n10846), .B(n10803), .C(n517), .Y(n5831) );
  OAI21X1 U12575 ( .A(n10848), .B(n10803), .C(n410), .Y(n5832) );
  OAI21X1 U12576 ( .A(n10850), .B(n10803), .C(n1192), .Y(n5833) );
  OAI21X1 U12577 ( .A(n10852), .B(n10803), .C(n1067), .Y(n5834) );
  OAI21X1 U12578 ( .A(n10854), .B(n10803), .C(n1443), .Y(n5835) );
  OAI21X1 U12579 ( .A(n10856), .B(n10803), .C(n1317), .Y(n5836) );
  OAI21X1 U12580 ( .A(n10858), .B(n10803), .C(n1743), .Y(n5837) );
  OAI21X1 U12581 ( .A(n10860), .B(n10803), .C(n1584), .Y(n5838) );
  OAI21X1 U12582 ( .A(n10862), .B(n10803), .C(n2058), .Y(n5839) );
  OAI21X1 U12583 ( .A(n10864), .B(n10803), .C(n1901), .Y(n5840) );
  OAI21X1 U12584 ( .A(n10866), .B(n10803), .C(n302), .Y(n5841) );
  OAI21X1 U12585 ( .A(n10868), .B(n10803), .C(n195), .Y(n5842) );
  OAI21X1 U12586 ( .A(n10870), .B(n10803), .C(n516), .Y(n5843) );
  OAI21X1 U12587 ( .A(n10872), .B(n10803), .C(n409), .Y(n5844) );
  OAI21X1 U12588 ( .A(n10874), .B(n10803), .C(n731), .Y(n5845) );
  OAI21X1 U12589 ( .A(n10876), .B(n10803), .C(n1191), .Y(n5846) );
  OAI21X1 U12590 ( .A(n10878), .B(n10803), .C(n1066), .Y(n5847) );
  OAI21X1 U12591 ( .A(n10880), .B(n10803), .C(n1442), .Y(n5848) );
  OAI21X1 U12592 ( .A(n10882), .B(n10803), .C(n1316), .Y(n5849) );
  OAI21X1 U12593 ( .A(n10884), .B(n10803), .C(n1742), .Y(n5850) );
  OAI21X1 U12594 ( .A(n10886), .B(n10803), .C(n1583), .Y(n5851) );
  OAI21X1 U12595 ( .A(n10888), .B(n10803), .C(n2057), .Y(n5852) );
  OAI21X1 U12596 ( .A(n10890), .B(n10803), .C(n1900), .Y(n5853) );
  OAI21X1 U12597 ( .A(n10892), .B(n10803), .C(n301), .Y(n5854) );
  OAI21X1 U12598 ( .A(n10894), .B(n10803), .C(n194), .Y(n5855) );
  OAI21X1 U12599 ( .A(n10896), .B(n10803), .C(n515), .Y(n5856) );
  OAI21X1 U12600 ( .A(n10898), .B(n10803), .C(n408), .Y(n5857) );
  OAI21X1 U12601 ( .A(n10900), .B(n10803), .C(n730), .Y(n5858) );
  OAI21X1 U12602 ( .A(n10902), .B(n10803), .C(n1190), .Y(n5859) );
  OAI21X1 U12603 ( .A(n10904), .B(n10803), .C(n1065), .Y(n5860) );
  OAI21X1 U12604 ( .A(n10906), .B(n10803), .C(n1441), .Y(n5861) );
  OAI21X1 U12605 ( .A(n10908), .B(n10803), .C(n1315), .Y(n5862) );
  OAI21X1 U12606 ( .A(n10910), .B(n10803), .C(n1741), .Y(n5863) );
  OAI21X1 U12607 ( .A(n10912), .B(n10803), .C(n1582), .Y(n5864) );
  OAI21X1 U12608 ( .A(n10914), .B(n10803), .C(n2056), .Y(n5865) );
  OAI21X1 U12609 ( .A(n10916), .B(n10803), .C(n1899), .Y(n5866) );
  OAI21X1 U12610 ( .A(n10918), .B(n10803), .C(n300), .Y(n5867) );
  OAI21X1 U12611 ( .A(n10920), .B(n10803), .C(n193), .Y(n5868) );
  OAI21X1 U12612 ( .A(n10922), .B(n10803), .C(n514), .Y(n5869) );
  OAI21X1 U12613 ( .A(n10924), .B(n10803), .C(n407), .Y(n5870) );
  OAI21X1 U12614 ( .A(n10926), .B(n10803), .C(n729), .Y(n5871) );
  OAI21X1 U12615 ( .A(n10928), .B(n10803), .C(n1189), .Y(n5872) );
  OAI21X1 U12616 ( .A(n10930), .B(n10803), .C(n1064), .Y(n5873) );
  OAI21X1 U12617 ( .A(n10932), .B(n10803), .C(n1440), .Y(n5874) );
  OAI21X1 U12618 ( .A(n10934), .B(n10803), .C(n1314), .Y(n5875) );
  OAI21X1 U12619 ( .A(n10936), .B(n10803), .C(n1740), .Y(n5876) );
  OAI21X1 U12620 ( .A(n10938), .B(n10803), .C(n1581), .Y(n5877) );
  OAI21X1 U12621 ( .A(n10940), .B(n10803), .C(n2055), .Y(n5878) );
  OAI21X1 U12622 ( .A(n10942), .B(n10803), .C(n1898), .Y(n5879) );
  OAI21X1 U12623 ( .A(n10944), .B(n10803), .C(n299), .Y(n5880) );
  OAI21X1 U12624 ( .A(n10946), .B(n10803), .C(n192), .Y(n5881) );
  OAI21X1 U12625 ( .A(n10948), .B(n10803), .C(n513), .Y(n5882) );
  OAI21X1 U12626 ( .A(n10950), .B(n10803), .C(n406), .Y(n5883) );
  OAI21X1 U12627 ( .A(n10954), .B(n10803), .C(n728), .Y(n5884) );
  OAI21X1 U12628 ( .A(n1144), .B(n1837), .C(n10956), .Y(n12369) );
  OAI21X1 U12629 ( .A(n10826), .B(n10805), .C(n1063), .Y(n5885) );
  OAI21X1 U12630 ( .A(n10828), .B(n10805), .C(n1188), .Y(n5886) );
  OAI21X1 U12631 ( .A(n10830), .B(n10805), .C(n1313), .Y(n5887) );
  OAI21X1 U12632 ( .A(n10832), .B(n10805), .C(n1439), .Y(n5888) );
  OAI21X1 U12633 ( .A(n10834), .B(n10805), .C(n1580), .Y(n5889) );
  OAI21X1 U12634 ( .A(n10836), .B(n10805), .C(n1739), .Y(n5890) );
  OAI21X1 U12635 ( .A(n10838), .B(n10805), .C(n1897), .Y(n5891) );
  OAI21X1 U12636 ( .A(n10840), .B(n10805), .C(n2054), .Y(n5892) );
  OAI21X1 U12637 ( .A(n10842), .B(n10805), .C(n191), .Y(n5893) );
  OAI21X1 U12638 ( .A(n10844), .B(n10805), .C(n298), .Y(n5894) );
  OAI21X1 U12639 ( .A(n10846), .B(n10805), .C(n405), .Y(n5895) );
  OAI21X1 U12640 ( .A(n10848), .B(n10805), .C(n512), .Y(n5896) );
  OAI21X1 U12641 ( .A(n10850), .B(n10805), .C(n1062), .Y(n5897) );
  OAI21X1 U12642 ( .A(n10852), .B(n10805), .C(n1187), .Y(n5898) );
  OAI21X1 U12643 ( .A(n10854), .B(n10805), .C(n1312), .Y(n5899) );
  OAI21X1 U12644 ( .A(n10856), .B(n10805), .C(n1438), .Y(n5900) );
  OAI21X1 U12645 ( .A(n10858), .B(n10805), .C(n1579), .Y(n5901) );
  OAI21X1 U12646 ( .A(n10860), .B(n10805), .C(n1738), .Y(n5902) );
  OAI21X1 U12647 ( .A(n10862), .B(n10805), .C(n1896), .Y(n5903) );
  OAI21X1 U12648 ( .A(n10864), .B(n10805), .C(n2053), .Y(n5904) );
  OAI21X1 U12649 ( .A(n10866), .B(n10805), .C(n190), .Y(n5905) );
  OAI21X1 U12650 ( .A(n10868), .B(n10805), .C(n297), .Y(n5906) );
  OAI21X1 U12651 ( .A(n10870), .B(n10805), .C(n404), .Y(n5907) );
  OAI21X1 U12652 ( .A(n10872), .B(n10805), .C(n511), .Y(n5908) );
  OAI21X1 U12653 ( .A(n10874), .B(n10805), .C(n619), .Y(n5909) );
  OAI21X1 U12654 ( .A(n10876), .B(n10805), .C(n1061), .Y(n5910) );
  OAI21X1 U12655 ( .A(n10878), .B(n10805), .C(n1186), .Y(n5911) );
  OAI21X1 U12656 ( .A(n10880), .B(n10805), .C(n1311), .Y(n5912) );
  OAI21X1 U12657 ( .A(n10882), .B(n10805), .C(n1437), .Y(n5913) );
  OAI21X1 U12658 ( .A(n10884), .B(n10805), .C(n1578), .Y(n5914) );
  OAI21X1 U12659 ( .A(n10886), .B(n10805), .C(n1737), .Y(n5915) );
  OAI21X1 U12660 ( .A(n10888), .B(n10805), .C(n1895), .Y(n5916) );
  OAI21X1 U12661 ( .A(n10890), .B(n10805), .C(n2052), .Y(n5917) );
  OAI21X1 U12662 ( .A(n10892), .B(n10805), .C(n189), .Y(n5918) );
  OAI21X1 U12663 ( .A(n10894), .B(n10805), .C(n296), .Y(n5919) );
  OAI21X1 U12664 ( .A(n10896), .B(n10805), .C(n403), .Y(n5920) );
  OAI21X1 U12665 ( .A(n10898), .B(n10805), .C(n510), .Y(n5921) );
  OAI21X1 U12666 ( .A(n10900), .B(n10805), .C(n618), .Y(n5922) );
  OAI21X1 U12667 ( .A(n10902), .B(n10805), .C(n1060), .Y(n5923) );
  OAI21X1 U12668 ( .A(n10904), .B(n10805), .C(n1185), .Y(n5924) );
  OAI21X1 U12669 ( .A(n10906), .B(n10805), .C(n1310), .Y(n5925) );
  OAI21X1 U12670 ( .A(n10908), .B(n10805), .C(n1436), .Y(n5926) );
  OAI21X1 U12671 ( .A(n10910), .B(n10805), .C(n1577), .Y(n5927) );
  OAI21X1 U12672 ( .A(n10912), .B(n10805), .C(n1736), .Y(n5928) );
  OAI21X1 U12673 ( .A(n10914), .B(n10805), .C(n1894), .Y(n5929) );
  OAI21X1 U12674 ( .A(n10916), .B(n10805), .C(n2051), .Y(n5930) );
  OAI21X1 U12675 ( .A(n10918), .B(n10805), .C(n188), .Y(n5931) );
  OAI21X1 U12676 ( .A(n10920), .B(n10805), .C(n295), .Y(n5932) );
  OAI21X1 U12677 ( .A(n10922), .B(n10805), .C(n402), .Y(n5933) );
  OAI21X1 U12678 ( .A(n10924), .B(n10805), .C(n509), .Y(n5934) );
  OAI21X1 U12679 ( .A(n10926), .B(n10805), .C(n617), .Y(n5935) );
  OAI21X1 U12680 ( .A(n10928), .B(n10805), .C(n1059), .Y(n5936) );
  OAI21X1 U12681 ( .A(n10930), .B(n10805), .C(n1184), .Y(n5937) );
  OAI21X1 U12682 ( .A(n10932), .B(n10805), .C(n1309), .Y(n5938) );
  OAI21X1 U12683 ( .A(n10934), .B(n10805), .C(n1435), .Y(n5939) );
  OAI21X1 U12684 ( .A(n10936), .B(n10805), .C(n1576), .Y(n5940) );
  OAI21X1 U12685 ( .A(n10938), .B(n10805), .C(n1735), .Y(n5941) );
  OAI21X1 U12686 ( .A(n10940), .B(n10805), .C(n1893), .Y(n5942) );
  OAI21X1 U12687 ( .A(n10942), .B(n10805), .C(n2050), .Y(n5943) );
  OAI21X1 U12688 ( .A(n10944), .B(n10805), .C(n187), .Y(n5944) );
  OAI21X1 U12689 ( .A(n10946), .B(n10805), .C(n294), .Y(n5945) );
  OAI21X1 U12690 ( .A(n10948), .B(n10805), .C(n401), .Y(n5946) );
  OAI21X1 U12691 ( .A(n10950), .B(n10805), .C(n508), .Y(n5947) );
  OAI21X1 U12692 ( .A(n10954), .B(n10805), .C(n616), .Y(n5948) );
  OAI21X1 U12693 ( .A(n1143), .B(n1837), .C(n10956), .Y(n12435) );
  OAI21X1 U12694 ( .A(n10826), .B(n10807), .C(n951), .Y(n5949) );
  OAI21X1 U12695 ( .A(n10828), .B(n10807), .C(n839), .Y(n5950) );
  OAI21X1 U12696 ( .A(n10830), .B(n10807), .C(n727), .Y(n5951) );
  OAI21X1 U12697 ( .A(n10832), .B(n10807), .C(n615), .Y(n5952) );
  OAI21X1 U12698 ( .A(n10834), .B(n10807), .C(n507), .Y(n5953) );
  OAI21X1 U12699 ( .A(n10836), .B(n10807), .C(n400), .Y(n5954) );
  OAI21X1 U12700 ( .A(n10838), .B(n10807), .C(n293), .Y(n5955) );
  OAI21X1 U12701 ( .A(n10840), .B(n10807), .C(n122), .Y(n5956) );
  OAI21X1 U12702 ( .A(n10842), .B(n10807), .C(n2049), .Y(n5957) );
  OAI21X1 U12703 ( .A(n10844), .B(n10807), .C(n1892), .Y(n5958) );
  OAI21X1 U12704 ( .A(n10846), .B(n10807), .C(n1734), .Y(n5959) );
  OAI21X1 U12705 ( .A(n10848), .B(n10807), .C(n1575), .Y(n5960) );
  OAI21X1 U12706 ( .A(n10850), .B(n10807), .C(n950), .Y(n5961) );
  OAI21X1 U12707 ( .A(n10852), .B(n10807), .C(n838), .Y(n5962) );
  OAI21X1 U12708 ( .A(n10854), .B(n10807), .C(n726), .Y(n5963) );
  OAI21X1 U12709 ( .A(n10856), .B(n10807), .C(n614), .Y(n5964) );
  OAI21X1 U12710 ( .A(n10858), .B(n10807), .C(n506), .Y(n5965) );
  OAI21X1 U12711 ( .A(n10860), .B(n10807), .C(n399), .Y(n5966) );
  OAI21X1 U12712 ( .A(n10862), .B(n10807), .C(n292), .Y(n5967) );
  OAI21X1 U12713 ( .A(n10864), .B(n10807), .C(n121), .Y(n5968) );
  OAI21X1 U12714 ( .A(n10866), .B(n10807), .C(n2048), .Y(n5969) );
  OAI21X1 U12715 ( .A(n10868), .B(n10807), .C(n1891), .Y(n5970) );
  OAI21X1 U12716 ( .A(n10870), .B(n10807), .C(n1733), .Y(n5971) );
  OAI21X1 U12717 ( .A(n10872), .B(n10807), .C(n1574), .Y(n5972) );
  OAI21X1 U12718 ( .A(n10874), .B(n10807), .C(n1434), .Y(n5973) );
  OAI21X1 U12719 ( .A(n10876), .B(n10807), .C(n949), .Y(n5974) );
  OAI21X1 U12720 ( .A(n10878), .B(n10807), .C(n837), .Y(n5975) );
  OAI21X1 U12721 ( .A(n10880), .B(n10807), .C(n725), .Y(n5976) );
  OAI21X1 U12722 ( .A(n10882), .B(n10807), .C(n613), .Y(n5977) );
  OAI21X1 U12723 ( .A(n10884), .B(n10807), .C(n505), .Y(n5978) );
  OAI21X1 U12724 ( .A(n10886), .B(n10807), .C(n398), .Y(n5979) );
  OAI21X1 U12725 ( .A(n10888), .B(n10807), .C(n291), .Y(n5980) );
  OAI21X1 U12726 ( .A(n10890), .B(n10807), .C(n120), .Y(n5981) );
  OAI21X1 U12727 ( .A(n10892), .B(n10807), .C(n2047), .Y(n5982) );
  OAI21X1 U12728 ( .A(n10894), .B(n10807), .C(n1890), .Y(n5983) );
  OAI21X1 U12729 ( .A(n10896), .B(n10807), .C(n1732), .Y(n5984) );
  OAI21X1 U12730 ( .A(n10898), .B(n10807), .C(n1573), .Y(n5985) );
  OAI21X1 U12731 ( .A(n10900), .B(n10807), .C(n1433), .Y(n5986) );
  OAI21X1 U12732 ( .A(n10902), .B(n10807), .C(n948), .Y(n5987) );
  OAI21X1 U12733 ( .A(n10904), .B(n10807), .C(n836), .Y(n5988) );
  OAI21X1 U12734 ( .A(n10906), .B(n10807), .C(n724), .Y(n5989) );
  OAI21X1 U12735 ( .A(n10908), .B(n10807), .C(n612), .Y(n5990) );
  OAI21X1 U12736 ( .A(n10910), .B(n10807), .C(n504), .Y(n5991) );
  OAI21X1 U12737 ( .A(n10912), .B(n10807), .C(n397), .Y(n5992) );
  OAI21X1 U12738 ( .A(n10914), .B(n10807), .C(n290), .Y(n5993) );
  OAI21X1 U12739 ( .A(n10916), .B(n10807), .C(n55), .Y(n5994) );
  OAI21X1 U12740 ( .A(n10918), .B(n10807), .C(n2046), .Y(n5995) );
  OAI21X1 U12741 ( .A(n10920), .B(n10807), .C(n1889), .Y(n5996) );
  OAI21X1 U12742 ( .A(n10922), .B(n10807), .C(n1731), .Y(n5997) );
  OAI21X1 U12743 ( .A(n10924), .B(n10807), .C(n1572), .Y(n5998) );
  OAI21X1 U12744 ( .A(n10926), .B(n10807), .C(n1432), .Y(n5999) );
  OAI21X1 U12745 ( .A(n10928), .B(n10807), .C(n947), .Y(n6000) );
  OAI21X1 U12746 ( .A(n10930), .B(n10807), .C(n835), .Y(n6001) );
  OAI21X1 U12747 ( .A(n10932), .B(n10807), .C(n723), .Y(n6002) );
  OAI21X1 U12748 ( .A(n10934), .B(n10807), .C(n611), .Y(n6003) );
  OAI21X1 U12749 ( .A(n10936), .B(n10807), .C(n503), .Y(n6004) );
  OAI21X1 U12750 ( .A(n10938), .B(n10807), .C(n396), .Y(n6005) );
  OAI21X1 U12751 ( .A(n10940), .B(n10807), .C(n289), .Y(n6006) );
  OAI21X1 U12752 ( .A(n10942), .B(n10807), .C(n54), .Y(n6007) );
  OAI21X1 U12753 ( .A(n10944), .B(n10807), .C(n2045), .Y(n6008) );
  OAI21X1 U12754 ( .A(n10946), .B(n10807), .C(n1888), .Y(n6009) );
  OAI21X1 U12755 ( .A(n10948), .B(n10807), .C(n1730), .Y(n6010) );
  OAI21X1 U12756 ( .A(n10950), .B(n10807), .C(n1571), .Y(n6011) );
  OAI21X1 U12757 ( .A(n10954), .B(n10807), .C(n1431), .Y(n6012) );
  OAI21X1 U12758 ( .A(n1268), .B(n1837), .C(n10956), .Y(n12501) );
  OAI21X1 U12759 ( .A(n10826), .B(n10809), .C(n834), .Y(n6013) );
  OAI21X1 U12760 ( .A(n10828), .B(n10809), .C(n946), .Y(n6014) );
  OAI21X1 U12761 ( .A(n10830), .B(n10809), .C(n610), .Y(n6015) );
  OAI21X1 U12762 ( .A(n10832), .B(n10809), .C(n722), .Y(n6016) );
  OAI21X1 U12763 ( .A(n10834), .B(n10809), .C(n395), .Y(n6017) );
  OAI21X1 U12764 ( .A(n10836), .B(n10809), .C(n502), .Y(n6018) );
  OAI21X1 U12765 ( .A(n10838), .B(n10809), .C(n53), .Y(n6019) );
  OAI21X1 U12766 ( .A(n10840), .B(n10809), .C(n288), .Y(n6020) );
  OAI21X1 U12767 ( .A(n10842), .B(n10809), .C(n1887), .Y(n6021) );
  OAI21X1 U12768 ( .A(n10844), .B(n10809), .C(n2044), .Y(n6022) );
  OAI21X1 U12769 ( .A(n10846), .B(n10809), .C(n1570), .Y(n6023) );
  OAI21X1 U12770 ( .A(n10848), .B(n10809), .C(n1729), .Y(n6024) );
  OAI21X1 U12771 ( .A(n10850), .B(n10809), .C(n833), .Y(n6025) );
  OAI21X1 U12772 ( .A(n10852), .B(n10809), .C(n945), .Y(n6026) );
  OAI21X1 U12773 ( .A(n10854), .B(n10809), .C(n609), .Y(n6027) );
  OAI21X1 U12774 ( .A(n10856), .B(n10809), .C(n721), .Y(n6028) );
  OAI21X1 U12775 ( .A(n10858), .B(n10809), .C(n394), .Y(n6029) );
  OAI21X1 U12776 ( .A(n10860), .B(n10809), .C(n501), .Y(n6030) );
  OAI21X1 U12777 ( .A(n10862), .B(n10809), .C(n52), .Y(n6031) );
  OAI21X1 U12778 ( .A(n10864), .B(n10809), .C(n287), .Y(n6032) );
  OAI21X1 U12779 ( .A(n10866), .B(n10809), .C(n1886), .Y(n6033) );
  OAI21X1 U12780 ( .A(n10868), .B(n10809), .C(n2043), .Y(n6034) );
  OAI21X1 U12781 ( .A(n10870), .B(n10809), .C(n1569), .Y(n6035) );
  OAI21X1 U12782 ( .A(n10872), .B(n10809), .C(n1728), .Y(n6036) );
  OAI21X1 U12783 ( .A(n10874), .B(n10809), .C(n1308), .Y(n6037) );
  OAI21X1 U12784 ( .A(n10876), .B(n10809), .C(n832), .Y(n6038) );
  OAI21X1 U12785 ( .A(n10878), .B(n10809), .C(n944), .Y(n6039) );
  OAI21X1 U12786 ( .A(n10880), .B(n10809), .C(n608), .Y(n6040) );
  OAI21X1 U12787 ( .A(n10882), .B(n10809), .C(n720), .Y(n6041) );
  OAI21X1 U12788 ( .A(n10884), .B(n10809), .C(n393), .Y(n6042) );
  OAI21X1 U12789 ( .A(n10886), .B(n10809), .C(n500), .Y(n6043) );
  OAI21X1 U12790 ( .A(n10888), .B(n10809), .C(n51), .Y(n6044) );
  OAI21X1 U12791 ( .A(n10890), .B(n10809), .C(n286), .Y(n6045) );
  OAI21X1 U12792 ( .A(n10892), .B(n10809), .C(n1885), .Y(n6046) );
  OAI21X1 U12793 ( .A(n10894), .B(n10809), .C(n2042), .Y(n6047) );
  OAI21X1 U12794 ( .A(n10896), .B(n10809), .C(n1568), .Y(n6048) );
  OAI21X1 U12795 ( .A(n10898), .B(n10809), .C(n1727), .Y(n6049) );
  OAI21X1 U12796 ( .A(n10900), .B(n10809), .C(n1307), .Y(n6050) );
  OAI21X1 U12797 ( .A(n10902), .B(n10809), .C(n831), .Y(n6051) );
  OAI21X1 U12798 ( .A(n10904), .B(n10809), .C(n943), .Y(n6052) );
  OAI21X1 U12799 ( .A(n10906), .B(n10809), .C(n607), .Y(n6053) );
  OAI21X1 U12800 ( .A(n10908), .B(n10809), .C(n719), .Y(n6054) );
  OAI21X1 U12801 ( .A(n10910), .B(n10809), .C(n392), .Y(n6055) );
  OAI21X1 U12802 ( .A(n10912), .B(n10809), .C(n499), .Y(n6056) );
  OAI21X1 U12803 ( .A(n10914), .B(n10809), .C(n50), .Y(n6057) );
  OAI21X1 U12804 ( .A(n10916), .B(n10809), .C(n285), .Y(n6058) );
  OAI21X1 U12805 ( .A(n10918), .B(n10809), .C(n1884), .Y(n6059) );
  OAI21X1 U12806 ( .A(n10920), .B(n10809), .C(n2041), .Y(n6060) );
  OAI21X1 U12807 ( .A(n10922), .B(n10809), .C(n1567), .Y(n6061) );
  OAI21X1 U12808 ( .A(n10924), .B(n10809), .C(n1726), .Y(n6062) );
  OAI21X1 U12809 ( .A(n10926), .B(n10809), .C(n1306), .Y(n6063) );
  OAI21X1 U12810 ( .A(n10928), .B(n10809), .C(n830), .Y(n6064) );
  OAI21X1 U12811 ( .A(n10930), .B(n10809), .C(n942), .Y(n6065) );
  OAI21X1 U12812 ( .A(n10932), .B(n10809), .C(n606), .Y(n6066) );
  OAI21X1 U12813 ( .A(n10934), .B(n10809), .C(n718), .Y(n6067) );
  OAI21X1 U12814 ( .A(n10936), .B(n10809), .C(n391), .Y(n6068) );
  OAI21X1 U12815 ( .A(n10938), .B(n10809), .C(n498), .Y(n6069) );
  OAI21X1 U12816 ( .A(n10940), .B(n10809), .C(n49), .Y(n6070) );
  OAI21X1 U12817 ( .A(n10942), .B(n10809), .C(n284), .Y(n6071) );
  OAI21X1 U12818 ( .A(n10944), .B(n10809), .C(n1883), .Y(n6072) );
  OAI21X1 U12819 ( .A(n10946), .B(n10809), .C(n2040), .Y(n6073) );
  OAI21X1 U12820 ( .A(n10948), .B(n10809), .C(n1566), .Y(n6074) );
  OAI21X1 U12821 ( .A(n10950), .B(n10809), .C(n1725), .Y(n6075) );
  OAI21X1 U12822 ( .A(n10954), .B(n10809), .C(n1305), .Y(n6076) );
  OAI21X1 U12823 ( .A(n1394), .B(n1837), .C(n10956), .Y(n12567) );
  OAI21X1 U12824 ( .A(n10826), .B(n10811), .C(n717), .Y(n6077) );
  OAI21X1 U12825 ( .A(n10828), .B(n10811), .C(n605), .Y(n6078) );
  OAI21X1 U12826 ( .A(n10830), .B(n10811), .C(n941), .Y(n6079) );
  OAI21X1 U12827 ( .A(n10832), .B(n10811), .C(n829), .Y(n6080) );
  OAI21X1 U12828 ( .A(n10834), .B(n10811), .C(n283), .Y(n6081) );
  OAI21X1 U12829 ( .A(n10836), .B(n10811), .C(n48), .Y(n6082) );
  OAI21X1 U12830 ( .A(n10838), .B(n10811), .C(n497), .Y(n6083) );
  OAI21X1 U12831 ( .A(n10840), .B(n10811), .C(n390), .Y(n6084) );
  OAI21X1 U12832 ( .A(n10842), .B(n10811), .C(n1724), .Y(n6085) );
  OAI21X1 U12833 ( .A(n10844), .B(n10811), .C(n1565), .Y(n6086) );
  OAI21X1 U12834 ( .A(n10846), .B(n10811), .C(n2039), .Y(n6087) );
  OAI21X1 U12835 ( .A(n10848), .B(n10811), .C(n1882), .Y(n6088) );
  OAI21X1 U12836 ( .A(n10850), .B(n10811), .C(n716), .Y(n6089) );
  OAI21X1 U12837 ( .A(n10852), .B(n10811), .C(n604), .Y(n6090) );
  OAI21X1 U12838 ( .A(n10854), .B(n10811), .C(n940), .Y(n6091) );
  OAI21X1 U12839 ( .A(n10856), .B(n10811), .C(n828), .Y(n6092) );
  OAI21X1 U12840 ( .A(n10858), .B(n10811), .C(n282), .Y(n6093) );
  OAI21X1 U12841 ( .A(n10860), .B(n10811), .C(n47), .Y(n6094) );
  OAI21X1 U12842 ( .A(n10862), .B(n10811), .C(n496), .Y(n6095) );
  OAI21X1 U12843 ( .A(n10864), .B(n10811), .C(n389), .Y(n6096) );
  OAI21X1 U12844 ( .A(n10866), .B(n10811), .C(n1723), .Y(n6097) );
  OAI21X1 U12845 ( .A(n10868), .B(n10811), .C(n1564), .Y(n6098) );
  OAI21X1 U12846 ( .A(n10870), .B(n10811), .C(n2038), .Y(n6099) );
  OAI21X1 U12847 ( .A(n10872), .B(n10811), .C(n1881), .Y(n6100) );
  OAI21X1 U12848 ( .A(n10874), .B(n10811), .C(n1183), .Y(n6101) );
  OAI21X1 U12849 ( .A(n10876), .B(n10811), .C(n715), .Y(n6102) );
  OAI21X1 U12850 ( .A(n10878), .B(n10811), .C(n603), .Y(n6103) );
  OAI21X1 U12851 ( .A(n10880), .B(n10811), .C(n939), .Y(n6104) );
  OAI21X1 U12852 ( .A(n10882), .B(n10811), .C(n827), .Y(n6105) );
  OAI21X1 U12853 ( .A(n10884), .B(n10811), .C(n281), .Y(n6106) );
  OAI21X1 U12854 ( .A(n10886), .B(n10811), .C(n46), .Y(n6107) );
  OAI21X1 U12855 ( .A(n10888), .B(n10811), .C(n495), .Y(n6108) );
  OAI21X1 U12856 ( .A(n10890), .B(n10811), .C(n388), .Y(n6109) );
  OAI21X1 U12857 ( .A(n10892), .B(n10811), .C(n1722), .Y(n6110) );
  OAI21X1 U12858 ( .A(n10894), .B(n10811), .C(n1563), .Y(n6111) );
  OAI21X1 U12859 ( .A(n10896), .B(n10811), .C(n2037), .Y(n6112) );
  OAI21X1 U12860 ( .A(n10898), .B(n10811), .C(n1880), .Y(n6113) );
  OAI21X1 U12861 ( .A(n10900), .B(n10811), .C(n1182), .Y(n6114) );
  OAI21X1 U12862 ( .A(n10902), .B(n10811), .C(n714), .Y(n6115) );
  OAI21X1 U12863 ( .A(n10904), .B(n10811), .C(n602), .Y(n6116) );
  OAI21X1 U12864 ( .A(n10906), .B(n10811), .C(n938), .Y(n6117) );
  OAI21X1 U12865 ( .A(n10908), .B(n10811), .C(n826), .Y(n6118) );
  OAI21X1 U12866 ( .A(n10910), .B(n10811), .C(n280), .Y(n6119) );
  OAI21X1 U12867 ( .A(n10912), .B(n10811), .C(n45), .Y(n6120) );
  OAI21X1 U12868 ( .A(n10914), .B(n10811), .C(n494), .Y(n6121) );
  OAI21X1 U12869 ( .A(n10916), .B(n10811), .C(n387), .Y(n6122) );
  OAI21X1 U12870 ( .A(n10918), .B(n10811), .C(n1721), .Y(n6123) );
  OAI21X1 U12871 ( .A(n10920), .B(n10811), .C(n1562), .Y(n6124) );
  OAI21X1 U12872 ( .A(n10922), .B(n10811), .C(n2036), .Y(n6125) );
  OAI21X1 U12873 ( .A(n10924), .B(n10811), .C(n1879), .Y(n6126) );
  OAI21X1 U12874 ( .A(n10926), .B(n10811), .C(n1181), .Y(n6127) );
  OAI21X1 U12875 ( .A(n10928), .B(n10811), .C(n713), .Y(n6128) );
  OAI21X1 U12876 ( .A(n10930), .B(n10811), .C(n601), .Y(n6129) );
  OAI21X1 U12877 ( .A(n10932), .B(n10811), .C(n937), .Y(n6130) );
  OAI21X1 U12878 ( .A(n10934), .B(n10811), .C(n825), .Y(n6131) );
  OAI21X1 U12879 ( .A(n10936), .B(n10811), .C(n279), .Y(n6132) );
  OAI21X1 U12880 ( .A(n10938), .B(n10811), .C(n44), .Y(n6133) );
  OAI21X1 U12881 ( .A(n10940), .B(n10811), .C(n493), .Y(n6134) );
  OAI21X1 U12882 ( .A(n10942), .B(n10811), .C(n386), .Y(n6135) );
  OAI21X1 U12883 ( .A(n10944), .B(n10811), .C(n1720), .Y(n6136) );
  OAI21X1 U12884 ( .A(n10946), .B(n10811), .C(n1561), .Y(n6137) );
  OAI21X1 U12885 ( .A(n10948), .B(n10811), .C(n2035), .Y(n6138) );
  OAI21X1 U12886 ( .A(n10950), .B(n10811), .C(n1878), .Y(n6139) );
  OAI21X1 U12887 ( .A(n10954), .B(n10811), .C(n1180), .Y(n6140) );
  OAI21X1 U12888 ( .A(n1678), .B(n1837), .C(n10956), .Y(n12634) );
  OAI21X1 U12889 ( .A(n10826), .B(n10813), .C(n600), .Y(n6141) );
  OAI21X1 U12890 ( .A(n10828), .B(n10813), .C(n712), .Y(n6142) );
  OAI21X1 U12891 ( .A(n10830), .B(n10813), .C(n824), .Y(n6143) );
  OAI21X1 U12892 ( .A(n10832), .B(n10813), .C(n936), .Y(n6144) );
  OAI21X1 U12893 ( .A(n10834), .B(n10813), .C(n43), .Y(n6145) );
  OAI21X1 U12894 ( .A(n10836), .B(n10813), .C(n278), .Y(n6146) );
  OAI21X1 U12895 ( .A(n10838), .B(n10813), .C(n385), .Y(n6147) );
  OAI21X1 U12896 ( .A(n10840), .B(n10813), .C(n492), .Y(n6148) );
  OAI21X1 U12897 ( .A(n10842), .B(n10813), .C(n1560), .Y(n6149) );
  OAI21X1 U12898 ( .A(n10844), .B(n10813), .C(n1719), .Y(n6150) );
  OAI21X1 U12899 ( .A(n10846), .B(n10813), .C(n1877), .Y(n6151) );
  OAI21X1 U12900 ( .A(n10848), .B(n10813), .C(n2034), .Y(n6152) );
  OAI21X1 U12901 ( .A(n10850), .B(n10813), .C(n599), .Y(n6153) );
  OAI21X1 U12902 ( .A(n10852), .B(n10813), .C(n711), .Y(n6154) );
  OAI21X1 U12903 ( .A(n10854), .B(n10813), .C(n823), .Y(n6155) );
  OAI21X1 U12904 ( .A(n10856), .B(n10813), .C(n935), .Y(n6156) );
  OAI21X1 U12905 ( .A(n10858), .B(n10813), .C(n42), .Y(n6157) );
  OAI21X1 U12906 ( .A(n10860), .B(n10813), .C(n277), .Y(n6158) );
  OAI21X1 U12907 ( .A(n10862), .B(n10813), .C(n384), .Y(n6159) );
  OAI21X1 U12908 ( .A(n10864), .B(n10813), .C(n491), .Y(n6160) );
  OAI21X1 U12909 ( .A(n10866), .B(n10813), .C(n1559), .Y(n6161) );
  OAI21X1 U12910 ( .A(n10868), .B(n10813), .C(n1718), .Y(n6162) );
  OAI21X1 U12911 ( .A(n10870), .B(n10813), .C(n1876), .Y(n6163) );
  OAI21X1 U12912 ( .A(n10872), .B(n10813), .C(n2033), .Y(n6164) );
  OAI21X1 U12913 ( .A(n10874), .B(n10813), .C(n1058), .Y(n6165) );
  OAI21X1 U12914 ( .A(n10876), .B(n10813), .C(n598), .Y(n6166) );
  OAI21X1 U12915 ( .A(n10878), .B(n10813), .C(n710), .Y(n6167) );
  OAI21X1 U12916 ( .A(n10880), .B(n10813), .C(n822), .Y(n6168) );
  OAI21X1 U12917 ( .A(n10882), .B(n10813), .C(n934), .Y(n6169) );
  OAI21X1 U12918 ( .A(n10884), .B(n10813), .C(n41), .Y(n6170) );
  OAI21X1 U12919 ( .A(n10886), .B(n10813), .C(n276), .Y(n6171) );
  OAI21X1 U12920 ( .A(n10888), .B(n10813), .C(n383), .Y(n6172) );
  OAI21X1 U12921 ( .A(n10890), .B(n10813), .C(n490), .Y(n6173) );
  OAI21X1 U12922 ( .A(n10892), .B(n10813), .C(n1558), .Y(n6174) );
  OAI21X1 U12923 ( .A(n10894), .B(n10813), .C(n1717), .Y(n6175) );
  OAI21X1 U12924 ( .A(n10896), .B(n10813), .C(n1875), .Y(n6176) );
  OAI21X1 U12925 ( .A(n10898), .B(n10813), .C(n2032), .Y(n6177) );
  OAI21X1 U12926 ( .A(n10900), .B(n10813), .C(n1057), .Y(n6178) );
  OAI21X1 U12927 ( .A(n10902), .B(n10813), .C(n597), .Y(n6179) );
  OAI21X1 U12928 ( .A(n10904), .B(n10813), .C(n709), .Y(n6180) );
  OAI21X1 U12929 ( .A(n10906), .B(n10813), .C(n821), .Y(n6181) );
  OAI21X1 U12930 ( .A(n10908), .B(n10813), .C(n933), .Y(n6182) );
  OAI21X1 U12931 ( .A(n10910), .B(n10813), .C(n40), .Y(n6183) );
  OAI21X1 U12932 ( .A(n10912), .B(n10813), .C(n275), .Y(n6184) );
  OAI21X1 U12933 ( .A(n10914), .B(n10813), .C(n382), .Y(n6185) );
  OAI21X1 U12934 ( .A(n10916), .B(n10813), .C(n489), .Y(n6186) );
  OAI21X1 U12935 ( .A(n10918), .B(n10813), .C(n1557), .Y(n6187) );
  OAI21X1 U12936 ( .A(n10920), .B(n10813), .C(n1716), .Y(n6188) );
  OAI21X1 U12937 ( .A(n10922), .B(n10813), .C(n1874), .Y(n6189) );
  OAI21X1 U12938 ( .A(n10924), .B(n10813), .C(n2031), .Y(n6190) );
  OAI21X1 U12939 ( .A(n10926), .B(n10813), .C(n1056), .Y(n6191) );
  OAI21X1 U12940 ( .A(n10928), .B(n10813), .C(n596), .Y(n6192) );
  OAI21X1 U12941 ( .A(n10930), .B(n10813), .C(n708), .Y(n6193) );
  OAI21X1 U12942 ( .A(n10932), .B(n10813), .C(n820), .Y(n6194) );
  OAI21X1 U12943 ( .A(n10934), .B(n10813), .C(n932), .Y(n6195) );
  OAI21X1 U12944 ( .A(n10936), .B(n10813), .C(n39), .Y(n6196) );
  OAI21X1 U12945 ( .A(n10938), .B(n10813), .C(n274), .Y(n6197) );
  OAI21X1 U12946 ( .A(n10940), .B(n10813), .C(n381), .Y(n6198) );
  OAI21X1 U12947 ( .A(n10942), .B(n10813), .C(n488), .Y(n6199) );
  OAI21X1 U12948 ( .A(n10944), .B(n10813), .C(n1556), .Y(n6200) );
  OAI21X1 U12949 ( .A(n10946), .B(n10813), .C(n1715), .Y(n6201) );
  OAI21X1 U12950 ( .A(n10948), .B(n10813), .C(n1873), .Y(n6202) );
  OAI21X1 U12951 ( .A(n10950), .B(n10813), .C(n2030), .Y(n6203) );
  OAI21X1 U12952 ( .A(n10954), .B(n10813), .C(n1055), .Y(n6204) );
  NAND3X1 U12953 ( .A(n10965), .B(n10964), .C(n11112), .Y(n13096) );
  OAI21X1 U12954 ( .A(n1520), .B(n1679), .C(n10956), .Y(n12700) );
  OAI21X1 U12955 ( .A(n10826), .B(n10815), .C(n2029), .Y(n6205) );
  OAI21X1 U12956 ( .A(n10828), .B(n10815), .C(n1872), .Y(n6206) );
  OAI21X1 U12957 ( .A(n10830), .B(n10815), .C(n1714), .Y(n6207) );
  OAI21X1 U12958 ( .A(n10832), .B(n10815), .C(n1555), .Y(n6208) );
  OAI21X1 U12959 ( .A(n10834), .B(n10815), .C(n1430), .Y(n6209) );
  OAI21X1 U12960 ( .A(n10836), .B(n10815), .C(n1304), .Y(n6210) );
  OAI21X1 U12961 ( .A(n10838), .B(n10815), .C(n1179), .Y(n6211) );
  OAI21X1 U12962 ( .A(n10840), .B(n10815), .C(n1054), .Y(n6212) );
  OAI21X1 U12963 ( .A(n10842), .B(n10815), .C(n931), .Y(n6213) );
  OAI21X1 U12964 ( .A(n10844), .B(n10815), .C(n819), .Y(n6214) );
  OAI21X1 U12965 ( .A(n10846), .B(n10815), .C(n707), .Y(n6215) );
  OAI21X1 U12966 ( .A(n10848), .B(n10815), .C(n595), .Y(n6216) );
  OAI21X1 U12967 ( .A(n10850), .B(n10815), .C(n2028), .Y(n6217) );
  OAI21X1 U12968 ( .A(n10852), .B(n10815), .C(n1871), .Y(n6218) );
  OAI21X1 U12969 ( .A(n10854), .B(n10815), .C(n1713), .Y(n6219) );
  OAI21X1 U12970 ( .A(n10856), .B(n10815), .C(n1554), .Y(n6220) );
  OAI21X1 U12971 ( .A(n10858), .B(n10815), .C(n1429), .Y(n6221) );
  OAI21X1 U12972 ( .A(n10860), .B(n10815), .C(n1303), .Y(n6222) );
  OAI21X1 U12973 ( .A(n10862), .B(n10815), .C(n1178), .Y(n6223) );
  OAI21X1 U12974 ( .A(n10864), .B(n10815), .C(n1053), .Y(n6224) );
  OAI21X1 U12975 ( .A(n10866), .B(n10815), .C(n930), .Y(n6225) );
  OAI21X1 U12976 ( .A(n10868), .B(n10815), .C(n818), .Y(n6226) );
  OAI21X1 U12977 ( .A(n10870), .B(n10815), .C(n706), .Y(n6227) );
  OAI21X1 U12978 ( .A(n10872), .B(n10815), .C(n594), .Y(n6228) );
  OAI21X1 U12979 ( .A(n10874), .B(n10815), .C(n487), .Y(n6229) );
  OAI21X1 U12980 ( .A(n10876), .B(n10815), .C(n2027), .Y(n6230) );
  OAI21X1 U12981 ( .A(n10878), .B(n10815), .C(n1870), .Y(n6231) );
  OAI21X1 U12982 ( .A(n10880), .B(n10815), .C(n1712), .Y(n6232) );
  OAI21X1 U12983 ( .A(n10882), .B(n10815), .C(n1553), .Y(n6233) );
  OAI21X1 U12984 ( .A(n10884), .B(n10815), .C(n1428), .Y(n6234) );
  OAI21X1 U12985 ( .A(n10886), .B(n10815), .C(n1302), .Y(n6235) );
  OAI21X1 U12986 ( .A(n10888), .B(n10815), .C(n1177), .Y(n6236) );
  OAI21X1 U12987 ( .A(n10890), .B(n10815), .C(n1052), .Y(n6237) );
  OAI21X1 U12988 ( .A(n10892), .B(n10815), .C(n929), .Y(n6238) );
  OAI21X1 U12989 ( .A(n10894), .B(n10815), .C(n817), .Y(n6239) );
  OAI21X1 U12990 ( .A(n10896), .B(n10815), .C(n705), .Y(n6240) );
  OAI21X1 U12991 ( .A(n10898), .B(n10815), .C(n593), .Y(n6241) );
  OAI21X1 U12992 ( .A(n10900), .B(n10815), .C(n486), .Y(n6242) );
  OAI21X1 U12993 ( .A(n10902), .B(n10815), .C(n2026), .Y(n6243) );
  OAI21X1 U12994 ( .A(n10904), .B(n10815), .C(n1869), .Y(n6244) );
  OAI21X1 U12995 ( .A(n10906), .B(n10815), .C(n1711), .Y(n6245) );
  OAI21X1 U12996 ( .A(n10908), .B(n10815), .C(n1552), .Y(n6246) );
  OAI21X1 U12997 ( .A(n10910), .B(n10815), .C(n1427), .Y(n6247) );
  OAI21X1 U12998 ( .A(n10912), .B(n10815), .C(n1301), .Y(n6248) );
  OAI21X1 U12999 ( .A(n10914), .B(n10815), .C(n1176), .Y(n6249) );
  OAI21X1 U13000 ( .A(n10916), .B(n10815), .C(n1051), .Y(n6250) );
  OAI21X1 U13001 ( .A(n10918), .B(n10815), .C(n928), .Y(n6251) );
  OAI21X1 U13002 ( .A(n10920), .B(n10815), .C(n816), .Y(n6252) );
  OAI21X1 U13003 ( .A(n10922), .B(n10815), .C(n704), .Y(n6253) );
  OAI21X1 U13004 ( .A(n10924), .B(n10815), .C(n592), .Y(n6254) );
  OAI21X1 U13005 ( .A(n10926), .B(n10815), .C(n485), .Y(n6255) );
  OAI21X1 U13006 ( .A(n10928), .B(n10815), .C(n2025), .Y(n6256) );
  OAI21X1 U13007 ( .A(n10930), .B(n10815), .C(n1868), .Y(n6257) );
  OAI21X1 U13008 ( .A(n10932), .B(n10815), .C(n1710), .Y(n6258) );
  OAI21X1 U13009 ( .A(n10934), .B(n10815), .C(n1551), .Y(n6259) );
  OAI21X1 U13010 ( .A(n10936), .B(n10815), .C(n1426), .Y(n6260) );
  OAI21X1 U13011 ( .A(n10938), .B(n10815), .C(n1300), .Y(n6261) );
  OAI21X1 U13012 ( .A(n10940), .B(n10815), .C(n1175), .Y(n6262) );
  OAI21X1 U13013 ( .A(n10942), .B(n10815), .C(n1050), .Y(n6263) );
  OAI21X1 U13014 ( .A(n10944), .B(n10815), .C(n927), .Y(n6264) );
  OAI21X1 U13015 ( .A(n10946), .B(n10815), .C(n815), .Y(n6265) );
  OAI21X1 U13016 ( .A(n10948), .B(n10815), .C(n703), .Y(n6266) );
  OAI21X1 U13017 ( .A(n10950), .B(n10815), .C(n591), .Y(n6267) );
  OAI21X1 U13018 ( .A(n10954), .B(n10815), .C(n484), .Y(n6268) );
  OAI21X1 U13019 ( .A(n1395), .B(n1679), .C(n10956), .Y(n12766) );
  OAI21X1 U13020 ( .A(n10826), .B(n10817), .C(n1867), .Y(n6269) );
  OAI21X1 U13021 ( .A(n10828), .B(n10817), .C(n2024), .Y(n6270) );
  OAI21X1 U13022 ( .A(n10830), .B(n10817), .C(n1550), .Y(n6271) );
  OAI21X1 U13023 ( .A(n10832), .B(n10817), .C(n1709), .Y(n6272) );
  OAI21X1 U13024 ( .A(n10834), .B(n10817), .C(n1299), .Y(n6273) );
  OAI21X1 U13025 ( .A(n10836), .B(n10817), .C(n1425), .Y(n6274) );
  OAI21X1 U13026 ( .A(n10838), .B(n10817), .C(n1049), .Y(n6275) );
  OAI21X1 U13027 ( .A(n10840), .B(n10817), .C(n1174), .Y(n6276) );
  OAI21X1 U13028 ( .A(n10842), .B(n10817), .C(n814), .Y(n6277) );
  OAI21X1 U13029 ( .A(n10844), .B(n10817), .C(n926), .Y(n6278) );
  OAI21X1 U13030 ( .A(n10846), .B(n10817), .C(n590), .Y(n6279) );
  OAI21X1 U13031 ( .A(n10848), .B(n10817), .C(n702), .Y(n6280) );
  OAI21X1 U13032 ( .A(n10850), .B(n10817), .C(n1866), .Y(n6281) );
  OAI21X1 U13033 ( .A(n10852), .B(n10817), .C(n2023), .Y(n6282) );
  OAI21X1 U13034 ( .A(n10854), .B(n10817), .C(n1549), .Y(n6283) );
  OAI21X1 U13035 ( .A(n10856), .B(n10817), .C(n1708), .Y(n6284) );
  OAI21X1 U13036 ( .A(n10858), .B(n10817), .C(n1298), .Y(n6285) );
  OAI21X1 U13037 ( .A(n10860), .B(n10817), .C(n1424), .Y(n6286) );
  OAI21X1 U13038 ( .A(n10862), .B(n10817), .C(n1048), .Y(n6287) );
  OAI21X1 U13039 ( .A(n10864), .B(n10817), .C(n1173), .Y(n6288) );
  OAI21X1 U13040 ( .A(n10866), .B(n10817), .C(n813), .Y(n6289) );
  OAI21X1 U13041 ( .A(n10868), .B(n10817), .C(n925), .Y(n6290) );
  OAI21X1 U13042 ( .A(n10870), .B(n10817), .C(n589), .Y(n6291) );
  OAI21X1 U13043 ( .A(n10872), .B(n10817), .C(n701), .Y(n6292) );
  OAI21X1 U13044 ( .A(n10874), .B(n10817), .C(n380), .Y(n6293) );
  OAI21X1 U13045 ( .A(n10876), .B(n10817), .C(n1865), .Y(n6294) );
  OAI21X1 U13046 ( .A(n10878), .B(n10817), .C(n2022), .Y(n6295) );
  OAI21X1 U13047 ( .A(n10880), .B(n10817), .C(n1548), .Y(n6296) );
  OAI21X1 U13048 ( .A(n10882), .B(n10817), .C(n1707), .Y(n6297) );
  OAI21X1 U13049 ( .A(n10884), .B(n10817), .C(n1297), .Y(n6298) );
  OAI21X1 U13050 ( .A(n10886), .B(n10817), .C(n1423), .Y(n6299) );
  OAI21X1 U13051 ( .A(n10888), .B(n10817), .C(n1047), .Y(n6300) );
  OAI21X1 U13052 ( .A(n10890), .B(n10817), .C(n1172), .Y(n6301) );
  OAI21X1 U13053 ( .A(n10892), .B(n10817), .C(n812), .Y(n6302) );
  OAI21X1 U13054 ( .A(n10894), .B(n10817), .C(n924), .Y(n6303) );
  OAI21X1 U13055 ( .A(n10896), .B(n10817), .C(n588), .Y(n6304) );
  OAI21X1 U13056 ( .A(n10898), .B(n10817), .C(n700), .Y(n6305) );
  OAI21X1 U13057 ( .A(n10900), .B(n10817), .C(n379), .Y(n6306) );
  OAI21X1 U13058 ( .A(n10902), .B(n10817), .C(n1864), .Y(n6307) );
  OAI21X1 U13059 ( .A(n10904), .B(n10817), .C(n2021), .Y(n6308) );
  OAI21X1 U13060 ( .A(n10906), .B(n10817), .C(n1547), .Y(n6309) );
  OAI21X1 U13061 ( .A(n10908), .B(n10817), .C(n1706), .Y(n6310) );
  OAI21X1 U13062 ( .A(n10910), .B(n10817), .C(n1296), .Y(n6311) );
  OAI21X1 U13063 ( .A(n10912), .B(n10817), .C(n1422), .Y(n6312) );
  OAI21X1 U13064 ( .A(n10914), .B(n10817), .C(n1046), .Y(n6313) );
  OAI21X1 U13065 ( .A(n10916), .B(n10817), .C(n1171), .Y(n6314) );
  OAI21X1 U13066 ( .A(n10918), .B(n10817), .C(n811), .Y(n6315) );
  OAI21X1 U13067 ( .A(n10920), .B(n10817), .C(n923), .Y(n6316) );
  OAI21X1 U13068 ( .A(n10922), .B(n10817), .C(n587), .Y(n6317) );
  OAI21X1 U13069 ( .A(n10924), .B(n10817), .C(n699), .Y(n6318) );
  OAI21X1 U13070 ( .A(n10926), .B(n10817), .C(n378), .Y(n6319) );
  OAI21X1 U13071 ( .A(n10928), .B(n10817), .C(n1863), .Y(n6320) );
  OAI21X1 U13072 ( .A(n10930), .B(n10817), .C(n2020), .Y(n6321) );
  OAI21X1 U13073 ( .A(n10932), .B(n10817), .C(n1546), .Y(n6322) );
  OAI21X1 U13074 ( .A(n10934), .B(n10817), .C(n1705), .Y(n6323) );
  OAI21X1 U13075 ( .A(n10936), .B(n10817), .C(n1295), .Y(n6324) );
  OAI21X1 U13076 ( .A(n10938), .B(n10817), .C(n1421), .Y(n6325) );
  OAI21X1 U13077 ( .A(n10940), .B(n10817), .C(n1045), .Y(n6326) );
  OAI21X1 U13078 ( .A(n10942), .B(n10817), .C(n1170), .Y(n6327) );
  OAI21X1 U13079 ( .A(n10944), .B(n10817), .C(n810), .Y(n6328) );
  OAI21X1 U13080 ( .A(n10946), .B(n10817), .C(n922), .Y(n6329) );
  OAI21X1 U13081 ( .A(n10948), .B(n10817), .C(n586), .Y(n6330) );
  OAI21X1 U13082 ( .A(n10950), .B(n10817), .C(n698), .Y(n6331) );
  OAI21X1 U13083 ( .A(n10954), .B(n10817), .C(n377), .Y(n6332) );
  OAI21X1 U13084 ( .A(n1269), .B(n1679), .C(n10956), .Y(n12832) );
  OAI21X1 U13085 ( .A(n10826), .B(n10819), .C(n1704), .Y(n6333) );
  OAI21X1 U13086 ( .A(n10828), .B(n10819), .C(n1545), .Y(n6334) );
  OAI21X1 U13087 ( .A(n10830), .B(n10819), .C(n2019), .Y(n6335) );
  OAI21X1 U13088 ( .A(n10832), .B(n10819), .C(n1862), .Y(n6336) );
  OAI21X1 U13089 ( .A(n10834), .B(n10819), .C(n1169), .Y(n6337) );
  OAI21X1 U13090 ( .A(n10836), .B(n10819), .C(n1044), .Y(n6338) );
  OAI21X1 U13091 ( .A(n10838), .B(n10819), .C(n1420), .Y(n6339) );
  OAI21X1 U13092 ( .A(n10840), .B(n10819), .C(n1294), .Y(n6340) );
  OAI21X1 U13093 ( .A(n10842), .B(n10819), .C(n697), .Y(n6341) );
  OAI21X1 U13094 ( .A(n10844), .B(n10819), .C(n585), .Y(n6342) );
  OAI21X1 U13095 ( .A(n10846), .B(n10819), .C(n921), .Y(n6343) );
  OAI21X1 U13096 ( .A(n10848), .B(n10819), .C(n809), .Y(n6344) );
  OAI21X1 U13097 ( .A(n10850), .B(n10819), .C(n1703), .Y(n6345) );
  OAI21X1 U13098 ( .A(n10852), .B(n10819), .C(n1544), .Y(n6346) );
  OAI21X1 U13099 ( .A(n10854), .B(n10819), .C(n2018), .Y(n6347) );
  OAI21X1 U13100 ( .A(n10856), .B(n10819), .C(n1861), .Y(n6348) );
  OAI21X1 U13101 ( .A(n10858), .B(n10819), .C(n1168), .Y(n6349) );
  OAI21X1 U13102 ( .A(n10860), .B(n10819), .C(n1043), .Y(n6350) );
  OAI21X1 U13103 ( .A(n10862), .B(n10819), .C(n1419), .Y(n6351) );
  OAI21X1 U13104 ( .A(n10864), .B(n10819), .C(n1293), .Y(n6352) );
  OAI21X1 U13105 ( .A(n10866), .B(n10819), .C(n696), .Y(n6353) );
  OAI21X1 U13106 ( .A(n10868), .B(n10819), .C(n584), .Y(n6354) );
  OAI21X1 U13107 ( .A(n10870), .B(n10819), .C(n920), .Y(n6355) );
  OAI21X1 U13108 ( .A(n10872), .B(n10819), .C(n808), .Y(n6356) );
  OAI21X1 U13109 ( .A(n10874), .B(n10819), .C(n273), .Y(n6357) );
  OAI21X1 U13110 ( .A(n10876), .B(n10819), .C(n1702), .Y(n6358) );
  OAI21X1 U13111 ( .A(n10878), .B(n10819), .C(n1543), .Y(n6359) );
  OAI21X1 U13112 ( .A(n10880), .B(n10819), .C(n2017), .Y(n6360) );
  OAI21X1 U13113 ( .A(n10882), .B(n10819), .C(n1860), .Y(n6361) );
  OAI21X1 U13114 ( .A(n10884), .B(n10819), .C(n1167), .Y(n6362) );
  OAI21X1 U13115 ( .A(n10886), .B(n10819), .C(n1042), .Y(n6363) );
  OAI21X1 U13116 ( .A(n10888), .B(n10819), .C(n1418), .Y(n6364) );
  OAI21X1 U13117 ( .A(n10890), .B(n10819), .C(n1292), .Y(n6365) );
  OAI21X1 U13118 ( .A(n10892), .B(n10819), .C(n695), .Y(n6366) );
  OAI21X1 U13119 ( .A(n10894), .B(n10819), .C(n583), .Y(n6367) );
  OAI21X1 U13120 ( .A(n10896), .B(n10819), .C(n919), .Y(n6368) );
  OAI21X1 U13121 ( .A(n10898), .B(n10819), .C(n807), .Y(n6369) );
  OAI21X1 U13122 ( .A(n10900), .B(n10819), .C(n272), .Y(n6370) );
  OAI21X1 U13123 ( .A(n10902), .B(n10819), .C(n1701), .Y(n6371) );
  OAI21X1 U13124 ( .A(n10904), .B(n10819), .C(n1542), .Y(n6372) );
  OAI21X1 U13125 ( .A(n10906), .B(n10819), .C(n2016), .Y(n6373) );
  OAI21X1 U13126 ( .A(n10908), .B(n10819), .C(n1859), .Y(n6374) );
  OAI21X1 U13127 ( .A(n10910), .B(n10819), .C(n1166), .Y(n6375) );
  OAI21X1 U13128 ( .A(n10912), .B(n10819), .C(n1041), .Y(n6376) );
  OAI21X1 U13129 ( .A(n10914), .B(n10819), .C(n1417), .Y(n6377) );
  OAI21X1 U13130 ( .A(n10916), .B(n10819), .C(n1291), .Y(n6378) );
  OAI21X1 U13131 ( .A(n10918), .B(n10819), .C(n694), .Y(n6379) );
  OAI21X1 U13132 ( .A(n10920), .B(n10819), .C(n582), .Y(n6380) );
  OAI21X1 U13133 ( .A(n10922), .B(n10819), .C(n918), .Y(n6381) );
  OAI21X1 U13134 ( .A(n10924), .B(n10819), .C(n806), .Y(n6382) );
  OAI21X1 U13135 ( .A(n10926), .B(n10819), .C(n271), .Y(n6383) );
  OAI21X1 U13136 ( .A(n10928), .B(n10819), .C(n1700), .Y(n6384) );
  OAI21X1 U13137 ( .A(n10930), .B(n10819), .C(n1541), .Y(n6385) );
  OAI21X1 U13138 ( .A(n10932), .B(n10819), .C(n2015), .Y(n6386) );
  OAI21X1 U13139 ( .A(n10934), .B(n10819), .C(n1858), .Y(n6387) );
  OAI21X1 U13140 ( .A(n10936), .B(n10819), .C(n1165), .Y(n6388) );
  OAI21X1 U13141 ( .A(n10938), .B(n10819), .C(n1040), .Y(n6389) );
  OAI21X1 U13142 ( .A(n10940), .B(n10819), .C(n1416), .Y(n6390) );
  OAI21X1 U13143 ( .A(n10942), .B(n10819), .C(n1290), .Y(n6391) );
  OAI21X1 U13144 ( .A(n10944), .B(n10819), .C(n693), .Y(n6392) );
  OAI21X1 U13145 ( .A(n10946), .B(n10819), .C(n581), .Y(n6393) );
  OAI21X1 U13146 ( .A(n10948), .B(n10819), .C(n917), .Y(n6394) );
  OAI21X1 U13147 ( .A(n10950), .B(n10819), .C(n805), .Y(n6395) );
  OAI21X1 U13148 ( .A(n10954), .B(n10819), .C(n270), .Y(n6396) );
  OAI21X1 U13149 ( .A(n1144), .B(n1679), .C(n10956), .Y(n12898) );
  OAI21X1 U13150 ( .A(n10826), .B(n10821), .C(n1540), .Y(n6397) );
  OAI21X1 U13151 ( .A(n10828), .B(n10821), .C(n1699), .Y(n6398) );
  OAI21X1 U13152 ( .A(n10830), .B(n10821), .C(n1857), .Y(n6399) );
  OAI21X1 U13153 ( .A(n10832), .B(n10821), .C(n2014), .Y(n6400) );
  OAI21X1 U13154 ( .A(n10834), .B(n10821), .C(n1039), .Y(n6401) );
  OAI21X1 U13155 ( .A(n10836), .B(n10821), .C(n1164), .Y(n6402) );
  OAI21X1 U13156 ( .A(n10838), .B(n10821), .C(n1289), .Y(n6403) );
  OAI21X1 U13157 ( .A(n10840), .B(n10821), .C(n1415), .Y(n6404) );
  OAI21X1 U13158 ( .A(n10842), .B(n10821), .C(n580), .Y(n6405) );
  OAI21X1 U13159 ( .A(n10844), .B(n10821), .C(n692), .Y(n6406) );
  OAI21X1 U13160 ( .A(n10846), .B(n10821), .C(n804), .Y(n6407) );
  OAI21X1 U13161 ( .A(n10848), .B(n10821), .C(n916), .Y(n6408) );
  OAI21X1 U13162 ( .A(n10850), .B(n10821), .C(n1539), .Y(n6409) );
  OAI21X1 U13163 ( .A(n10852), .B(n10821), .C(n1698), .Y(n6410) );
  OAI21X1 U13164 ( .A(n10854), .B(n10821), .C(n1856), .Y(n6411) );
  OAI21X1 U13165 ( .A(n10856), .B(n10821), .C(n2013), .Y(n6412) );
  OAI21X1 U13166 ( .A(n10858), .B(n10821), .C(n1038), .Y(n6413) );
  OAI21X1 U13167 ( .A(n10860), .B(n10821), .C(n1163), .Y(n6414) );
  OAI21X1 U13168 ( .A(n10862), .B(n10821), .C(n1288), .Y(n6415) );
  OAI21X1 U13169 ( .A(n10864), .B(n10821), .C(n1414), .Y(n6416) );
  OAI21X1 U13170 ( .A(n10866), .B(n10821), .C(n579), .Y(n6417) );
  OAI21X1 U13171 ( .A(n10868), .B(n10821), .C(n691), .Y(n6418) );
  OAI21X1 U13172 ( .A(n10870), .B(n10821), .C(n803), .Y(n6419) );
  OAI21X1 U13173 ( .A(n10872), .B(n10821), .C(n915), .Y(n6420) );
  OAI21X1 U13174 ( .A(n10874), .B(n10821), .C(n38), .Y(n6421) );
  OAI21X1 U13175 ( .A(n10876), .B(n10821), .C(n1538), .Y(n6422) );
  OAI21X1 U13176 ( .A(n10878), .B(n10821), .C(n1697), .Y(n6423) );
  OAI21X1 U13177 ( .A(n10880), .B(n10821), .C(n1855), .Y(n6424) );
  OAI21X1 U13178 ( .A(n10882), .B(n10821), .C(n2012), .Y(n6425) );
  OAI21X1 U13179 ( .A(n10884), .B(n10821), .C(n1037), .Y(n6426) );
  OAI21X1 U13180 ( .A(n10886), .B(n10821), .C(n1162), .Y(n6427) );
  OAI21X1 U13181 ( .A(n10888), .B(n10821), .C(n1287), .Y(n6428) );
  OAI21X1 U13182 ( .A(n10890), .B(n10821), .C(n1413), .Y(n6429) );
  OAI21X1 U13183 ( .A(n10892), .B(n10821), .C(n578), .Y(n6430) );
  OAI21X1 U13184 ( .A(n10894), .B(n10821), .C(n690), .Y(n6431) );
  OAI21X1 U13185 ( .A(n10896), .B(n10821), .C(n802), .Y(n6432) );
  OAI21X1 U13186 ( .A(n10898), .B(n10821), .C(n914), .Y(n6433) );
  OAI21X1 U13187 ( .A(n10900), .B(n10821), .C(n37), .Y(n6434) );
  OAI21X1 U13188 ( .A(n10902), .B(n10821), .C(n1537), .Y(n6435) );
  OAI21X1 U13189 ( .A(n10904), .B(n10821), .C(n1696), .Y(n6436) );
  OAI21X1 U13190 ( .A(n10906), .B(n10821), .C(n1854), .Y(n6437) );
  OAI21X1 U13191 ( .A(n10908), .B(n10821), .C(n2011), .Y(n6438) );
  OAI21X1 U13192 ( .A(n10910), .B(n10821), .C(n1036), .Y(n6439) );
  OAI21X1 U13193 ( .A(n10912), .B(n10821), .C(n1161), .Y(n6440) );
  OAI21X1 U13194 ( .A(n10914), .B(n10821), .C(n1286), .Y(n6441) );
  OAI21X1 U13195 ( .A(n10916), .B(n10821), .C(n1412), .Y(n6442) );
  OAI21X1 U13196 ( .A(n10918), .B(n10821), .C(n577), .Y(n6443) );
  OAI21X1 U13197 ( .A(n10920), .B(n10821), .C(n689), .Y(n6444) );
  OAI21X1 U13198 ( .A(n10922), .B(n10821), .C(n801), .Y(n6445) );
  OAI21X1 U13199 ( .A(n10924), .B(n10821), .C(n913), .Y(n6446) );
  OAI21X1 U13200 ( .A(n10926), .B(n10821), .C(n36), .Y(n6447) );
  OAI21X1 U13201 ( .A(n10928), .B(n10821), .C(n1536), .Y(n6448) );
  OAI21X1 U13202 ( .A(n10930), .B(n10821), .C(n1695), .Y(n6449) );
  OAI21X1 U13203 ( .A(n10932), .B(n10821), .C(n1853), .Y(n6450) );
  OAI21X1 U13204 ( .A(n10934), .B(n10821), .C(n2010), .Y(n6451) );
  OAI21X1 U13205 ( .A(n10936), .B(n10821), .C(n1035), .Y(n6452) );
  OAI21X1 U13206 ( .A(n10938), .B(n10821), .C(n1160), .Y(n6453) );
  OAI21X1 U13207 ( .A(n10940), .B(n10821), .C(n1285), .Y(n6454) );
  OAI21X1 U13208 ( .A(n10942), .B(n10821), .C(n1411), .Y(n6455) );
  OAI21X1 U13209 ( .A(n10944), .B(n10821), .C(n576), .Y(n6456) );
  OAI21X1 U13210 ( .A(n10946), .B(n10821), .C(n688), .Y(n6457) );
  OAI21X1 U13211 ( .A(n10948), .B(n10821), .C(n800), .Y(n6458) );
  OAI21X1 U13212 ( .A(n10950), .B(n10821), .C(n912), .Y(n6459) );
  OAI21X1 U13213 ( .A(n10954), .B(n10821), .C(n35), .Y(n6460) );
  OAI21X1 U13214 ( .A(n1143), .B(n1679), .C(n10956), .Y(n12964) );
  OAI21X1 U13215 ( .A(n10826), .B(n10823), .C(n1410), .Y(n6461) );
  OAI21X1 U13216 ( .A(n10828), .B(n10823), .C(n1284), .Y(n6462) );
  OAI21X1 U13217 ( .A(n10830), .B(n10823), .C(n1159), .Y(n6463) );
  OAI21X1 U13218 ( .A(n10832), .B(n10823), .C(n1034), .Y(n6464) );
  OAI21X1 U13219 ( .A(n10834), .B(n10823), .C(n2009), .Y(n6465) );
  OAI21X1 U13220 ( .A(n10836), .B(n10823), .C(n1852), .Y(n6466) );
  OAI21X1 U13221 ( .A(n10838), .B(n10823), .C(n1694), .Y(n6467) );
  OAI21X1 U13222 ( .A(n10840), .B(n10823), .C(n1535), .Y(n6468) );
  OAI21X1 U13223 ( .A(n10842), .B(n10823), .C(n483), .Y(n6469) );
  OAI21X1 U13224 ( .A(n10844), .B(n10823), .C(n376), .Y(n6470) );
  OAI21X1 U13225 ( .A(n10846), .B(n10823), .C(n269), .Y(n6471) );
  OAI21X1 U13226 ( .A(n10848), .B(n10823), .C(n34), .Y(n6472) );
  OAI21X1 U13227 ( .A(n10850), .B(n10823), .C(n1409), .Y(n6473) );
  OAI21X1 U13228 ( .A(n10852), .B(n10823), .C(n1283), .Y(n6474) );
  OAI21X1 U13229 ( .A(n10854), .B(n10823), .C(n1158), .Y(n6475) );
  OAI21X1 U13230 ( .A(n10856), .B(n10823), .C(n1033), .Y(n6476) );
  OAI21X1 U13231 ( .A(n10858), .B(n10823), .C(n2008), .Y(n6477) );
  OAI21X1 U13232 ( .A(n10860), .B(n10823), .C(n1851), .Y(n6478) );
  OAI21X1 U13233 ( .A(n10862), .B(n10823), .C(n1693), .Y(n6479) );
  OAI21X1 U13234 ( .A(n10864), .B(n10823), .C(n1534), .Y(n6480) );
  OAI21X1 U13235 ( .A(n10866), .B(n10823), .C(n482), .Y(n6481) );
  OAI21X1 U13236 ( .A(n10868), .B(n10823), .C(n375), .Y(n6482) );
  OAI21X1 U13237 ( .A(n10870), .B(n10823), .C(n268), .Y(n6483) );
  OAI21X1 U13238 ( .A(n10872), .B(n10823), .C(n18), .Y(n6484) );
  OAI21X1 U13239 ( .A(n10874), .B(n10823), .C(n911), .Y(n6485) );
  OAI21X1 U13240 ( .A(n10876), .B(n10823), .C(n1408), .Y(n6486) );
  OAI21X1 U13241 ( .A(n10878), .B(n10823), .C(n1282), .Y(n6487) );
  OAI21X1 U13242 ( .A(n10880), .B(n10823), .C(n1157), .Y(n6488) );
  OAI21X1 U13243 ( .A(n10882), .B(n10823), .C(n1032), .Y(n6489) );
  OAI21X1 U13244 ( .A(n10884), .B(n10823), .C(n2007), .Y(n6490) );
  OAI21X1 U13245 ( .A(n10886), .B(n10823), .C(n1850), .Y(n6491) );
  OAI21X1 U13246 ( .A(n10888), .B(n10823), .C(n1692), .Y(n6492) );
  OAI21X1 U13247 ( .A(n10890), .B(n10823), .C(n1533), .Y(n6493) );
  OAI21X1 U13248 ( .A(n10892), .B(n10823), .C(n481), .Y(n6494) );
  OAI21X1 U13249 ( .A(n10894), .B(n10823), .C(n374), .Y(n6495) );
  OAI21X1 U13250 ( .A(n10896), .B(n10823), .C(n267), .Y(n6496) );
  OAI21X1 U13251 ( .A(n10898), .B(n10823), .C(n17), .Y(n6497) );
  OAI21X1 U13252 ( .A(n10900), .B(n10823), .C(n910), .Y(n6498) );
  OAI21X1 U13253 ( .A(n10902), .B(n10823), .C(n1407), .Y(n6499) );
  OAI21X1 U13254 ( .A(n10904), .B(n10823), .C(n1281), .Y(n6500) );
  OAI21X1 U13255 ( .A(n10906), .B(n10823), .C(n1156), .Y(n6501) );
  OAI21X1 U13256 ( .A(n10908), .B(n10823), .C(n1031), .Y(n6502) );
  OAI21X1 U13257 ( .A(n10910), .B(n10823), .C(n2006), .Y(n6503) );
  OAI21X1 U13258 ( .A(n10912), .B(n10823), .C(n1849), .Y(n6504) );
  OAI21X1 U13259 ( .A(n10914), .B(n10823), .C(n1691), .Y(n6505) );
  OAI21X1 U13260 ( .A(n10916), .B(n10823), .C(n1532), .Y(n6506) );
  OAI21X1 U13261 ( .A(n10918), .B(n10823), .C(n480), .Y(n6507) );
  OAI21X1 U13262 ( .A(n10920), .B(n10823), .C(n373), .Y(n6508) );
  OAI21X1 U13263 ( .A(n10922), .B(n10823), .C(n266), .Y(n6509) );
  OAI21X1 U13264 ( .A(n10924), .B(n10823), .C(n16), .Y(n6510) );
  OAI21X1 U13265 ( .A(n10926), .B(n10823), .C(n909), .Y(n6511) );
  OAI21X1 U13266 ( .A(n10928), .B(n10823), .C(n1406), .Y(n6512) );
  OAI21X1 U13267 ( .A(n10930), .B(n10823), .C(n1280), .Y(n6513) );
  OAI21X1 U13268 ( .A(n10932), .B(n10823), .C(n1155), .Y(n6514) );
  OAI21X1 U13269 ( .A(n10934), .B(n10823), .C(n1030), .Y(n6515) );
  OAI21X1 U13270 ( .A(n10936), .B(n10823), .C(n2005), .Y(n6516) );
  OAI21X1 U13271 ( .A(n10938), .B(n10823), .C(n1848), .Y(n6517) );
  OAI21X1 U13272 ( .A(n10940), .B(n10823), .C(n1690), .Y(n6518) );
  OAI21X1 U13273 ( .A(n10942), .B(n10823), .C(n1531), .Y(n6519) );
  OAI21X1 U13274 ( .A(n10944), .B(n10823), .C(n479), .Y(n6520) );
  OAI21X1 U13275 ( .A(n10946), .B(n10823), .C(n372), .Y(n6521) );
  OAI21X1 U13276 ( .A(n10948), .B(n10823), .C(n265), .Y(n6522) );
  OAI21X1 U13277 ( .A(n10950), .B(n10823), .C(n15), .Y(n6523) );
  OAI21X1 U13278 ( .A(n10954), .B(n10823), .C(n908), .Y(n6524) );
  OAI21X1 U13279 ( .A(n1268), .B(n1679), .C(n10956), .Y(n13030) );
  OAI21X1 U13280 ( .A(n10826), .B(n10825), .C(n1279), .Y(n6525) );
  OAI21X1 U13281 ( .A(n10828), .B(n10825), .C(n1405), .Y(n6526) );
  OAI21X1 U13282 ( .A(n10830), .B(n10825), .C(n1029), .Y(n6527) );
  OAI21X1 U13283 ( .A(n10832), .B(n10825), .C(n1154), .Y(n6528) );
  OAI21X1 U13284 ( .A(n10834), .B(n10825), .C(n1847), .Y(n6529) );
  OAI21X1 U13285 ( .A(n10836), .B(n10825), .C(n2004), .Y(n6530) );
  OAI21X1 U13286 ( .A(n10838), .B(n10825), .C(n1530), .Y(n6531) );
  OAI21X1 U13287 ( .A(n10840), .B(n10825), .C(n1689), .Y(n6532) );
  OAI21X1 U13288 ( .A(n10842), .B(n10825), .C(n371), .Y(n6533) );
  OAI21X1 U13289 ( .A(n10844), .B(n10825), .C(n478), .Y(n6534) );
  OAI21X1 U13290 ( .A(n10846), .B(n10825), .C(n14), .Y(n6535) );
  OAI21X1 U13291 ( .A(n10848), .B(n10825), .C(n264), .Y(n6536) );
  OAI21X1 U13292 ( .A(n10850), .B(n10825), .C(n1278), .Y(n6537) );
  OAI21X1 U13293 ( .A(n10852), .B(n10825), .C(n1404), .Y(n6538) );
  OAI21X1 U13294 ( .A(n10854), .B(n10825), .C(n1028), .Y(n6539) );
  OAI21X1 U13295 ( .A(n10856), .B(n10825), .C(n1153), .Y(n6540) );
  OAI21X1 U13296 ( .A(n10858), .B(n10825), .C(n1846), .Y(n6541) );
  OAI21X1 U13297 ( .A(n10860), .B(n10825), .C(n2003), .Y(n6542) );
  OAI21X1 U13298 ( .A(n10862), .B(n10825), .C(n1529), .Y(n6543) );
  OAI21X1 U13299 ( .A(n10864), .B(n10825), .C(n1688), .Y(n6544) );
  OAI21X1 U13300 ( .A(n10866), .B(n10825), .C(n370), .Y(n6545) );
  OAI21X1 U13301 ( .A(n10868), .B(n10825), .C(n477), .Y(n6546) );
  OAI21X1 U13302 ( .A(n10870), .B(n10825), .C(n13), .Y(n6547) );
  OAI21X1 U13303 ( .A(n10872), .B(n10825), .C(n263), .Y(n6548) );
  OAI21X1 U13304 ( .A(n10874), .B(n10825), .C(n799), .Y(n6549) );
  OAI21X1 U13305 ( .A(n10876), .B(n10825), .C(n1277), .Y(n6550) );
  OAI21X1 U13306 ( .A(n10878), .B(n10825), .C(n1403), .Y(n6551) );
  OAI21X1 U13307 ( .A(n10880), .B(n10825), .C(n1027), .Y(n6552) );
  OAI21X1 U13308 ( .A(n10882), .B(n10825), .C(n1152), .Y(n6553) );
  OAI21X1 U13309 ( .A(n10884), .B(n10825), .C(n1845), .Y(n6554) );
  OAI21X1 U13310 ( .A(n10886), .B(n10825), .C(n2002), .Y(n6555) );
  OAI21X1 U13311 ( .A(n10888), .B(n10825), .C(n1528), .Y(n6556) );
  OAI21X1 U13312 ( .A(n10890), .B(n10825), .C(n1687), .Y(n6557) );
  OAI21X1 U13313 ( .A(n10892), .B(n10825), .C(n369), .Y(n6558) );
  OAI21X1 U13314 ( .A(n10894), .B(n10825), .C(n476), .Y(n6559) );
  OAI21X1 U13315 ( .A(n10896), .B(n10825), .C(n12), .Y(n6560) );
  OAI21X1 U13316 ( .A(n10898), .B(n10825), .C(n262), .Y(n6561) );
  OAI21X1 U13317 ( .A(n10900), .B(n10825), .C(n798), .Y(n6562) );
  OAI21X1 U13318 ( .A(n10902), .B(n10825), .C(n1276), .Y(n6563) );
  OAI21X1 U13319 ( .A(n10904), .B(n10825), .C(n1402), .Y(n6564) );
  OAI21X1 U13320 ( .A(n10906), .B(n10825), .C(n1026), .Y(n6565) );
  OAI21X1 U13321 ( .A(n10908), .B(n10825), .C(n1151), .Y(n6566) );
  OAI21X1 U13322 ( .A(n10910), .B(n10825), .C(n1844), .Y(n6567) );
  OAI21X1 U13323 ( .A(n10912), .B(n10825), .C(n2001), .Y(n6568) );
  OAI21X1 U13324 ( .A(n10914), .B(n10825), .C(n1527), .Y(n6569) );
  OAI21X1 U13325 ( .A(n10916), .B(n10825), .C(n1686), .Y(n6570) );
  OAI21X1 U13326 ( .A(n10918), .B(n10825), .C(n368), .Y(n6571) );
  OAI21X1 U13327 ( .A(n10920), .B(n10825), .C(n475), .Y(n6572) );
  OAI21X1 U13328 ( .A(n10922), .B(n10825), .C(n11), .Y(n6573) );
  OAI21X1 U13329 ( .A(n10924), .B(n10825), .C(n261), .Y(n6574) );
  OAI21X1 U13330 ( .A(n10926), .B(n10825), .C(n797), .Y(n6575) );
  OAI21X1 U13331 ( .A(n10928), .B(n10825), .C(n1275), .Y(n6576) );
  OAI21X1 U13332 ( .A(n10930), .B(n10825), .C(n1401), .Y(n6577) );
  OAI21X1 U13333 ( .A(n10932), .B(n10825), .C(n1025), .Y(n6578) );
  OAI21X1 U13334 ( .A(n10934), .B(n10825), .C(n1150), .Y(n6579) );
  OAI21X1 U13335 ( .A(n10936), .B(n10825), .C(n1843), .Y(n6580) );
  OAI21X1 U13336 ( .A(n10938), .B(n10825), .C(n2000), .Y(n6581) );
  OAI21X1 U13337 ( .A(n10940), .B(n10825), .C(n1526), .Y(n6582) );
  OAI21X1 U13338 ( .A(n10942), .B(n10825), .C(n1685), .Y(n6583) );
  OAI21X1 U13339 ( .A(n10944), .B(n10825), .C(n367), .Y(n6584) );
  OAI21X1 U13340 ( .A(n10946), .B(n10825), .C(n474), .Y(n6585) );
  OAI21X1 U13341 ( .A(n10948), .B(n10825), .C(n10), .Y(n6586) );
  OAI21X1 U13342 ( .A(n10950), .B(n10825), .C(n260), .Y(n6587) );
  OAI21X1 U13343 ( .A(n10954), .B(n10825), .C(n796), .Y(n6588) );
  OAI21X1 U13344 ( .A(n1394), .B(n1679), .C(n10956), .Y(n13097) );
  OAI21X1 U13345 ( .A(n10826), .B(n10953), .C(n1149), .Y(n6589) );
  OAI21X1 U13346 ( .A(n10828), .B(n10953), .C(n1024), .Y(n6590) );
  OAI21X1 U13347 ( .A(n10830), .B(n10953), .C(n1400), .Y(n6591) );
  OAI21X1 U13348 ( .A(n10832), .B(n10953), .C(n1274), .Y(n6592) );
  OAI21X1 U13349 ( .A(n10834), .B(n10953), .C(n1684), .Y(n6593) );
  OAI21X1 U13350 ( .A(n10836), .B(n10953), .C(n1525), .Y(n6594) );
  OAI21X1 U13351 ( .A(n10838), .B(n10953), .C(n1999), .Y(n6595) );
  OAI21X1 U13352 ( .A(n10840), .B(n10953), .C(n1842), .Y(n6596) );
  OAI21X1 U13353 ( .A(n10842), .B(n10953), .C(n259), .Y(n6597) );
  OAI21X1 U13354 ( .A(n10844), .B(n10953), .C(n9), .Y(n6598) );
  OAI21X1 U13355 ( .A(n10846), .B(n10953), .C(n473), .Y(n6599) );
  OAI21X1 U13356 ( .A(n10848), .B(n10953), .C(n366), .Y(n6600) );
  OAI21X1 U13357 ( .A(n10850), .B(n10953), .C(n1148), .Y(n6601) );
  OAI21X1 U13358 ( .A(n10852), .B(n10953), .C(n1023), .Y(n6602) );
  OAI21X1 U13359 ( .A(n10854), .B(n10953), .C(n1399), .Y(n6603) );
  OAI21X1 U13360 ( .A(n10856), .B(n10953), .C(n1273), .Y(n6604) );
  OAI21X1 U13361 ( .A(n10858), .B(n10953), .C(n1683), .Y(n6605) );
  OAI21X1 U13362 ( .A(n10860), .B(n10953), .C(n1524), .Y(n6606) );
  OAI21X1 U13363 ( .A(n10862), .B(n10953), .C(n1998), .Y(n6607) );
  OAI21X1 U13364 ( .A(n10864), .B(n10953), .C(n1841), .Y(n6608) );
  OAI21X1 U13365 ( .A(n10866), .B(n10953), .C(n258), .Y(n6609) );
  OAI21X1 U13366 ( .A(n10868), .B(n10953), .C(n8), .Y(n6610) );
  OAI21X1 U13367 ( .A(n10870), .B(n10953), .C(n472), .Y(n6611) );
  OAI21X1 U13368 ( .A(n10872), .B(n10953), .C(n365), .Y(n6612) );
  OAI21X1 U13369 ( .A(n10874), .B(n10953), .C(n687), .Y(n6613) );
  OAI21X1 U13370 ( .A(n10876), .B(n10953), .C(n1147), .Y(n6614) );
  OAI21X1 U13371 ( .A(n10878), .B(n10953), .C(n1022), .Y(n6615) );
  OAI21X1 U13372 ( .A(n10880), .B(n10953), .C(n1398), .Y(n6616) );
  OAI21X1 U13373 ( .A(n10882), .B(n10953), .C(n1272), .Y(n6617) );
  OAI21X1 U13374 ( .A(n10884), .B(n10953), .C(n1682), .Y(n6618) );
  OAI21X1 U13375 ( .A(n10886), .B(n10953), .C(n1523), .Y(n6619) );
  OAI21X1 U13376 ( .A(n10888), .B(n10953), .C(n1997), .Y(n6620) );
  OAI21X1 U13377 ( .A(n10890), .B(n10953), .C(n1840), .Y(n6621) );
  OAI21X1 U13378 ( .A(n10892), .B(n10953), .C(n257), .Y(n6622) );
  OAI21X1 U13379 ( .A(n10894), .B(n10953), .C(n7), .Y(n6623) );
  OAI21X1 U13380 ( .A(n10896), .B(n10953), .C(n471), .Y(n6624) );
  OAI21X1 U13381 ( .A(n10898), .B(n10953), .C(n364), .Y(n6625) );
  OAI21X1 U13382 ( .A(n10900), .B(n10953), .C(n686), .Y(n6626) );
  OAI21X1 U13383 ( .A(n10902), .B(n10953), .C(n1146), .Y(n6627) );
  OAI21X1 U13384 ( .A(n10904), .B(n10953), .C(n1021), .Y(n6628) );
  OAI21X1 U13385 ( .A(n10906), .B(n10953), .C(n1397), .Y(n6629) );
  OAI21X1 U13386 ( .A(n10908), .B(n10953), .C(n1271), .Y(n6630) );
  OAI21X1 U13387 ( .A(n10910), .B(n10953), .C(n1681), .Y(n6631) );
  OAI21X1 U13388 ( .A(n10912), .B(n10953), .C(n1522), .Y(n6632) );
  OAI21X1 U13389 ( .A(n10914), .B(n10953), .C(n1996), .Y(n6633) );
  OAI21X1 U13390 ( .A(n10916), .B(n10953), .C(n1839), .Y(n6634) );
  OAI21X1 U13391 ( .A(n10918), .B(n10953), .C(n256), .Y(n6635) );
  OAI21X1 U13392 ( .A(n10920), .B(n10953), .C(n6), .Y(n6636) );
  OAI21X1 U13393 ( .A(n10922), .B(n10953), .C(n470), .Y(n6637) );
  OAI21X1 U13394 ( .A(n10924), .B(n10953), .C(n363), .Y(n6638) );
  OAI21X1 U13395 ( .A(n10926), .B(n10953), .C(n685), .Y(n6639) );
  OAI21X1 U13396 ( .A(n10928), .B(n10953), .C(n1145), .Y(n6640) );
  OAI21X1 U13397 ( .A(n10930), .B(n10953), .C(n1020), .Y(n6641) );
  OAI21X1 U13398 ( .A(n10932), .B(n10953), .C(n1396), .Y(n6642) );
  OAI21X1 U13399 ( .A(n10934), .B(n10953), .C(n1270), .Y(n6643) );
  OAI21X1 U13400 ( .A(n10936), .B(n10953), .C(n1680), .Y(n6644) );
  OAI21X1 U13401 ( .A(n10938), .B(n10953), .C(n1521), .Y(n6645) );
  OAI21X1 U13402 ( .A(n10940), .B(n10953), .C(n1995), .Y(n6646) );
  OAI21X1 U13403 ( .A(n10942), .B(n10953), .C(n1838), .Y(n6647) );
  OAI21X1 U13404 ( .A(n10944), .B(n10953), .C(n255), .Y(n6648) );
  OAI21X1 U13405 ( .A(n10946), .B(n10953), .C(n5), .Y(n6649) );
  OAI21X1 U13406 ( .A(n10948), .B(n10953), .C(n469), .Y(n6650) );
  OAI21X1 U13407 ( .A(n10950), .B(n10953), .C(n362), .Y(n6651) );
  OAI21X1 U13408 ( .A(n10954), .B(n10953), .C(n684), .Y(n6652) );
endmodule


module alu_DW_mult_tc_1 ( a, b, product, ALU1ALU_MUL32_CLK );
  input [32:0] a;
  input [32:0] b;
  output [65:0] product;
  input ALU1ALU_MUL32_CLK;
  wire   n4, n9, n12, n16, n22, n24, n28, n34, n36, n40, n46, n48, n52, n58,
         n60, n64, n70, n72, n76, n82, n84, n88, n94, n96, n100, n106, n108,
         n112, n118, n120, n124, n127, n129, n227, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n294, n295, n296, n298, n300, n301, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n338,
         n339, n340, n341, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n360, n361, n362,
         n363, n365, n366, n367, n368, n369, n370, n371, n373, n376, n377,
         n379, n381, n382, n383, n384, n388, n390, n391, n393, n394, n395,
         n396, n397, n399, n400, n401, n403, n405, n406, n407, n408, n412,
         n414, n415, n417, n418, n419, n420, n421, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n434, n435, n436, n437, n439, n440,
         n441, n442, n443, n447, n449, n450, n451, n452, n456, n457, n458,
         n460, n462, n463, n465, n467, n468, n469, n470, n472, n475, n476,
         n477, n478, n480, n482, n483, n485, n487, n488, n489, n490, n492,
         n493, n494, n496, n498, n499, n501, n502, n503, n504, n506, n507,
         n508, n513, n514, n518, n519, n520, n523, n524, n525, n527, n528,
         n529, n530, n533, n534, n535, n536, n537, n541, n543, n544, n547,
         n548, n549, n550, n551, n552, n553, n556, n557, n558, n559, n560,
         n562, n563, n564, n565, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n593, n594, n595, n597,
         n599, n600, n602, n604, n605, n606, n607, n608, n609, n610, n612,
         n614, n615, n617, n619, n620, n621, n622, n624, n626, n627, n628,
         n629, n631, n634, n635, n636, n637, n639, n641, n642, n643, n644,
         n645, n646, n647, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n668, n669, n673,
         n675, n676, n677, n678, n679, n680, n681, n682, n686, n687, n688,
         n689, n694, n695, n696, n697, n701, n702, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n723,
         n724, n728, n729, n730, n734, n735, n736, n737, n738, n742, n743,
         n744, n745, n746, n750, n751, n753, n754, n758, n760, n761, n762,
         n763, n764, n765, n770, n771, n778, n783, n786, n788, n789, n790,
         n791, n797, n799, n800, n821, n822, n823, n824, n825, n826, n827,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2268, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2302, n2303, n2304, n2305, n2306, n2308,
         n2309, n2310, n2315, n2316, n2317, n2318, n2319, n2320, n2323, n2324,
         n2325, n2326, n2328, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2343, n2344, n2347, n2348, n2349, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2361, n2362, n2365, n2366, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2381, n2382, n2383,
         n2384, n2386, n2389, n2390, n2391, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2409, n2410,
         n2411, n2412, n2413, n2414, n2417, n2418, n2419, n2420, n2423, n2424,
         n2425, n2426, n2427, n2432, n2433, n2434, n2435, n2436, n2439, n2440,
         n2441, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3625, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068;

  XOR2X1 U232 ( .A(n294), .B(n4902), .Y(product[63]) );
  XNOR2X1 U234 ( .A(n301), .B(n4644), .Y(product[62]) );
  OAI21X1 U235 ( .A(n3954), .B(n4922), .C(n3948), .Y(n294) );
  AOI21X1 U237 ( .A(n305), .B(n4919), .C(n298), .Y(n296) );
  XNOR2X1 U244 ( .A(n312), .B(n4711), .Y(product[61]) );
  OAI21X1 U245 ( .A(n304), .B(n3940), .C(n303), .Y(n301) );
  OAI21X1 U249 ( .A(n4420), .B(n4758), .C(n4341), .Y(n305) );
  AOI21X1 U251 ( .A(n230), .B(n4557), .C(n309), .Y(n307) );
  OAI21X1 U253 ( .A(n4900), .B(n4608), .C(n4899), .Y(n309) );
  XNOR2X1 U258 ( .A(n323), .B(n4709), .Y(product[60]) );
  OAI21X1 U259 ( .A(n4357), .B(n4922), .C(n4340), .Y(n312) );
  AOI21X1 U261 ( .A(n419), .B(n317), .C(n316), .Y(n314) );
  AOI21X1 U265 ( .A(n371), .B(n4409), .C(n320), .Y(n318) );
  OAI21X1 U267 ( .A(n4898), .B(n4664), .C(n4897), .Y(n320) );
  XNOR2X1 U272 ( .A(n334), .B(n4585), .Y(product[59]) );
  OAI21X1 U273 ( .A(n3953), .B(n3940), .C(n4339), .Y(n323) );
  AOI21X1 U275 ( .A(n367), .B(n326), .C(n327), .Y(n325) );
  AOI21X1 U279 ( .A(n353), .B(n4732), .C(n331), .Y(n329) );
  OAI21X1 U281 ( .A(n4896), .B(n4893), .C(n4895), .Y(n331) );
  XNOR2X1 U286 ( .A(n341), .B(n4710), .Y(product[58]) );
  OAI21X1 U287 ( .A(n3952), .B(n4922), .C(n4337), .Y(n334) );
  AOI21X1 U289 ( .A(n345), .B(n763), .C(n338), .Y(n336) );
  XNOR2X1 U296 ( .A(n356), .B(n4712), .Y(product[57]) );
  OAI21X1 U297 ( .A(n344), .B(n4763), .C(n343), .Y(n341) );
  OAI21X1 U301 ( .A(n4419), .B(n4758), .C(n4335), .Y(n345) );
  AOI21X1 U303 ( .A(n230), .B(n4556), .C(n349), .Y(n347) );
  OAI21X1 U305 ( .A(n350), .B(n373), .C(n351), .Y(n349) );
  OAI21X1 U309 ( .A(n4892), .B(n4889), .C(n4891), .Y(n353) );
  XNOR2X1 U314 ( .A(n363), .B(n4648), .Y(product[56]) );
  OAI21X1 U315 ( .A(n3946), .B(n4763), .C(n4334), .Y(n356) );
  AOI21X1 U317 ( .A(n367), .B(n765), .C(n360), .Y(n358) );
  XNOR2X1 U324 ( .A(n382), .B(n4589), .Y(product[55]) );
  OAI21X1 U325 ( .A(n366), .B(n4763), .C(n365), .Y(n363) );
  OAI21X1 U329 ( .A(n4413), .B(n4758), .C(n4332), .Y(n367) );
  AOI21X1 U331 ( .A(n230), .B(n4628), .C(n371), .Y(n369) );
  OAI21X1 U337 ( .A(n4736), .B(n4666), .C(n4331), .Y(n371) );
  AOI21X1 U339 ( .A(n4918), .B(n388), .C(n379), .Y(n377) );
  XNOR2X1 U346 ( .A(n391), .B(n4588), .Y(product[54]) );
  OAI21X1 U347 ( .A(n3951), .B(n4763), .C(n4330), .Y(n382) );
  AOI21X1 U349 ( .A(n395), .B(n4917), .C(n388), .Y(n384) );
  XNOR2X1 U358 ( .A(n406), .B(n4715), .Y(product[53]) );
  OAI21X1 U359 ( .A(n394), .B(n3940), .C(n393), .Y(n391) );
  OAI21X1 U363 ( .A(n4418), .B(n4758), .C(n4328), .Y(n395) );
  AOI21X1 U365 ( .A(n230), .B(n400), .C(n399), .Y(n397) );
  AOI21X1 U369 ( .A(n4916), .B(n412), .C(n403), .Y(n401) );
  XNOR2X1 U376 ( .A(n415), .B(n4536), .Y(product[52]) );
  OAI21X1 U377 ( .A(n4469), .B(n4922), .C(n4327), .Y(n406) );
  AOI21X1 U379 ( .A(n419), .B(n4915), .C(n412), .Y(n408) );
  XNOR2X1 U388 ( .A(n430), .B(n4647), .Y(product[51]) );
  OAI21X1 U389 ( .A(n418), .B(n3940), .C(n417), .Y(n415) );
  OAI21X1 U393 ( .A(n420), .B(n4758), .C(n421), .Y(n419) );
  OAI21X1 U397 ( .A(n4663), .B(n4615), .C(n4326), .Y(n230) );
  AOI21X1 U399 ( .A(n4731), .B(n447), .C(n427), .Y(n425) );
  OAI21X1 U401 ( .A(n4884), .B(n4881), .C(n4883), .Y(n427) );
  XNOR2X1 U406 ( .A(n437), .B(n4590), .Y(product[50]) );
  OAI21X1 U407 ( .A(n4356), .B(n4922), .C(n4325), .Y(n430) );
  AOI21X1 U409 ( .A(n441), .B(n771), .C(n434), .Y(n432) );
  XNOR2X1 U416 ( .A(n450), .B(n4499), .Y(product[49]) );
  OAI21X1 U417 ( .A(n440), .B(n3940), .C(n439), .Y(n437) );
  OAI21X1 U421 ( .A(n4559), .B(n4758), .C(n4324), .Y(n441) );
  AOI21X1 U423 ( .A(n456), .B(n4914), .C(n447), .Y(n443) );
  OAI21X1 U433 ( .A(n4923), .B(n4455), .C(n4323), .Y(n450) );
  AOI21X1 U435 ( .A(n472), .B(n457), .C(n456), .Y(n452) );
  AOI21X1 U441 ( .A(n4913), .B(n465), .C(n460), .Y(n458) );
  XNOR2X1 U448 ( .A(n3931), .B(n4479), .Y(product[47]) );
  AOI21X1 U449 ( .A(n468), .B(n4912), .C(n465), .Y(n463) );
  XOR2X1 U456 ( .A(n4458), .B(n4656), .Y(product[46]) );
  OAI21X1 U457 ( .A(n4689), .B(n4923), .C(n4758), .Y(n468) );
  AOI21X1 U463 ( .A(n4482), .B(n508), .C(n476), .Y(n470) );
  OAI21X1 U465 ( .A(n4614), .B(n4665), .C(n4759), .Y(n476) );
  AOI21X1 U467 ( .A(n4911), .B(n485), .C(n480), .Y(n478) );
  XNOR2X1 U474 ( .A(n488), .B(n4478), .Y(product[45]) );
  AOI21X1 U475 ( .A(n488), .B(n4910), .C(n485), .Y(n483) );
  XOR2X1 U482 ( .A(n4582), .B(n4717), .Y(product[44]) );
  OAI21X1 U483 ( .A(n4450), .B(n4763), .C(n4451), .Y(n488) );
  AOI21X1 U485 ( .A(n508), .B(n493), .C(n492), .Y(n490) );
  AOI21X1 U489 ( .A(n4909), .B(n501), .C(n496), .Y(n494) );
  XNOR2X1 U496 ( .A(n504), .B(n4646), .Y(product[43]) );
  AOI21X1 U497 ( .A(n504), .B(n778), .C(n501), .Y(n499) );
  OAI21X1 U505 ( .A(n507), .B(n4923), .C(n506), .Y(n504) );
  OAI21X1 U513 ( .A(n4625), .B(n4678), .C(n4550), .Y(n508) );
  XOR2X1 U526 ( .A(n3960), .B(n4389), .Y(product[40]) );
  AOI21X1 U528 ( .A(n4760), .B(n3938), .C(n523), .Y(n227) );
  OAI21X1 U530 ( .A(n4670), .B(n4417), .C(n4322), .Y(n523) );
  AOI21X1 U532 ( .A(n541), .B(n3925), .C(n527), .Y(n525) );
  OAI21X1 U534 ( .A(n4677), .B(n4751), .C(n4607), .Y(n527) );
  XNOR2X1 U539 ( .A(n3934), .B(n4388), .Y(product[39]) );
  AOI21X1 U540 ( .A(n535), .B(n3929), .C(n534), .Y(n530) );
  XOR2X1 U547 ( .A(n4502), .B(n4501), .Y(product[38]) );
  OAI21X1 U548 ( .A(n4358), .B(n3933), .C(n4320), .Y(n535) );
  AOI21X1 U550 ( .A(n553), .B(n4764), .C(n541), .Y(n537) );
  OAI21X1 U554 ( .A(n4739), .B(n4609), .C(n4549), .Y(n541) );
  XNOR2X1 U559 ( .A(n549), .B(n4535), .Y(product[37]) );
  AOI21X1 U560 ( .A(n549), .B(n3935), .C(n548), .Y(n544) );
  XOR2X1 U567 ( .A(n4538), .B(n4537), .Y(product[36]) );
  OAI21X1 U568 ( .A(n575), .B(n4621), .C(n4670), .Y(n549) );
  AOI21X1 U574 ( .A(n569), .B(n4553), .C(n557), .Y(n551) );
  OAI21X1 U576 ( .A(n4871), .B(n4743), .C(n4606), .Y(n557) );
  XNOR2X1 U581 ( .A(n4761), .B(n4716), .Y(product[35]) );
  AOI21X1 U582 ( .A(n565), .B(n786), .C(n562), .Y(n560) );
  XNOR2X1 U589 ( .A(n572), .B(n4645), .Y(product[34]) );
  OAI21X1 U590 ( .A(n568), .B(n3933), .C(n567), .Y(n565) );
  OAI21X1 U594 ( .A(n4869), .B(n4742), .C(n4599), .Y(n569) );
  XOR2X1 U599 ( .A(n3928), .B(n4722), .Y(product[33]) );
  OAI21X1 U600 ( .A(n4870), .B(n3933), .C(n4869), .Y(n572) );
  OAI21X1 U607 ( .A(n4610), .B(n4733), .C(n4611), .Y(n576) );
  AOI21X1 U609 ( .A(n588), .B(n4612), .C(n580), .Y(n578) );
  OAI21X1 U611 ( .A(n4865), .B(n4868), .C(n4867), .Y(n580) );
  XOR2X1 U616 ( .A(n4668), .B(n4723), .Y(product[31]) );
  OAI21X1 U617 ( .A(n4866), .B(n4668), .C(n4865), .Y(n583) );
  XOR2X1 U622 ( .A(n4470), .B(n4721), .Y(product[30]) );
  AOI21X1 U623 ( .A(n605), .B(n4552), .C(n588), .Y(n586) );
  OAI21X1 U625 ( .A(n4864), .B(n4730), .C(n4863), .Y(n588) );
  XOR2X1 U630 ( .A(n4581), .B(n4657), .Y(product[29]) );
  AOI21X1 U631 ( .A(n605), .B(n594), .C(n593), .Y(n591) );
  AOI21X1 U635 ( .A(n4908), .B(n602), .C(n597), .Y(n595) );
  XNOR2X1 U642 ( .A(n605), .B(n4713), .Y(product[28]) );
  AOI21X1 U643 ( .A(n605), .B(n4907), .C(n602), .Y(n600) );
  XOR2X1 U650 ( .A(n4580), .B(n4655), .Y(product[27]) );
  AOI21X1 U652 ( .A(n635), .B(n4734), .C(n608), .Y(n606) );
  OAI21X1 U654 ( .A(n4555), .B(n4735), .C(n4468), .Y(n608) );
  AOI21X1 U656 ( .A(n4906), .B(n617), .C(n612), .Y(n610) );
  XNOR2X1 U663 ( .A(n620), .B(n4643), .Y(product[26]) );
  AOI21X1 U664 ( .A(n620), .B(n4905), .C(n617), .Y(n615) );
  XNOR2X1 U671 ( .A(n627), .B(n4714), .Y(product[25]) );
  OAI21X1 U672 ( .A(n4667), .B(n634), .C(n4555), .Y(n620) );
  AOI21X1 U674 ( .A(n4904), .B(n631), .C(n624), .Y(n622) );
  XOR2X1 U681 ( .A(n634), .B(n4720), .Y(product[24]) );
  OAI21X1 U682 ( .A(n4857), .B(n634), .C(n4856), .Y(n627) );
  XOR2X1 U691 ( .A(n4654), .B(n4653), .Y(product[23]) );
  OAI21X1 U693 ( .A(n4849), .B(n4490), .C(n4489), .Y(n635) );
  AOI21X1 U695 ( .A(n644), .B(n4903), .C(n639), .Y(n637) );
  XOR2X1 U702 ( .A(n4718), .B(n4719), .Y(product[22]) );
  AOI21X1 U703 ( .A(n652), .B(n4707), .C(n644), .Y(n642) );
  OAI21X1 U705 ( .A(n4851), .B(n4854), .C(n4853), .Y(n644) );
  XNOR2X1 U710 ( .A(n652), .B(n4583), .Y(product[21]) );
  AOI21X1 U711 ( .A(n652), .B(n800), .C(n649), .Y(n647) );
  XNOR2X1 U718 ( .A(n4848), .B(n4850), .Y(product[20]) );
  AOI21X1 U720 ( .A(n662), .B(n4351), .C(n655), .Y(n653) );
  OAI21X1 U722 ( .A(n4753), .B(n4623), .C(n4546), .Y(n655) );
  XOR2X1 U727 ( .A(n661), .B(n4593), .Y(product[19]) );
  OAI21X1 U728 ( .A(n4680), .B(n661), .C(n4753), .Y(n658) );
  XOR2X1 U733 ( .A(n4652), .B(n4651), .Y(product[18]) );
  OAI21X1 U735 ( .A(n4355), .B(n4402), .C(n4319), .Y(n662) );
  AOI21X1 U737 ( .A(n4808), .B(n673), .C(n668), .Y(n664) );
  XNOR2X1 U744 ( .A(n4401), .B(n4708), .Y(product[17]) );
  AOI21X1 U745 ( .A(n4401), .B(n4805), .C(n673), .Y(n669) );
  XNOR2X1 U752 ( .A(n680), .B(n4460), .Y(product[16]) );
  AOI21X1 U754 ( .A(n3945), .B(n695), .C(n677), .Y(n675) );
  OAI21X1 U756 ( .A(n4740), .B(n4558), .C(n4661), .Y(n677) );
  XNOR2X1 U761 ( .A(n687), .B(n4472), .Y(product[15]) );
  OAI21X1 U762 ( .A(n4613), .B(n694), .C(n4558), .Y(n680) );
  AOI21X1 U764 ( .A(n4806), .B(n689), .C(n686), .Y(n682) );
  XOR2X1 U771 ( .A(n694), .B(n4500), .Y(product[14]) );
  OAI21X1 U772 ( .A(n4662), .B(n694), .C(n4738), .Y(n687) );
  XOR2X1 U781 ( .A(n4650), .B(n4649), .Y(product[13]) );
  OAI21X1 U783 ( .A(n4354), .B(n4511), .C(n4318), .Y(n695) );
  AOI21X1 U785 ( .A(n4807), .B(n706), .C(n701), .Y(n697) );
  XNOR2X1 U792 ( .A(n707), .B(n4584), .Y(product[12]) );
  AOI21X1 U793 ( .A(n707), .B(n4816), .C(n706), .Y(n702) );
  XNOR2X1 U800 ( .A(n713), .B(n4471), .Y(product[11]) );
  AOI21X1 U802 ( .A(n4512), .B(n717), .C(n710), .Y(n708) );
  OAI21X1 U804 ( .A(n4752), .B(n4681), .C(n4547), .Y(n710) );
  XOR2X1 U809 ( .A(n4641), .B(n716), .Y(product[10]) );
  OAI21X1 U810 ( .A(n4619), .B(n716), .C(n4752), .Y(n713) );
  XOR2X1 U815 ( .A(n4591), .B(n4592), .Y(product[9]) );
  OAI21X1 U817 ( .A(n4551), .B(n4457), .C(n4456), .Y(n717) );
  AOI21X1 U819 ( .A(n4817), .B(n728), .C(n723), .Y(n719) );
  XNOR2X1 U826 ( .A(n729), .B(n4642), .Y(product[8]) );
  AOI21X1 U827 ( .A(n729), .B(n4815), .C(n728), .Y(n724) );
  XNOR2X1 U834 ( .A(n4491), .B(n735), .Y(product[7]) );
  AOI21X1 U836 ( .A(n4820), .B(n735), .C(n734), .Y(n730) );
  XOR2X1 U843 ( .A(n4529), .B(n4617), .Y(product[6]) );
  OAI21X1 U844 ( .A(n4617), .B(n4729), .C(n4660), .Y(n735) );
  XNOR2X1 U849 ( .A(n4492), .B(n743), .Y(product[5]) );
  AOI21X1 U850 ( .A(n743), .B(n4819), .C(n742), .Y(n738) );
  XOR2X1 U857 ( .A(n4493), .B(n4669), .Y(product[4]) );
  OAI21X1 U858 ( .A(n4728), .B(n4669), .C(n4545), .Y(n743) );
  XNOR2X1 U863 ( .A(n4527), .B(n4737), .Y(product[3]) );
  AOI21X1 U864 ( .A(n4818), .B(n4737), .C(n750), .Y(n746) );
  XOR2X1 U871 ( .A(n4827), .B(n4616), .Y(product[2]) );
  FAX1 U886 ( .A(n5068), .B(n2517), .C(n827), .YC(n823), .YS(n824) );
  FAX1 U887 ( .A(n2518), .B(n831), .C(n2541), .YC(n825), .YS(n826) );
  FAX1 U889 ( .A(n831), .B(n2542), .C(n834), .YC(n829), .YS(n830) );
  FAX1 U891 ( .A(n2543), .B(n835), .C(n838), .YC(n832), .YS(n833) );
  FAX1 U892 ( .A(n5065), .B(n840), .C(n2519), .YC(n834), .YS(n835) );
  FAX1 U893 ( .A(n2544), .B(n839), .C(n844), .YC(n836), .YS(n837) );
  FAX1 U894 ( .A(n2520), .B(n846), .C(n2576), .YC(n838), .YS(n839) );
  FAX1 U896 ( .A(n851), .B(n845), .C(n849), .YC(n842), .YS(n843) );
  FAX1 U897 ( .A(n846), .B(n2545), .C(n2577), .YC(n844), .YS(n845) );
  FAX1 U899 ( .A(n857), .B(n850), .C(n855), .YC(n847), .YS(n848) );
  FAX1 U900 ( .A(n2578), .B(n2546), .C(n852), .YC(n849), .YS(n850) );
  FAX1 U901 ( .A(n5062), .B(n859), .C(n2521), .YC(n851), .YS(n852) );
  FAX1 U902 ( .A(n865), .B(n856), .C(n863), .YC(n853), .YS(n854) );
  FAX1 U903 ( .A(n2579), .B(n2547), .C(n858), .YC(n855), .YS(n856) );
  FAX1 U904 ( .A(n2522), .B(n867), .C(n2611), .YC(n857), .YS(n858) );
  FAX1 U906 ( .A(n866), .B(n870), .C(n864), .YC(n861), .YS(n862) );
  FAX1 U907 ( .A(n2612), .B(n874), .C(n872), .YC(n863), .YS(n864) );
  FAX1 U908 ( .A(n867), .B(n2580), .C(n2548), .YC(n865), .YS(n866) );
  FAX1 U910 ( .A(n873), .B(n871), .C(n878), .YC(n868), .YS(n869) );
  FAX1 U911 ( .A(n875), .B(n882), .C(n880), .YC(n870), .YS(n871) );
  FAX1 U912 ( .A(n2549), .B(n2581), .C(n2613), .YC(n872), .YS(n873) );
  FAX1 U913 ( .A(n5059), .B(n884), .C(n2523), .YC(n874), .YS(n875) );
  FAX1 U914 ( .A(n890), .B(n879), .C(n888), .YC(n876), .YS(n877) );
  FAX1 U915 ( .A(n883), .B(n892), .C(n881), .YC(n878), .YS(n879) );
  FAX1 U916 ( .A(n2550), .B(n2582), .C(n2614), .YC(n880), .YS(n881) );
  FAX1 U917 ( .A(n2524), .B(n894), .C(n2646), .YC(n882), .YS(n883) );
  FAX1 U919 ( .A(n899), .B(n889), .C(n897), .YC(n886), .YS(n887) );
  FAX1 U920 ( .A(n901), .B(n893), .C(n891), .YC(n888), .YS(n889) );
  FAX1 U921 ( .A(n2551), .B(n2647), .C(n903), .YC(n890), .YS(n891) );
  FAX1 U922 ( .A(n894), .B(n2615), .C(n2583), .YC(n892), .YS(n893) );
  FAX1 U924 ( .A(n909), .B(n898), .C(n907), .YC(n895), .YS(n896) );
  FAX1 U925 ( .A(n911), .B(n902), .C(n900), .YC(n897), .YS(n898) );
  FAX1 U926 ( .A(n2616), .B(n904), .C(n913), .YC(n899), .YS(n900) );
  FAX1 U927 ( .A(n2584), .B(n2648), .C(n2552), .YC(n901), .YS(n902) );
  FAX1 U928 ( .A(n5056), .B(n915), .C(n2525), .YC(n903), .YS(n904) );
  FAX1 U929 ( .A(n921), .B(n908), .C(n919), .YC(n905), .YS(n906) );
  FAX1 U930 ( .A(n923), .B(n912), .C(n910), .YC(n907), .YS(n908) );
  FAX1 U931 ( .A(n2617), .B(n914), .C(n925), .YC(n909), .YS(n910) );
  FAX1 U932 ( .A(n2585), .B(n2649), .C(n2553), .YC(n911), .YS(n912) );
  FAX1 U933 ( .A(n2526), .B(n927), .C(n2681), .YC(n913), .YS(n914) );
  FAX1 U935 ( .A(n922), .B(n930), .C(n920), .YC(n917), .YS(n918) );
  FAX1 U936 ( .A(n926), .B(n924), .C(n932), .YC(n919), .YS(n920) );
  FAX1 U937 ( .A(n2586), .B(n936), .C(n934), .YC(n921), .YS(n922) );
  FAX1 U938 ( .A(n2650), .B(n2554), .C(n2682), .YC(n923), .YS(n924) );
  FAX1 U939 ( .A(n927), .B(n938), .C(n2618), .YC(n925), .YS(n926) );
  FAX1 U941 ( .A(n933), .B(n942), .C(n931), .YC(n928), .YS(n929) );
  FAX1 U942 ( .A(n937), .B(n946), .C(n944), .YC(n930), .YS(n931) );
  FAX1 U943 ( .A(n950), .B(n948), .C(n935), .YC(n932), .YS(n933) );
  FAX1 U944 ( .A(n2619), .B(n2651), .C(n2683), .YC(n934), .YS(n935) );
  FAX1 U945 ( .A(n2587), .B(n2555), .C(n939), .YC(n936), .YS(n937) );
  FAX1 U946 ( .A(n5053), .B(n2527), .C(n952), .YC(n938), .YS(n939) );
  FAX1 U947 ( .A(n945), .B(n956), .C(n943), .YC(n940), .YS(n941) );
  FAX1 U948 ( .A(n947), .B(n960), .C(n958), .YC(n942), .YS(n943) );
  FAX1 U949 ( .A(n964), .B(n962), .C(n949), .YC(n944), .YS(n945) );
  FAX1 U950 ( .A(n2620), .B(n2556), .C(n951), .YC(n946), .YS(n947) );
  FAX1 U951 ( .A(n2588), .B(n2684), .C(n2652), .YC(n948), .YS(n949) );
  FAX1 U952 ( .A(n966), .B(n2528), .C(n2716), .YC(n950), .YS(n951) );
  FAX1 U954 ( .A(n959), .B(n969), .C(n957), .YC(n954), .YS(n955) );
  FAX1 U955 ( .A(n961), .B(n973), .C(n971), .YC(n956), .YS(n957) );
  FAX1 U956 ( .A(n975), .B(n965), .C(n963), .YC(n958), .YS(n959) );
  FAX1 U957 ( .A(n2557), .B(n979), .C(n977), .YC(n960), .YS(n961) );
  FAX1 U958 ( .A(n2589), .B(n2685), .C(n2717), .YC(n962), .YS(n963) );
  FAX1 U959 ( .A(n966), .B(n2653), .C(n2621), .YC(n964), .YS(n965) );
  FAX1 U961 ( .A(n972), .B(n983), .C(n970), .YC(n967), .YS(n968) );
  FAX1 U962 ( .A(n987), .B(n974), .C(n985), .YC(n969), .YS(n970) );
  FAX1 U963 ( .A(n989), .B(n978), .C(n976), .YC(n971), .YS(n972) );
  FAX1 U964 ( .A(n980), .B(n993), .C(n991), .YC(n973), .YS(n974) );
  FAX1 U965 ( .A(n2718), .B(n2590), .C(n2686), .YC(n975), .YS(n976) );
  FAX1 U966 ( .A(n2529), .B(n2622), .C(n2654), .YC(n977), .YS(n978) );
  FAX1 U967 ( .A(n5050), .B(n995), .C(n2558), .YC(n979), .YS(n980) );
  FAX1 U968 ( .A(n986), .B(n984), .C(n999), .YC(n981), .YS(n982) );
  FAX1 U969 ( .A(n1003), .B(n988), .C(n1001), .YC(n983), .YS(n984) );
  FAX1 U970 ( .A(n1005), .B(n990), .C(n992), .YC(n985), .YS(n986) );
  FAX1 U971 ( .A(n1009), .B(n994), .C(n1007), .YC(n987), .YS(n988) );
  FAX1 U972 ( .A(n2719), .B(n2655), .C(n2687), .YC(n989), .YS(n990) );
  FAX1 U973 ( .A(n2623), .B(n2591), .C(n2559), .YC(n991), .YS(n992) );
  FAX1 U974 ( .A(n996), .B(n1011), .C(n2751), .YC(n993), .YS(n994) );
  FAX1 U976 ( .A(n1017), .B(n1000), .C(n1015), .YC(n997), .YS(n998) );
  FAX1 U977 ( .A(n1019), .B(n1004), .C(n1002), .YC(n999), .YS(n1000) );
  FAX1 U978 ( .A(n1006), .B(n1008), .C(n1021), .YC(n1001), .YS(n1002) );
  FAX1 U979 ( .A(n1010), .B(n1025), .C(n1023), .YC(n1003), .YS(n1004) );
  FAX1 U980 ( .A(n2688), .B(n2592), .C(n2624), .YC(n1005), .YS(n1006) );
  FAX1 U981 ( .A(n2656), .B(n2720), .C(n2752), .YC(n1007), .YS(n1008) );
  FAX1 U982 ( .A(n2560), .B(n1012), .C(n1027), .YC(n1009), .YS(n1010) );
  FAX1 U984 ( .A(n1033), .B(n1016), .C(n1031), .YC(n1013), .YS(n1014) );
  FAX1 U985 ( .A(n1035), .B(n1020), .C(n1018), .YC(n1015), .YS(n1016) );
  FAX1 U986 ( .A(n1039), .B(n1022), .C(n1037), .YC(n1017), .YS(n1018) );
  FAX1 U987 ( .A(n1041), .B(n1026), .C(n1024), .YC(n1019), .YS(n1020) );
  FAX1 U988 ( .A(n2721), .B(n2689), .C(n1043), .YC(n1021), .YS(n1022) );
  FAX1 U989 ( .A(n2753), .B(n1028), .C(n2561), .YC(n1023), .YS(n1024) );
  FAX1 U990 ( .A(n2593), .B(n2657), .C(n2625), .YC(n1025), .YS(n1026) );
  FAX1 U991 ( .A(n5047), .B(n1045), .C(n2530), .YC(n1027), .YS(n1028) );
  FAX1 U992 ( .A(n1051), .B(n1032), .C(n1049), .YC(n1029), .YS(n1030) );
  FAX1 U993 ( .A(n1053), .B(n1036), .C(n1034), .YC(n1031), .YS(n1032) );
  FAX1 U994 ( .A(n1057), .B(n1038), .C(n1055), .YC(n1033), .YS(n1034) );
  FAX1 U995 ( .A(n1059), .B(n1042), .C(n1040), .YC(n1035), .YS(n1036) );
  FAX1 U996 ( .A(n2690), .B(n1044), .C(n1061), .YC(n1037), .YS(n1038) );
  FAX1 U997 ( .A(n2722), .B(n2626), .C(n2658), .YC(n1039), .YS(n1040) );
  FAX1 U998 ( .A(n2786), .B(n2754), .C(n2594), .YC(n1041), .YS(n1042) );
  FAX1 U999 ( .A(n1063), .B(n2531), .C(n2562), .YC(n1043), .YS(n1044) );
  FAX1 U1001 ( .A(n4839), .B(n4838), .C(n4840), .YC(n1047), .YS(n1048) );
  FAX1 U1002 ( .A(n1070), .B(n1054), .C(n1068), .YC(n1049), .YS(n1050) );
  FAX1 U1003 ( .A(n1058), .B(n1072), .C(n1056), .YC(n1051), .YS(n1052) );
  FAX1 U1004 ( .A(n1076), .B(n1074), .C(n1060), .YC(n1053), .YS(n1054) );
  FAX1 U1005 ( .A(n2723), .B(n1078), .C(n1062), .YC(n1055), .YS(n1056) );
  FAX1 U1006 ( .A(n2755), .B(n2627), .C(n2691), .YC(n1057), .YS(n1058) );
  FAX1 U1007 ( .A(n2659), .B(n2787), .C(n2563), .YC(n1059), .YS(n1060) );
  FAX1 U1008 ( .A(n1063), .B(n2595), .C(n1080), .YC(n1061), .YS(n1062) );
  FAX1 U1010 ( .A(n4836), .B(n4833), .C(n4837), .YC(n1064), .YS(n1065) );
  FAX1 U1011 ( .A(n1088), .B(n1071), .C(n1086), .YC(n1066), .YS(n1067) );
  FAX1 U1012 ( .A(n1075), .B(n1090), .C(n1073), .YC(n1068), .YS(n1069) );
  FAX1 U1013 ( .A(n1094), .B(n1092), .C(n1077), .YC(n1070), .YS(n1071) );
  FAX1 U1014 ( .A(n1098), .B(n1096), .C(n1079), .YC(n1072), .YS(n1073) );
  FAX1 U1015 ( .A(n2756), .B(n2692), .C(n2724), .YC(n1074), .YS(n1075) );
  FAX1 U1016 ( .A(n2660), .B(n2788), .C(n2596), .YC(n1076), .YS(n1077) );
  FAX1 U1017 ( .A(n2628), .B(n2564), .C(n1081), .YC(n1078), .YS(n1079) );
  FAX1 U1018 ( .A(n5044), .B(n5040), .C(n2532), .YC(n1080), .YS(n1081) );
  FAX1 U1019 ( .A(n1087), .B(n1102), .C(n1085), .YC(n1082), .YS(n1083) );
  FAX1 U1020 ( .A(n1106), .B(n1089), .C(n1104), .YC(n1084), .YS(n1085) );
  FAX1 U1021 ( .A(n1093), .B(n1108), .C(n1091), .YC(n1086), .YS(n1087) );
  FAX1 U1022 ( .A(n1112), .B(n1110), .C(n1095), .YC(n1088), .YS(n1089) );
  FAX1 U1023 ( .A(n1099), .B(n1114), .C(n1097), .YC(n1090), .YS(n1091) );
  FAX1 U1024 ( .A(n2789), .B(n2725), .C(n2757), .YC(n1092), .YS(n1093) );
  FAX1 U1025 ( .A(n2661), .B(n2693), .C(n2629), .YC(n1094), .YS(n1095) );
  FAX1 U1026 ( .A(n2565), .B(n2821), .C(n1116), .YC(n1096), .YS(n1097) );
  FAX1 U1027 ( .A(n5038), .B(n2533), .C(n2597), .YC(n1098), .YS(n1099) );
  FAX1 U1028 ( .A(n1105), .B(n1120), .C(n1103), .YC(n1100), .YS(n1101) );
  FAX1 U1029 ( .A(n1124), .B(n1107), .C(n1122), .YC(n1102), .YS(n1103) );
  FAX1 U1030 ( .A(n1113), .B(n1126), .C(n1109), .YC(n1104), .YS(n1105) );
  FAX1 U1031 ( .A(n1115), .B(n1111), .C(n1128), .YC(n1106), .YS(n1107) );
  FAX1 U1032 ( .A(n1134), .B(n1132), .C(n1130), .YC(n1108), .YS(n1109) );
  FAX1 U1033 ( .A(n2758), .B(n2726), .C(n2822), .YC(n1110), .YS(n1111) );
  FAX1 U1034 ( .A(n2790), .B(n1117), .C(n2598), .YC(n1112), .YS(n1113) );
  FAX1 U1035 ( .A(n2630), .B(n2694), .C(n2662), .YC(n1114), .YS(n1115) );
  FAX1 U1036 ( .A(n5038), .B(n2534), .C(n2566), .YC(n1116), .YS(n1117) );
  FAX1 U1037 ( .A(n1123), .B(n1138), .C(n1121), .YC(n1118), .YS(n1119) );
  FAX1 U1038 ( .A(n1142), .B(n1125), .C(n1140), .YC(n1120), .YS(n1121) );
  FAX1 U1039 ( .A(n1129), .B(n1144), .C(n1127), .YC(n1122), .YS(n1123) );
  FAX1 U1040 ( .A(n1148), .B(n1146), .C(n1131), .YC(n1124), .YS(n1125) );
  FAX1 U1041 ( .A(n1135), .B(n1150), .C(n1133), .YC(n1126), .YS(n1127) );
  FAX1 U1042 ( .A(n2791), .B(n2759), .C(n1152), .YC(n1128), .YS(n1129) );
  FAX1 U1043 ( .A(n2823), .B(n2727), .C(n2631), .YC(n1130), .YS(n1131) );
  FAX1 U1044 ( .A(n2663), .B(n2599), .C(n2695), .YC(n1132), .YS(n1133) );
  FAX1 U1045 ( .A(n5038), .B(n2535), .C(n2567), .YC(n1134), .YS(n1135) );
  FAX1 U1046 ( .A(n1141), .B(n1156), .C(n1139), .YC(n1136), .YS(n1137) );
  FAX1 U1047 ( .A(n1160), .B(n1143), .C(n1158), .YC(n1138), .YS(n1139) );
  FAX1 U1048 ( .A(n1147), .B(n1162), .C(n1145), .YC(n1140), .YS(n1141) );
  FAX1 U1049 ( .A(n1166), .B(n1164), .C(n1149), .YC(n1142), .YS(n1143) );
  FAX1 U1050 ( .A(n1153), .B(n1168), .C(n1151), .YC(n1144), .YS(n1145) );
  FAX1 U1051 ( .A(n2792), .B(n2728), .C(n2760), .YC(n1146), .YS(n1147) );
  FAX1 U1052 ( .A(n2824), .B(n1170), .C(n2664), .YC(n1148), .YS(n1149) );
  FAX1 U1053 ( .A(n2632), .B(n2696), .C(n2856), .YC(n1150), .YS(n1151) );
  FAX1 U1054 ( .A(n2536), .B(n2568), .C(n2600), .YC(n1152), .YS(n1153) );
  FAX1 U1055 ( .A(n1159), .B(n1174), .C(n1157), .YC(n1154), .YS(n1155) );
  FAX1 U1056 ( .A(n1178), .B(n1161), .C(n1176), .YC(n1156), .YS(n1157) );
  FAX1 U1057 ( .A(n1165), .B(n1180), .C(n1163), .YC(n1158), .YS(n1159) );
  FAX1 U1058 ( .A(n1182), .B(n1169), .C(n1167), .YC(n1160), .YS(n1161) );
  FAX1 U1059 ( .A(n1188), .B(n1186), .C(n1184), .YC(n1162), .YS(n1163) );
  FAX1 U1060 ( .A(n2825), .B(n2793), .C(n2857), .YC(n1164), .YS(n1165) );
  FAX1 U1061 ( .A(n2761), .B(n2633), .C(n1171), .YC(n1166), .YS(n1167) );
  FAX1 U1062 ( .A(n2665), .B(n2729), .C(n2697), .YC(n1168), .YS(n1169) );
  FAX1 U1063 ( .A(n2537), .B(n2569), .C(n2601), .YC(n1170), .YS(n1171) );
  FAX1 U1064 ( .A(n1177), .B(n1192), .C(n1175), .YC(n1172), .YS(n1173) );
  FAX1 U1065 ( .A(n1196), .B(n1179), .C(n1194), .YC(n1174), .YS(n1175) );
  FAX1 U1066 ( .A(n1183), .B(n1198), .C(n1181), .YC(n1176), .YS(n1177) );
  FAX1 U1067 ( .A(n1202), .B(n1200), .C(n1185), .YC(n1178), .YS(n1179) );
  FAX1 U1068 ( .A(n1189), .B(n1204), .C(n1187), .YC(n1180), .YS(n1181) );
  FAX1 U1069 ( .A(n2858), .B(n2794), .C(n2826), .YC(n1182), .YS(n1183) );
  FAX1 U1070 ( .A(n2730), .B(n2762), .C(n2666), .YC(n1184), .YS(n1185) );
  FAX1 U1071 ( .A(n2698), .B(n2634), .C(n1206), .YC(n1186), .YS(n1187) );
  FAX1 U1072 ( .A(n2538), .B(n2570), .C(n2602), .YC(n1188), .YS(n1189) );
  FAX1 U1073 ( .A(n1195), .B(n1210), .C(n1193), .YC(n1190), .YS(n1191) );
  FAX1 U1074 ( .A(n1214), .B(n1197), .C(n1212), .YC(n1192), .YS(n1193) );
  FAX1 U1075 ( .A(n1218), .B(n1216), .C(n1199), .YC(n1194), .YS(n1195) );
  FAX1 U1076 ( .A(n1220), .B(n1203), .C(n1201), .YC(n1196), .YS(n1197) );
  FAX1 U1077 ( .A(n2795), .B(n2731), .C(n1205), .YC(n1198), .YS(n1199) );
  FAX1 U1078 ( .A(n2827), .B(n1222), .C(n2699), .YC(n1200), .YS(n1201) );
  FAX1 U1079 ( .A(n1207), .B(n2763), .C(n2859), .YC(n1202), .YS(n1203) );
  FAX1 U1080 ( .A(n2603), .B(n2667), .C(n2635), .YC(n1204), .YS(n1205) );
  FAX1 U1081 ( .A(n2539), .B(n2571), .C(n1224), .YC(n1206), .YS(n1207) );
  FAX1 U1082 ( .A(n1213), .B(n1228), .C(n1211), .YC(n1208), .YS(n1209) );
  FAX1 U1083 ( .A(n1232), .B(n1215), .C(n1230), .YC(n1210), .YS(n1211) );
  FAX1 U1084 ( .A(n1219), .B(n1234), .C(n1217), .YC(n1212), .YS(n1213) );
  FAX1 U1085 ( .A(n1238), .B(n1236), .C(n1221), .YC(n1214), .YS(n1215) );
  FAX1 U1086 ( .A(n2828), .B(n2796), .C(n1240), .YC(n1216), .YS(n1217) );
  FAX1 U1087 ( .A(n2860), .B(n2668), .C(n1223), .YC(n1218), .YS(n1219) );
  FAX1 U1088 ( .A(n2700), .B(n2764), .C(n2732), .YC(n1220), .YS(n1221) );
  FAX1 U1089 ( .A(n1225), .B(n2604), .C(n2636), .YC(n1222), .YS(n1223) );
  HAX1 U1090 ( .A(n2572), .B(n1242), .YC(n1224), .YS(n1225) );
  FAX1 U1091 ( .A(n1231), .B(n1246), .C(n1229), .YC(n1226), .YS(n1227) );
  FAX1 U1092 ( .A(n1250), .B(n1233), .C(n1248), .YC(n1228), .YS(n1229) );
  FAX1 U1093 ( .A(n1252), .B(n1237), .C(n1235), .YC(n1230), .YS(n1231) );
  FAX1 U1094 ( .A(n1256), .B(n1239), .C(n1254), .YC(n1232), .YS(n1233) );
  FAX1 U1095 ( .A(n2829), .B(n2797), .C(n1241), .YC(n1234), .YS(n1235) );
  FAX1 U1096 ( .A(n2861), .B(n2765), .C(n2701), .YC(n1236), .YS(n1237) );
  FAX1 U1097 ( .A(n2733), .B(n2669), .C(n1258), .YC(n1238), .YS(n1239) );
  FAX1 U1098 ( .A(n1243), .B(n2605), .C(n2637), .YC(n1240), .YS(n1241) );
  HAX1 U1099 ( .A(n2573), .B(n1260), .YC(n1242), .YS(n1243) );
  FAX1 U1100 ( .A(n1249), .B(n1264), .C(n1247), .YC(n1244), .YS(n1245) );
  FAX1 U1101 ( .A(n1268), .B(n1251), .C(n1266), .YC(n1246), .YS(n1247) );
  FAX1 U1102 ( .A(n1270), .B(n1255), .C(n1253), .YC(n1248), .YS(n1249) );
  FAX1 U1103 ( .A(n2830), .B(n1257), .C(n1272), .YC(n1250), .YS(n1251) );
  FAX1 U1104 ( .A(n2862), .B(n1274), .C(n2734), .YC(n1252), .YS(n1253) );
  FAX1 U1105 ( .A(n1259), .B(n2766), .C(n2798), .YC(n1254), .YS(n1255) );
  FAX1 U1106 ( .A(n2638), .B(n2670), .C(n2702), .YC(n1256), .YS(n1257) );
  FAX1 U1107 ( .A(n1261), .B(n2606), .C(n1276), .YC(n1258), .YS(n1259) );
  HAX1 U1108 ( .A(n5066), .B(n2574), .YC(n1260), .YS(n1261) );
  FAX1 U1109 ( .A(n1267), .B(n1280), .C(n1265), .YC(n1262), .YS(n1263) );
  FAX1 U1110 ( .A(n1284), .B(n1269), .C(n1282), .YC(n1264), .YS(n1265) );
  FAX1 U1111 ( .A(n1286), .B(n1273), .C(n1271), .YC(n1266), .YS(n1267) );
  FAX1 U1112 ( .A(n2799), .B(n1290), .C(n1288), .YC(n1268), .YS(n1269) );
  FAX1 U1113 ( .A(n2831), .B(n2703), .C(n1275), .YC(n1270), .YS(n1271) );
  FAX1 U1114 ( .A(n2735), .B(n2767), .C(n2863), .YC(n1272), .YS(n1273) );
  FAX1 U1115 ( .A(n1277), .B(n2639), .C(n2671), .YC(n1274), .YS(n1275) );
  HAX1 U1116 ( .A(n2607), .B(n1292), .YC(n1276), .YS(n1277) );
  FAX1 U1117 ( .A(n1283), .B(n1296), .C(n1281), .YC(n1278), .YS(n1279) );
  FAX1 U1118 ( .A(n1287), .B(n1285), .C(n1298), .YC(n1280), .YS(n1281) );
  FAX1 U1119 ( .A(n1289), .B(n1302), .C(n1300), .YC(n1282), .YS(n1283) );
  FAX1 U1120 ( .A(n2832), .B(n1291), .C(n1304), .YC(n1284), .YS(n1285) );
  FAX1 U1121 ( .A(n2864), .B(n2800), .C(n2736), .YC(n1286), .YS(n1287) );
  FAX1 U1122 ( .A(n2768), .B(n2704), .C(n1306), .YC(n1288), .YS(n1289) );
  FAX1 U1123 ( .A(n1293), .B(n2640), .C(n2672), .YC(n1290), .YS(n1291) );
  HAX1 U1124 ( .A(n2608), .B(n1308), .YC(n1292), .YS(n1293) );
  FAX1 U1125 ( .A(n1299), .B(n1312), .C(n1297), .YC(n1294), .YS(n1295) );
  FAX1 U1126 ( .A(n1303), .B(n1301), .C(n1314), .YC(n1296), .YS(n1297) );
  FAX1 U1127 ( .A(n1305), .B(n1318), .C(n1316), .YC(n1298), .YS(n1299) );
  FAX1 U1128 ( .A(n2833), .B(n1320), .C(n2769), .YC(n1300), .YS(n1301) );
  FAX1 U1129 ( .A(n1307), .B(n2801), .C(n2865), .YC(n1302), .YS(n1303) );
  FAX1 U1130 ( .A(n2673), .B(n2737), .C(n2705), .YC(n1304), .YS(n1305) );
  FAX1 U1131 ( .A(n1309), .B(n2641), .C(n1322), .YC(n1306), .YS(n1307) );
  HAX1 U1132 ( .A(n5063), .B(n2609), .YC(n1308), .YS(n1309) );
  FAX1 U1133 ( .A(n1315), .B(n1326), .C(n1313), .YC(n1310), .YS(n1311) );
  FAX1 U1134 ( .A(n1319), .B(n1317), .C(n1328), .YC(n1312), .YS(n1313) );
  FAX1 U1135 ( .A(n1334), .B(n1332), .C(n1330), .YC(n1314), .YS(n1315) );
  FAX1 U1136 ( .A(n2866), .B(n2738), .C(n1321), .YC(n1316), .YS(n1317) );
  FAX1 U1137 ( .A(n2770), .B(n2802), .C(n2834), .YC(n1318), .YS(n1319) );
  FAX1 U1138 ( .A(n1323), .B(n2674), .C(n2706), .YC(n1320), .YS(n1321) );
  HAX1 U1139 ( .A(n2642), .B(n1336), .YC(n1322), .YS(n1323) );
  FAX1 U1140 ( .A(n1329), .B(n1340), .C(n1327), .YC(n1324), .YS(n1325) );
  FAX1 U1141 ( .A(n1344), .B(n1331), .C(n1342), .YC(n1326), .YS(n1327) );
  FAX1 U1142 ( .A(n1335), .B(n1346), .C(n1333), .YC(n1328), .YS(n1329) );
  FAX1 U1143 ( .A(n2867), .B(n2835), .C(n2771), .YC(n1330), .YS(n1331) );
  FAX1 U1144 ( .A(n2803), .B(n2739), .C(n1348), .YC(n1332), .YS(n1333) );
  FAX1 U1145 ( .A(n1337), .B(n2675), .C(n2707), .YC(n1334), .YS(n1335) );
  HAX1 U1146 ( .A(n2643), .B(n1350), .YC(n1336), .YS(n1337) );
  FAX1 U1147 ( .A(n1343), .B(n1354), .C(n1341), .YC(n1338), .YS(n1339) );
  FAX1 U1148 ( .A(n1358), .B(n1345), .C(n1356), .YC(n1340), .YS(n1341) );
  FAX1 U1149 ( .A(n1360), .B(n2804), .C(n1347), .YC(n1342), .YS(n1343) );
  FAX1 U1150 ( .A(n1349), .B(n2868), .C(n2836), .YC(n1344), .YS(n1345) );
  FAX1 U1151 ( .A(n2708), .B(n2740), .C(n2772), .YC(n1346), .YS(n1347) );
  FAX1 U1152 ( .A(n1351), .B(n2676), .C(n1362), .YC(n1348), .YS(n1349) );
  HAX1 U1153 ( .A(n5060), .B(n2644), .YC(n1350), .YS(n1351) );
  FAX1 U1154 ( .A(n1357), .B(n1366), .C(n1355), .YC(n1352), .YS(n1353) );
  FAX1 U1155 ( .A(n1370), .B(n1359), .C(n1368), .YC(n1354), .YS(n1355) );
  FAX1 U1156 ( .A(n2773), .B(n1361), .C(n1372), .YC(n1356), .YS(n1357) );
  FAX1 U1157 ( .A(n2805), .B(n2869), .C(n2837), .YC(n1358), .YS(n1359) );
  FAX1 U1158 ( .A(n1363), .B(n2709), .C(n2741), .YC(n1360), .YS(n1361) );
  HAX1 U1159 ( .A(n2677), .B(n1374), .YC(n1362), .YS(n1363) );
  FAX1 U1160 ( .A(n1369), .B(n1378), .C(n1367), .YC(n1364), .YS(n1365) );
  FAX1 U1161 ( .A(n1382), .B(n1371), .C(n1380), .YC(n1366), .YS(n1367) );
  FAX1 U1162 ( .A(n2870), .B(n2806), .C(n1373), .YC(n1368), .YS(n1369) );
  FAX1 U1163 ( .A(n2742), .B(n2774), .C(n1384), .YC(n1370), .YS(n1371) );
  FAX1 U1164 ( .A(n1375), .B(n2710), .C(n2838), .YC(n1372), .YS(n1373) );
  HAX1 U1165 ( .A(n2678), .B(n1386), .YC(n1374), .YS(n1375) );
  FAX1 U1166 ( .A(n1381), .B(n1390), .C(n1379), .YC(n1376), .YS(n1377) );
  FAX1 U1167 ( .A(n2839), .B(n1383), .C(n1392), .YC(n1378), .YS(n1379) );
  FAX1 U1168 ( .A(n1385), .B(n2871), .C(n1394), .YC(n1380), .YS(n1381) );
  FAX1 U1169 ( .A(n2743), .B(n2807), .C(n2775), .YC(n1382), .YS(n1383) );
  FAX1 U1170 ( .A(n1387), .B(n2711), .C(n1396), .YC(n1384), .YS(n1385) );
  HAX1 U1171 ( .A(n5057), .B(n2679), .YC(n1386), .YS(n1387) );
  FAX1 U1172 ( .A(n1393), .B(n1400), .C(n1391), .YC(n1388), .YS(n1389) );
  FAX1 U1173 ( .A(n1395), .B(n1404), .C(n1402), .YC(n1390), .YS(n1391) );
  FAX1 U1174 ( .A(n2840), .B(n2872), .C(n2808), .YC(n1392), .YS(n1393) );
  FAX1 U1175 ( .A(n1397), .B(n2744), .C(n2776), .YC(n1394), .YS(n1395) );
  HAX1 U1176 ( .A(n2712), .B(n1406), .YC(n1396), .YS(n1397) );
  FAX1 U1177 ( .A(n1403), .B(n1410), .C(n1401), .YC(n1398), .YS(n1399) );
  FAX1 U1178 ( .A(n2841), .B(n1405), .C(n1412), .YC(n1400), .YS(n1401) );
  FAX1 U1179 ( .A(n2777), .B(n2809), .C(n1414), .YC(n1402), .YS(n1403) );
  FAX1 U1180 ( .A(n1407), .B(n2745), .C(n2873), .YC(n1404), .YS(n1405) );
  HAX1 U1181 ( .A(n2713), .B(n1416), .YC(n1406), .YS(n1407) );
  FAX1 U1182 ( .A(n1413), .B(n1420), .C(n1411), .YC(n1408), .YS(n1409) );
  FAX1 U1183 ( .A(n1415), .B(n1422), .C(n2874), .YC(n1410), .YS(n1411) );
  FAX1 U1184 ( .A(n2778), .B(n2842), .C(n2810), .YC(n1412), .YS(n1413) );
  FAX1 U1185 ( .A(n1417), .B(n2746), .C(n1424), .YC(n1414), .YS(n1415) );
  HAX1 U1186 ( .A(n5054), .B(n2714), .YC(n1416), .YS(n1417) );
  FAX1 U1187 ( .A(n1430), .B(n1428), .C(n1421), .YC(n1418), .YS(n1419) );
  FAX1 U1188 ( .A(n2875), .B(n2843), .C(n1423), .YC(n1420), .YS(n1421) );
  FAX1 U1189 ( .A(n1425), .B(n2779), .C(n2811), .YC(n1422), .YS(n1423) );
  HAX1 U1190 ( .A(n2747), .B(n1432), .YC(n1424), .YS(n1425) );
  FAX1 U1191 ( .A(n1431), .B(n1436), .C(n1429), .YC(n1426), .YS(n1427) );
  FAX1 U1192 ( .A(n2844), .B(n1438), .C(n2876), .YC(n1428), .YS(n1429) );
  FAX1 U1193 ( .A(n1433), .B(n2780), .C(n2812), .YC(n1430), .YS(n1431) );
  HAX1 U1194 ( .A(n2748), .B(n1440), .YC(n1432), .YS(n1433) );
  FAX1 U1195 ( .A(n1439), .B(n1444), .C(n1437), .YC(n1434), .YS(n1435) );
  FAX1 U1196 ( .A(n2813), .B(n2877), .C(n2845), .YC(n1436), .YS(n1437) );
  FAX1 U1197 ( .A(n1441), .B(n2781), .C(n1446), .YC(n1438), .YS(n1439) );
  HAX1 U1198 ( .A(n5051), .B(n2749), .YC(n1440), .YS(n1441) );
  FAX1 U1199 ( .A(n2878), .B(n1445), .C(n1450), .YC(n1442), .YS(n1443) );
  FAX1 U1200 ( .A(n1447), .B(n2814), .C(n2846), .YC(n1444), .YS(n1445) );
  HAX1 U1201 ( .A(n2782), .B(n1452), .YC(n1446), .YS(n1447) );
  FAX1 U1202 ( .A(n2879), .B(n1456), .C(n1451), .YC(n1448), .YS(n1449) );
  FAX1 U1203 ( .A(n1453), .B(n2815), .C(n2847), .YC(n1450), .YS(n1451) );
  HAX1 U1204 ( .A(n2783), .B(n1458), .YC(n1452), .YS(n1453) );
  FAX1 U1205 ( .A(n2848), .B(n2880), .C(n1457), .YC(n1454), .YS(n1455) );
  FAX1 U1206 ( .A(n1459), .B(n2816), .C(n1462), .YC(n1456), .YS(n1457) );
  HAX1 U1207 ( .A(n5048), .B(n2784), .YC(n1458), .YS(n1459) );
  FAX1 U1208 ( .A(n1463), .B(n2849), .C(n2881), .YC(n1460), .YS(n1461) );
  HAX1 U1209 ( .A(n2817), .B(n1466), .YC(n1462), .YS(n1463) );
  FAX1 U1210 ( .A(n1467), .B(n2850), .C(n2882), .YC(n1464), .YS(n1465) );
  HAX1 U1211 ( .A(n2818), .B(n1470), .YC(n1466), .YS(n1467) );
  FAX1 U1212 ( .A(n1471), .B(n2851), .C(n1472), .YC(n1468), .YS(n1469) );
  HAX1 U1213 ( .A(n5045), .B(n2819), .YC(n1470), .YS(n1471) );
  HAX1 U1214 ( .A(n2852), .B(n1474), .YC(n1472), .YS(n1473) );
  HAX1 U1215 ( .A(n2853), .B(n1476), .YC(n1474), .YS(n1475) );
  HAX1 U1216 ( .A(n5042), .B(n2854), .YC(n1476), .YS(n1477) );
  OAI21X1 U1217 ( .A(n127), .B(n3593), .C(n4443), .Y(n2516) );
  OAI21X1 U1219 ( .A(n127), .B(n4809), .C(n4526), .Y(n821) );
  AOI21X1 U1220 ( .A(n5033), .B(n129), .C(n1478), .Y(n2891) );
  AND2X1 U1221 ( .A(n124), .B(n5036), .Y(n1478) );
  OAI21X1 U1222 ( .A(n4924), .B(n4779), .C(n4317), .Y(n2517) );
  AOI21X1 U1223 ( .A(n5031), .B(n129), .C(n1480), .Y(n2892) );
  OAI21X1 U1226 ( .A(n4924), .B(n4780), .C(n4316), .Y(n2518) );
  AOI21X1 U1227 ( .A(n5029), .B(n129), .C(n1482), .Y(n2893) );
  OAI21X1 U1230 ( .A(n4924), .B(n4776), .C(n4315), .Y(n827) );
  AOI21X1 U1231 ( .A(n5027), .B(n129), .C(n1484), .Y(n2894) );
  OAI21X1 U1234 ( .A(n4924), .B(n4769), .C(n4314), .Y(n2519) );
  AOI21X1 U1235 ( .A(n5025), .B(n129), .C(n1486), .Y(n2895) );
  OAI21X1 U1238 ( .A(n4924), .B(n4778), .C(n4313), .Y(n2520) );
  AOI21X1 U1239 ( .A(n5023), .B(n129), .C(n1488), .Y(n2896) );
  OAI21X1 U1242 ( .A(n4924), .B(n3914), .C(n4312), .Y(n840) );
  AOI21X1 U1243 ( .A(n5021), .B(n129), .C(n1490), .Y(n2897) );
  OAI21X1 U1246 ( .A(n4924), .B(n4767), .C(n4311), .Y(n2521) );
  AOI21X1 U1247 ( .A(n5019), .B(n129), .C(n1492), .Y(n2898) );
  OAI21X1 U1250 ( .A(n4924), .B(n4775), .C(n4310), .Y(n2522) );
  AOI21X1 U1251 ( .A(b[22]), .B(n129), .C(n1494), .Y(n2899) );
  OAI21X1 U1254 ( .A(n127), .B(n4774), .C(n4309), .Y(n859) );
  AOI21X1 U1255 ( .A(n5017), .B(n129), .C(n1496), .Y(n2900) );
  OAI21X1 U1258 ( .A(n127), .B(n4772), .C(n4308), .Y(n2523) );
  AOI21X1 U1259 ( .A(b[20]), .B(n129), .C(n1498), .Y(n2901) );
  OAI21X1 U1262 ( .A(n4924), .B(n4804), .C(n4307), .Y(n2524) );
  AOI21X1 U1263 ( .A(n5015), .B(n129), .C(n1500), .Y(n2902) );
  OAI21X1 U1266 ( .A(n4924), .B(n4803), .C(n4306), .Y(n884) );
  AOI21X1 U1267 ( .A(n5013), .B(n129), .C(n1502), .Y(n2903) );
  OAI21X1 U1270 ( .A(n4924), .B(n4766), .C(n4305), .Y(n2525) );
  AOI21X1 U1271 ( .A(b[17]), .B(n129), .C(n1504), .Y(n2904) );
  OAI21X1 U1274 ( .A(n4924), .B(n4773), .C(n4304), .Y(n2526) );
  AOI21X1 U1275 ( .A(n5011), .B(n129), .C(n1506), .Y(n2905) );
  OAI21X1 U1278 ( .A(n4924), .B(n4768), .C(n4303), .Y(n915) );
  AOI21X1 U1279 ( .A(n5009), .B(n129), .C(n1508), .Y(n2906) );
  OAI21X1 U1282 ( .A(n4924), .B(n3923), .C(n4302), .Y(n2527) );
  AOI21X1 U1283 ( .A(n5007), .B(n129), .C(n1510), .Y(n2907) );
  OAI21X1 U1286 ( .A(n4924), .B(n4783), .C(n4301), .Y(n2528) );
  AOI21X1 U1287 ( .A(n5005), .B(n129), .C(n1512), .Y(n2908) );
  OAI21X1 U1290 ( .A(n4924), .B(n3917), .C(n4300), .Y(n952) );
  AOI21X1 U1291 ( .A(n5003), .B(n129), .C(n1514), .Y(n2909) );
  OAI21X1 U1294 ( .A(n4924), .B(n3913), .C(n4299), .Y(n2529) );
  AOI21X1 U1295 ( .A(n5001), .B(n129), .C(n1516), .Y(n2910) );
  OAI21X1 U1298 ( .A(n4924), .B(n3918), .C(n4298), .Y(n995) );
  AOI21X1 U1299 ( .A(n4999), .B(n129), .C(n1518), .Y(n2911) );
  OAI21X1 U1302 ( .A(n4924), .B(n4782), .C(n4297), .Y(n1011) );
  AOI21X1 U1303 ( .A(n4997), .B(n129), .C(n1520), .Y(n2912) );
  OAI21X1 U1306 ( .A(n4924), .B(n3916), .C(n4296), .Y(n2530) );
  AOI21X1 U1307 ( .A(n4995), .B(n129), .C(n1522), .Y(n2913) );
  OAI21X1 U1310 ( .A(n127), .B(n3921), .C(n4295), .Y(n2531) );
  AOI21X1 U1311 ( .A(n4993), .B(n129), .C(n1524), .Y(n2914) );
  OAI21X1 U1314 ( .A(n127), .B(n4784), .C(n4294), .Y(n1045) );
  AOI21X1 U1315 ( .A(n4991), .B(n129), .C(n1526), .Y(n2915) );
  OAI21X1 U1318 ( .A(n127), .B(n3920), .C(n4293), .Y(n2532) );
  AOI21X1 U1319 ( .A(n4989), .B(n129), .C(n1528), .Y(n2916) );
  OAI21X1 U1322 ( .A(n127), .B(n4802), .C(n4292), .Y(n2533) );
  AOI21X1 U1323 ( .A(n4987), .B(n129), .C(n1530), .Y(n2917) );
  OAI21X1 U1326 ( .A(n127), .B(n4801), .C(n4291), .Y(n2534) );
  AOI21X1 U1327 ( .A(n4985), .B(n129), .C(n1532), .Y(n2918) );
  OAI21X1 U1330 ( .A(n127), .B(n3922), .C(n4290), .Y(n2535) );
  AOI21X1 U1331 ( .A(b[2]), .B(n129), .C(n1534), .Y(n2919) );
  OAI21X1 U1334 ( .A(n127), .B(n3919), .C(n4289), .Y(n2536) );
  AOI21X1 U1335 ( .A(b[1]), .B(n129), .C(n1536), .Y(n2920) );
  OAI21X1 U1338 ( .A(n127), .B(n4765), .C(n4288), .Y(n2537) );
  AOI21X1 U1339 ( .A(b[0]), .B(n129), .C(n1538), .Y(n2921) );
  OAI21X1 U1342 ( .A(n127), .B(n4359), .C(n3977), .Y(n2538) );
  OAI21X1 U1344 ( .A(n127), .B(n4982), .C(n2922), .Y(n2539) );
  AND2X1 U1346 ( .A(n4928), .B(n4981), .Y(n1540) );
  XOR2X1 U1348 ( .A(n2923), .B(n5066), .Y(n2541) );
  OAI21X1 U1349 ( .A(n4929), .B(n3593), .C(n4486), .Y(n2923) );
  XOR2X1 U1351 ( .A(n2924), .B(n5066), .Y(n2542) );
  OAI21X1 U1352 ( .A(n4929), .B(n4809), .C(n4447), .Y(n2924) );
  AOI21X1 U1353 ( .A(n5033), .B(n120), .C(n1541), .Y(n2958) );
  AND2X1 U1354 ( .A(n112), .B(n5036), .Y(n1541) );
  XOR2X1 U1355 ( .A(n2925), .B(n5066), .Y(n2543) );
  OAI21X1 U1356 ( .A(n4929), .B(n4779), .C(n4287), .Y(n2925) );
  AOI21X1 U1357 ( .A(n5031), .B(n120), .C(n1543), .Y(n2959) );
  XOR2X1 U1360 ( .A(n2926), .B(n5066), .Y(n2544) );
  OAI21X1 U1361 ( .A(n4929), .B(n4780), .C(n4286), .Y(n2926) );
  AOI21X1 U1362 ( .A(n5029), .B(n120), .C(n1545), .Y(n2960) );
  XOR2X1 U1365 ( .A(n2927), .B(n5066), .Y(n2545) );
  OAI21X1 U1366 ( .A(n4929), .B(n4776), .C(n4285), .Y(n2927) );
  AOI21X1 U1367 ( .A(n5027), .B(n120), .C(n1547), .Y(n2961) );
  XOR2X1 U1370 ( .A(n2928), .B(n5066), .Y(n2546) );
  OAI21X1 U1371 ( .A(n4929), .B(n4769), .C(n4284), .Y(n2928) );
  AOI21X1 U1372 ( .A(n5025), .B(n120), .C(n1549), .Y(n2962) );
  XOR2X1 U1375 ( .A(n2929), .B(n5066), .Y(n2547) );
  OAI21X1 U1376 ( .A(n4929), .B(n4778), .C(n4283), .Y(n2929) );
  AOI21X1 U1377 ( .A(n5023), .B(n120), .C(n1551), .Y(n2963) );
  XOR2X1 U1380 ( .A(n2930), .B(n5067), .Y(n2548) );
  OAI21X1 U1381 ( .A(n4929), .B(n3914), .C(n4282), .Y(n2930) );
  AOI21X1 U1382 ( .A(n5021), .B(n120), .C(n1553), .Y(n2964) );
  XOR2X1 U1385 ( .A(n2931), .B(n5066), .Y(n2549) );
  OAI21X1 U1386 ( .A(n4929), .B(n4767), .C(n4281), .Y(n2931) );
  AOI21X1 U1387 ( .A(n5019), .B(n120), .C(n1555), .Y(n2965) );
  XOR2X1 U1390 ( .A(n2932), .B(n5066), .Y(n2550) );
  OAI21X1 U1391 ( .A(n4929), .B(n4775), .C(n4280), .Y(n2932) );
  AOI21X1 U1392 ( .A(b[22]), .B(n120), .C(n1557), .Y(n2966) );
  XOR2X1 U1395 ( .A(n2933), .B(n5066), .Y(n2551) );
  OAI21X1 U1396 ( .A(n118), .B(n4774), .C(n4279), .Y(n2933) );
  AOI21X1 U1397 ( .A(n5017), .B(n120), .C(n1559), .Y(n2967) );
  XOR2X1 U1400 ( .A(n2934), .B(n5067), .Y(n2552) );
  OAI21X1 U1401 ( .A(n118), .B(n4772), .C(n4278), .Y(n2934) );
  AOI21X1 U1402 ( .A(b[20]), .B(n120), .C(n1561), .Y(n2968) );
  XOR2X1 U1405 ( .A(n2935), .B(a[29]), .Y(n2553) );
  OAI21X1 U1406 ( .A(n4929), .B(n4804), .C(n4277), .Y(n2935) );
  AOI21X1 U1407 ( .A(n5015), .B(n120), .C(n1563), .Y(n2969) );
  XOR2X1 U1410 ( .A(n2936), .B(a[29]), .Y(n2554) );
  OAI21X1 U1411 ( .A(n4929), .B(n4803), .C(n4276), .Y(n2936) );
  AOI21X1 U1412 ( .A(n5013), .B(n120), .C(n1565), .Y(n2970) );
  XOR2X1 U1415 ( .A(n2937), .B(n5066), .Y(n2555) );
  OAI21X1 U1416 ( .A(n4929), .B(n4766), .C(n4275), .Y(n2937) );
  AOI21X1 U1417 ( .A(b[17]), .B(n120), .C(n1567), .Y(n2971) );
  XOR2X1 U1420 ( .A(n2938), .B(n5066), .Y(n2556) );
  OAI21X1 U1421 ( .A(n4929), .B(n4773), .C(n4274), .Y(n2938) );
  AOI21X1 U1422 ( .A(n5011), .B(n120), .C(n1569), .Y(n2972) );
  XOR2X1 U1425 ( .A(n2939), .B(n5066), .Y(n2557) );
  OAI21X1 U1426 ( .A(n4929), .B(n4768), .C(n4273), .Y(n2939) );
  AOI21X1 U1427 ( .A(b[15]), .B(n120), .C(n1571), .Y(n2973) );
  XOR2X1 U1430 ( .A(n2940), .B(n5066), .Y(n2558) );
  OAI21X1 U1431 ( .A(n4929), .B(n3923), .C(n4272), .Y(n2940) );
  AOI21X1 U1432 ( .A(n5007), .B(n120), .C(n1573), .Y(n2974) );
  XOR2X1 U1435 ( .A(n2941), .B(n5066), .Y(n2559) );
  OAI21X1 U1436 ( .A(n4929), .B(n4783), .C(n4271), .Y(n2941) );
  AOI21X1 U1437 ( .A(n5005), .B(n120), .C(n1575), .Y(n2975) );
  XOR2X1 U1440 ( .A(n2942), .B(n5067), .Y(n2560) );
  OAI21X1 U1441 ( .A(n4929), .B(n3917), .C(n4270), .Y(n2942) );
  AOI21X1 U1442 ( .A(n5003), .B(n120), .C(n1577), .Y(n2976) );
  XOR2X1 U1445 ( .A(n2943), .B(n5067), .Y(n2561) );
  OAI21X1 U1446 ( .A(n4929), .B(n3913), .C(n4269), .Y(n2943) );
  AOI21X1 U1447 ( .A(n5001), .B(n120), .C(n1579), .Y(n2977) );
  XOR2X1 U1450 ( .A(n2944), .B(n5067), .Y(n2562) );
  OAI21X1 U1451 ( .A(n4929), .B(n3918), .C(n4268), .Y(n2944) );
  AOI21X1 U1452 ( .A(n4999), .B(n120), .C(n1581), .Y(n2978) );
  XOR2X1 U1455 ( .A(n2945), .B(n5066), .Y(n2563) );
  OAI21X1 U1456 ( .A(n4929), .B(n4782), .C(n4267), .Y(n2945) );
  AOI21X1 U1457 ( .A(n4997), .B(n120), .C(n1583), .Y(n2979) );
  XOR2X1 U1460 ( .A(n2946), .B(n5066), .Y(n2564) );
  OAI21X1 U1461 ( .A(n4929), .B(n3916), .C(n4266), .Y(n2946) );
  AOI21X1 U1462 ( .A(n4995), .B(n120), .C(n1585), .Y(n2980) );
  XOR2X1 U1465 ( .A(n2947), .B(n5066), .Y(n2565) );
  OAI21X1 U1466 ( .A(n118), .B(n3921), .C(n4265), .Y(n2947) );
  AOI21X1 U1467 ( .A(n4993), .B(n120), .C(n1587), .Y(n2981) );
  XOR2X1 U1470 ( .A(n2948), .B(n5067), .Y(n2566) );
  OAI21X1 U1471 ( .A(n118), .B(n4784), .C(n4264), .Y(n2948) );
  AOI21X1 U1472 ( .A(n4991), .B(n120), .C(n1589), .Y(n2982) );
  XOR2X1 U1475 ( .A(n2949), .B(n5067), .Y(n2567) );
  OAI21X1 U1476 ( .A(n118), .B(n3920), .C(n4263), .Y(n2949) );
  AOI21X1 U1477 ( .A(n4989), .B(n120), .C(n1591), .Y(n2983) );
  XOR2X1 U1480 ( .A(n2950), .B(n5067), .Y(n2568) );
  OAI21X1 U1481 ( .A(n118), .B(n4802), .C(n4262), .Y(n2950) );
  AOI21X1 U1482 ( .A(n4987), .B(n120), .C(n1593), .Y(n2984) );
  XOR2X1 U1485 ( .A(n2951), .B(n5067), .Y(n2569) );
  OAI21X1 U1486 ( .A(n118), .B(n4801), .C(n4261), .Y(n2951) );
  AOI21X1 U1487 ( .A(b[3]), .B(n120), .C(n1595), .Y(n2985) );
  XOR2X1 U1490 ( .A(n2952), .B(n5067), .Y(n2570) );
  OAI21X1 U1491 ( .A(n118), .B(n3922), .C(n4260), .Y(n2952) );
  AOI21X1 U1492 ( .A(b[2]), .B(n120), .C(n1597), .Y(n2986) );
  XOR2X1 U1495 ( .A(n2953), .B(n5067), .Y(n2571) );
  OAI21X1 U1496 ( .A(n118), .B(n3919), .C(n4259), .Y(n2953) );
  AOI21X1 U1497 ( .A(b[1]), .B(n120), .C(n1599), .Y(n2987) );
  XOR2X1 U1500 ( .A(n2954), .B(n5067), .Y(n2572) );
  OAI21X1 U1501 ( .A(n118), .B(n4765), .C(n4258), .Y(n2954) );
  AOI21X1 U1502 ( .A(n4981), .B(n120), .C(n1601), .Y(n2988) );
  XOR2X1 U1505 ( .A(n2955), .B(n5067), .Y(n2573) );
  OAI21X1 U1506 ( .A(n118), .B(n4359), .C(n3976), .Y(n2955) );
  XOR2X1 U1508 ( .A(n2956), .B(n5067), .Y(n2574) );
  OAI21X1 U1509 ( .A(n118), .B(n4982), .C(n2989), .Y(n2956) );
  AND2X1 U1511 ( .A(n4932), .B(n4981), .Y(n1603) );
  XOR2X1 U1513 ( .A(n2990), .B(n5063), .Y(n2576) );
  OAI21X1 U1514 ( .A(n4933), .B(n3593), .C(n4704), .Y(n2990) );
  XOR2X1 U1516 ( .A(n2991), .B(n5063), .Y(n2577) );
  OAI21X1 U1517 ( .A(n4933), .B(n4809), .C(n4257), .Y(n2991) );
  AOI21X1 U1518 ( .A(n5033), .B(n108), .C(n1604), .Y(n3025) );
  AND2X1 U1519 ( .A(n100), .B(n5036), .Y(n1604) );
  XOR2X1 U1520 ( .A(n2992), .B(n5063), .Y(n2578) );
  OAI21X1 U1521 ( .A(n4933), .B(n4779), .C(n4256), .Y(n2992) );
  AOI21X1 U1522 ( .A(n5031), .B(n108), .C(n1606), .Y(n3026) );
  XOR2X1 U1525 ( .A(n2993), .B(n5063), .Y(n2579) );
  OAI21X1 U1526 ( .A(n4933), .B(n4780), .C(n4255), .Y(n2993) );
  AOI21X1 U1527 ( .A(n5029), .B(n108), .C(n1608), .Y(n3027) );
  XOR2X1 U1530 ( .A(n2994), .B(n5063), .Y(n2580) );
  OAI21X1 U1531 ( .A(n4933), .B(n4776), .C(n4254), .Y(n2994) );
  AOI21X1 U1532 ( .A(n5027), .B(n108), .C(n1610), .Y(n3028) );
  XOR2X1 U1535 ( .A(n2995), .B(n5063), .Y(n2581) );
  OAI21X1 U1536 ( .A(n4933), .B(n4769), .C(n4253), .Y(n2995) );
  AOI21X1 U1537 ( .A(n5025), .B(n108), .C(n1612), .Y(n3029) );
  XOR2X1 U1540 ( .A(n2996), .B(n5063), .Y(n2582) );
  OAI21X1 U1541 ( .A(n4933), .B(n4778), .C(n4252), .Y(n2996) );
  AOI21X1 U1542 ( .A(n5023), .B(n108), .C(n1614), .Y(n3030) );
  XOR2X1 U1545 ( .A(n2997), .B(n5064), .Y(n2583) );
  OAI21X1 U1546 ( .A(n4933), .B(n3914), .C(n4251), .Y(n2997) );
  AOI21X1 U1547 ( .A(n5021), .B(n108), .C(n1616), .Y(n3031) );
  XOR2X1 U1550 ( .A(n2998), .B(n5063), .Y(n2584) );
  OAI21X1 U1551 ( .A(n4933), .B(n4767), .C(n4250), .Y(n2998) );
  AOI21X1 U1552 ( .A(n5019), .B(n108), .C(n1618), .Y(n3032) );
  XOR2X1 U1555 ( .A(n2999), .B(n5063), .Y(n2585) );
  OAI21X1 U1556 ( .A(n4933), .B(n4775), .C(n4249), .Y(n2999) );
  AOI21X1 U1557 ( .A(b[22]), .B(n108), .C(n1620), .Y(n3033) );
  XOR2X1 U1560 ( .A(n3000), .B(n5063), .Y(n2586) );
  OAI21X1 U1561 ( .A(n106), .B(n4774), .C(n4248), .Y(n3000) );
  AOI21X1 U1562 ( .A(n5017), .B(n108), .C(n1622), .Y(n3034) );
  XOR2X1 U1565 ( .A(n3001), .B(n5063), .Y(n2587) );
  OAI21X1 U1566 ( .A(n106), .B(n4772), .C(n4247), .Y(n3001) );
  AOI21X1 U1567 ( .A(b[20]), .B(n108), .C(n1624), .Y(n3035) );
  XOR2X1 U1570 ( .A(n3002), .B(n5063), .Y(n2588) );
  OAI21X1 U1571 ( .A(n4933), .B(n4804), .C(n4246), .Y(n3002) );
  AOI21X1 U1572 ( .A(n5015), .B(n108), .C(n1626), .Y(n3036) );
  XOR2X1 U1575 ( .A(n3003), .B(n5063), .Y(n2589) );
  OAI21X1 U1576 ( .A(n4933), .B(n4803), .C(n4245), .Y(n3003) );
  AOI21X1 U1577 ( .A(n5013), .B(n108), .C(n1628), .Y(n3037) );
  XOR2X1 U1580 ( .A(n3004), .B(n5064), .Y(n2590) );
  OAI21X1 U1581 ( .A(n4933), .B(n4766), .C(n4244), .Y(n3004) );
  AOI21X1 U1582 ( .A(b[17]), .B(n108), .C(n1630), .Y(n3038) );
  XOR2X1 U1585 ( .A(n3005), .B(n5063), .Y(n2591) );
  OAI21X1 U1586 ( .A(n4933), .B(n4773), .C(n4243), .Y(n3005) );
  AOI21X1 U1587 ( .A(n5011), .B(n108), .C(n1632), .Y(n3039) );
  XOR2X1 U1590 ( .A(n3006), .B(n5063), .Y(n2592) );
  OAI21X1 U1591 ( .A(n4933), .B(n4768), .C(n4242), .Y(n3006) );
  AOI21X1 U1592 ( .A(n5009), .B(n108), .C(n1634), .Y(n3040) );
  XOR2X1 U1595 ( .A(n3007), .B(n5063), .Y(n2593) );
  OAI21X1 U1596 ( .A(n4933), .B(n3923), .C(n4241), .Y(n3007) );
  AOI21X1 U1597 ( .A(n5007), .B(n108), .C(n1636), .Y(n3041) );
  XOR2X1 U1600 ( .A(n3008), .B(n5064), .Y(n2594) );
  OAI21X1 U1601 ( .A(n4933), .B(n4783), .C(n4240), .Y(n3008) );
  AOI21X1 U1602 ( .A(n5005), .B(n108), .C(n1638), .Y(n3042) );
  XOR2X1 U1605 ( .A(n3009), .B(n5064), .Y(n2595) );
  OAI21X1 U1606 ( .A(n4933), .B(n3917), .C(n4239), .Y(n3009) );
  AOI21X1 U1607 ( .A(n5003), .B(n108), .C(n1640), .Y(n3043) );
  XOR2X1 U1610 ( .A(n3010), .B(n5064), .Y(n2596) );
  OAI21X1 U1611 ( .A(n4933), .B(n3913), .C(n4238), .Y(n3010) );
  AOI21X1 U1612 ( .A(n5001), .B(n108), .C(n1642), .Y(n3044) );
  XOR2X1 U1615 ( .A(n3011), .B(n5064), .Y(n2597) );
  OAI21X1 U1616 ( .A(n4933), .B(n3918), .C(n4237), .Y(n3011) );
  AOI21X1 U1617 ( .A(n4999), .B(n108), .C(n1644), .Y(n3045) );
  XOR2X1 U1620 ( .A(n3012), .B(n5063), .Y(n2598) );
  OAI21X1 U1621 ( .A(n4933), .B(n4782), .C(n4236), .Y(n3012) );
  AOI21X1 U1622 ( .A(n4997), .B(n108), .C(n1646), .Y(n3046) );
  XOR2X1 U1625 ( .A(n3013), .B(n5063), .Y(n2599) );
  OAI21X1 U1626 ( .A(n4933), .B(n3916), .C(n4235), .Y(n3013) );
  AOI21X1 U1627 ( .A(n4995), .B(n108), .C(n1648), .Y(n3047) );
  XOR2X1 U1630 ( .A(n3014), .B(n5063), .Y(n2600) );
  OAI21X1 U1631 ( .A(n106), .B(n3921), .C(n4234), .Y(n3014) );
  AOI21X1 U1632 ( .A(n4993), .B(n108), .C(n1650), .Y(n3048) );
  XOR2X1 U1635 ( .A(n3015), .B(n5064), .Y(n2601) );
  OAI21X1 U1636 ( .A(n106), .B(n4784), .C(n4233), .Y(n3015) );
  AOI21X1 U1637 ( .A(n4991), .B(n108), .C(n1652), .Y(n3049) );
  XOR2X1 U1640 ( .A(n3016), .B(n5064), .Y(n2602) );
  OAI21X1 U1641 ( .A(n106), .B(n3920), .C(n4232), .Y(n3016) );
  AOI21X1 U1642 ( .A(n4989), .B(n108), .C(n1654), .Y(n3050) );
  XOR2X1 U1645 ( .A(n3017), .B(n5064), .Y(n2603) );
  OAI21X1 U1646 ( .A(n106), .B(n4802), .C(n4231), .Y(n3017) );
  AOI21X1 U1647 ( .A(n4987), .B(n108), .C(n1656), .Y(n3051) );
  XOR2X1 U1650 ( .A(n3018), .B(n5064), .Y(n2604) );
  OAI21X1 U1651 ( .A(n106), .B(n4801), .C(n4230), .Y(n3018) );
  AOI21X1 U1652 ( .A(b[3]), .B(n108), .C(n1658), .Y(n3052) );
  XOR2X1 U1655 ( .A(n3019), .B(n5064), .Y(n2605) );
  OAI21X1 U1656 ( .A(n106), .B(n3922), .C(n4229), .Y(n3019) );
  AOI21X1 U1657 ( .A(b[2]), .B(n108), .C(n1660), .Y(n3053) );
  XOR2X1 U1660 ( .A(n3020), .B(n5064), .Y(n2606) );
  OAI21X1 U1661 ( .A(n106), .B(n3919), .C(n4228), .Y(n3020) );
  AOI21X1 U1662 ( .A(b[1]), .B(n108), .C(n1662), .Y(n3054) );
  XOR2X1 U1665 ( .A(n3021), .B(n5064), .Y(n2607) );
  OAI21X1 U1666 ( .A(n106), .B(n4765), .C(n4227), .Y(n3021) );
  AOI21X1 U1667 ( .A(b[0]), .B(n108), .C(n1664), .Y(n3055) );
  XOR2X1 U1670 ( .A(n3022), .B(n5064), .Y(n2608) );
  OAI21X1 U1671 ( .A(n106), .B(n4359), .C(n3975), .Y(n3022) );
  XOR2X1 U1673 ( .A(n3023), .B(n5064), .Y(n2609) );
  OAI21X1 U1674 ( .A(n106), .B(n4982), .C(n3056), .Y(n3023) );
  AND2X1 U1676 ( .A(n4935), .B(n4981), .Y(n1666) );
  XOR2X1 U1678 ( .A(n3057), .B(n5060), .Y(n2611) );
  OAI21X1 U1679 ( .A(n4936), .B(n3593), .C(n4444), .Y(n3057) );
  XOR2X1 U1681 ( .A(n3058), .B(n5060), .Y(n2612) );
  OAI21X1 U1682 ( .A(n4936), .B(n4809), .C(n4488), .Y(n3058) );
  AOI21X1 U1683 ( .A(n5033), .B(n96), .C(n1667), .Y(n3092) );
  AND2X1 U1684 ( .A(n88), .B(n5036), .Y(n1667) );
  XOR2X1 U1685 ( .A(n3059), .B(n5060), .Y(n2613) );
  OAI21X1 U1686 ( .A(n4936), .B(n4779), .C(n4226), .Y(n3059) );
  AOI21X1 U1687 ( .A(n5031), .B(n96), .C(n1669), .Y(n3093) );
  XOR2X1 U1690 ( .A(n3060), .B(n5060), .Y(n2614) );
  OAI21X1 U1691 ( .A(n4936), .B(n4780), .C(n4225), .Y(n3060) );
  AOI21X1 U1692 ( .A(n5029), .B(n96), .C(n1671), .Y(n3094) );
  XOR2X1 U1695 ( .A(n3061), .B(n5060), .Y(n2615) );
  OAI21X1 U1696 ( .A(n4936), .B(n4776), .C(n4224), .Y(n3061) );
  AOI21X1 U1697 ( .A(n5027), .B(n96), .C(n1673), .Y(n3095) );
  XOR2X1 U1700 ( .A(n3062), .B(n5060), .Y(n2616) );
  OAI21X1 U1701 ( .A(n4936), .B(n4769), .C(n4223), .Y(n3062) );
  AOI21X1 U1702 ( .A(n5025), .B(n96), .C(n1675), .Y(n3096) );
  XOR2X1 U1705 ( .A(n3063), .B(n5060), .Y(n2617) );
  OAI21X1 U1706 ( .A(n4936), .B(n4778), .C(n4222), .Y(n3063) );
  AOI21X1 U1707 ( .A(n5023), .B(n96), .C(n1677), .Y(n3097) );
  XOR2X1 U1710 ( .A(n3064), .B(n5061), .Y(n2618) );
  OAI21X1 U1711 ( .A(n4936), .B(n3914), .C(n4221), .Y(n3064) );
  AOI21X1 U1712 ( .A(n5021), .B(n96), .C(n1679), .Y(n3098) );
  XOR2X1 U1715 ( .A(n3065), .B(n5060), .Y(n2619) );
  OAI21X1 U1716 ( .A(n4936), .B(n4767), .C(n4220), .Y(n3065) );
  AOI21X1 U1717 ( .A(n5019), .B(n96), .C(n1681), .Y(n3099) );
  XOR2X1 U1720 ( .A(n3066), .B(n5060), .Y(n2620) );
  OAI21X1 U1721 ( .A(n4936), .B(n4775), .C(n4219), .Y(n3066) );
  AOI21X1 U1722 ( .A(b[22]), .B(n96), .C(n1683), .Y(n3100) );
  XOR2X1 U1725 ( .A(n3067), .B(n5060), .Y(n2621) );
  OAI21X1 U1726 ( .A(n94), .B(n4774), .C(n4218), .Y(n3067) );
  AOI21X1 U1727 ( .A(n5017), .B(n96), .C(n1685), .Y(n3101) );
  XOR2X1 U1730 ( .A(n3068), .B(n5060), .Y(n2622) );
  OAI21X1 U1731 ( .A(n94), .B(n4772), .C(n4217), .Y(n3068) );
  AOI21X1 U1732 ( .A(b[20]), .B(n96), .C(n1687), .Y(n3102) );
  XOR2X1 U1735 ( .A(n3069), .B(n5060), .Y(n2623) );
  OAI21X1 U1736 ( .A(n4936), .B(n4804), .C(n4216), .Y(n3069) );
  AOI21X1 U1737 ( .A(n5015), .B(n96), .C(n1689), .Y(n3103) );
  XOR2X1 U1740 ( .A(n3070), .B(n5060), .Y(n2624) );
  OAI21X1 U1741 ( .A(n4936), .B(n4803), .C(n4215), .Y(n3070) );
  AOI21X1 U1742 ( .A(n5013), .B(n96), .C(n1691), .Y(n3104) );
  XOR2X1 U1745 ( .A(n3071), .B(n5061), .Y(n2625) );
  OAI21X1 U1746 ( .A(n4936), .B(n4766), .C(n4214), .Y(n3071) );
  AOI21X1 U1747 ( .A(b[17]), .B(n96), .C(n1693), .Y(n3105) );
  XOR2X1 U1750 ( .A(n3072), .B(n5060), .Y(n2626) );
  OAI21X1 U1751 ( .A(n4936), .B(n4773), .C(n4213), .Y(n3072) );
  AOI21X1 U1752 ( .A(n5011), .B(n96), .C(n1695), .Y(n3106) );
  XOR2X1 U1755 ( .A(n3073), .B(n5061), .Y(n2627) );
  OAI21X1 U1756 ( .A(n4936), .B(n4768), .C(n4212), .Y(n3073) );
  AOI21X1 U1757 ( .A(n5009), .B(n96), .C(n1697), .Y(n3107) );
  XOR2X1 U1760 ( .A(n3074), .B(n5060), .Y(n2628) );
  OAI21X1 U1761 ( .A(n4936), .B(n3923), .C(n4211), .Y(n3074) );
  AOI21X1 U1762 ( .A(n5007), .B(n96), .C(n1699), .Y(n3108) );
  XOR2X1 U1765 ( .A(n3075), .B(n5060), .Y(n2629) );
  OAI21X1 U1766 ( .A(n4936), .B(n4783), .C(n4210), .Y(n3075) );
  AOI21X1 U1767 ( .A(n5005), .B(n96), .C(n1701), .Y(n3109) );
  XOR2X1 U1770 ( .A(n3076), .B(n5061), .Y(n2630) );
  OAI21X1 U1771 ( .A(n4936), .B(n3917), .C(n4209), .Y(n3076) );
  AOI21X1 U1772 ( .A(n5003), .B(n96), .C(n1703), .Y(n3110) );
  XOR2X1 U1775 ( .A(n3077), .B(n5061), .Y(n2631) );
  OAI21X1 U1776 ( .A(n4936), .B(n3913), .C(n4208), .Y(n3077) );
  AOI21X1 U1777 ( .A(n5001), .B(n96), .C(n1705), .Y(n3111) );
  XOR2X1 U1780 ( .A(n3078), .B(n5061), .Y(n2632) );
  OAI21X1 U1781 ( .A(n4936), .B(n3918), .C(n4207), .Y(n3078) );
  AOI21X1 U1782 ( .A(n4999), .B(n96), .C(n1707), .Y(n3112) );
  XOR2X1 U1785 ( .A(n3079), .B(n5060), .Y(n2633) );
  OAI21X1 U1786 ( .A(n4936), .B(n4782), .C(n4206), .Y(n3079) );
  AOI21X1 U1787 ( .A(n4997), .B(n96), .C(n1709), .Y(n3113) );
  XOR2X1 U1790 ( .A(n3080), .B(n5060), .Y(n2634) );
  OAI21X1 U1791 ( .A(n4936), .B(n3916), .C(n4205), .Y(n3080) );
  AOI21X1 U1792 ( .A(n4995), .B(n96), .C(n1711), .Y(n3114) );
  XOR2X1 U1795 ( .A(n3081), .B(n5060), .Y(n2635) );
  OAI21X1 U1796 ( .A(n94), .B(n3921), .C(n4204), .Y(n3081) );
  AOI21X1 U1797 ( .A(n4993), .B(n96), .C(n1713), .Y(n3115) );
  XOR2X1 U1800 ( .A(n3082), .B(n5061), .Y(n2636) );
  OAI21X1 U1801 ( .A(n94), .B(n4784), .C(n4203), .Y(n3082) );
  AOI21X1 U1802 ( .A(n4991), .B(n96), .C(n1715), .Y(n3116) );
  XOR2X1 U1805 ( .A(n3083), .B(n5061), .Y(n2637) );
  OAI21X1 U1806 ( .A(n94), .B(n3920), .C(n4202), .Y(n3083) );
  AOI21X1 U1807 ( .A(n4989), .B(n96), .C(n1717), .Y(n3117) );
  XOR2X1 U1810 ( .A(n3084), .B(n5061), .Y(n2638) );
  OAI21X1 U1811 ( .A(n94), .B(n4802), .C(n4201), .Y(n3084) );
  AOI21X1 U1812 ( .A(n4987), .B(n96), .C(n1719), .Y(n3118) );
  XOR2X1 U1815 ( .A(n3085), .B(n5061), .Y(n2639) );
  OAI21X1 U1816 ( .A(n94), .B(n4801), .C(n4200), .Y(n3085) );
  AOI21X1 U1817 ( .A(b[3]), .B(n96), .C(n1721), .Y(n3119) );
  XOR2X1 U1820 ( .A(n3086), .B(n5061), .Y(n2640) );
  OAI21X1 U1821 ( .A(n94), .B(n3922), .C(n4199), .Y(n3086) );
  AOI21X1 U1822 ( .A(b[2]), .B(n96), .C(n1723), .Y(n3120) );
  XOR2X1 U1825 ( .A(n3087), .B(n5061), .Y(n2641) );
  OAI21X1 U1826 ( .A(n94), .B(n3919), .C(n4198), .Y(n3087) );
  AOI21X1 U1827 ( .A(b[1]), .B(n96), .C(n1725), .Y(n3121) );
  XOR2X1 U1830 ( .A(n3088), .B(n5061), .Y(n2642) );
  OAI21X1 U1831 ( .A(n94), .B(n4765), .C(n4197), .Y(n3088) );
  AOI21X1 U1832 ( .A(b[0]), .B(n96), .C(n1727), .Y(n3122) );
  XOR2X1 U1835 ( .A(n3089), .B(n5061), .Y(n2643) );
  OAI21X1 U1836 ( .A(n94), .B(n4359), .C(n3974), .Y(n3089) );
  XOR2X1 U1838 ( .A(n3090), .B(n5061), .Y(n2644) );
  OAI21X1 U1839 ( .A(n94), .B(n4982), .C(n3123), .Y(n3090) );
  AND2X1 U1841 ( .A(n4938), .B(n4981), .Y(n1729) );
  XOR2X1 U1843 ( .A(n3124), .B(n5057), .Y(n2646) );
  OAI21X1 U1844 ( .A(n4939), .B(n3593), .C(n4446), .Y(n3124) );
  XOR2X1 U1846 ( .A(n3125), .B(n5057), .Y(n2647) );
  OAI21X1 U1847 ( .A(n4939), .B(n4809), .C(n4445), .Y(n3125) );
  AOI21X1 U1848 ( .A(n5033), .B(n84), .C(n1730), .Y(n3159) );
  AND2X1 U1849 ( .A(n76), .B(n5036), .Y(n1730) );
  XOR2X1 U1850 ( .A(n3126), .B(n5057), .Y(n2648) );
  OAI21X1 U1851 ( .A(n4779), .B(n4939), .C(n4196), .Y(n3126) );
  AOI21X1 U1852 ( .A(n5031), .B(n84), .C(n1732), .Y(n3160) );
  XOR2X1 U1855 ( .A(n3127), .B(n5057), .Y(n2649) );
  OAI21X1 U1856 ( .A(n4939), .B(n4780), .C(n4195), .Y(n3127) );
  AOI21X1 U1857 ( .A(n5029), .B(n84), .C(n1734), .Y(n3161) );
  XOR2X1 U1860 ( .A(n3128), .B(n5057), .Y(n2650) );
  OAI21X1 U1861 ( .A(n4939), .B(n4776), .C(n4194), .Y(n3128) );
  AOI21X1 U1862 ( .A(n5027), .B(n84), .C(n1736), .Y(n3162) );
  XOR2X1 U1865 ( .A(n3129), .B(n5057), .Y(n2651) );
  OAI21X1 U1866 ( .A(n4939), .B(n4769), .C(n4193), .Y(n3129) );
  AOI21X1 U1867 ( .A(n5025), .B(n84), .C(n1738), .Y(n3163) );
  XOR2X1 U1870 ( .A(n3130), .B(n5057), .Y(n2652) );
  OAI21X1 U1871 ( .A(n4939), .B(n4778), .C(n4192), .Y(n3130) );
  AOI21X1 U1872 ( .A(n5023), .B(n84), .C(n1740), .Y(n3164) );
  XOR2X1 U1875 ( .A(n3131), .B(n5058), .Y(n2653) );
  OAI21X1 U1876 ( .A(n4939), .B(n3914), .C(n4191), .Y(n3131) );
  AOI21X1 U1877 ( .A(n5021), .B(n84), .C(n1742), .Y(n3165) );
  XOR2X1 U1880 ( .A(n3132), .B(n5057), .Y(n2654) );
  OAI21X1 U1881 ( .A(n4939), .B(n4767), .C(n4190), .Y(n3132) );
  AOI21X1 U1882 ( .A(n5019), .B(n84), .C(n1744), .Y(n3166) );
  XOR2X1 U1885 ( .A(n3133), .B(n5057), .Y(n2655) );
  OAI21X1 U1886 ( .A(n4939), .B(n4775), .C(n4189), .Y(n3133) );
  AOI21X1 U1887 ( .A(b[22]), .B(n84), .C(n1746), .Y(n3167) );
  XOR2X1 U1890 ( .A(n3134), .B(n5057), .Y(n2656) );
  OAI21X1 U1891 ( .A(n82), .B(n4774), .C(n4188), .Y(n3134) );
  AOI21X1 U1892 ( .A(n5017), .B(n84), .C(n1748), .Y(n3168) );
  XOR2X1 U1895 ( .A(n3135), .B(n5058), .Y(n2657) );
  OAI21X1 U1896 ( .A(n82), .B(n4772), .C(n4187), .Y(n3135) );
  AOI21X1 U1897 ( .A(b[20]), .B(n84), .C(n1750), .Y(n3169) );
  XOR2X1 U1900 ( .A(n3136), .B(a[20]), .Y(n2658) );
  OAI21X1 U1901 ( .A(n4939), .B(n4804), .C(n4186), .Y(n3136) );
  AOI21X1 U1902 ( .A(n5015), .B(n84), .C(n1752), .Y(n3170) );
  XOR2X1 U1905 ( .A(n3137), .B(n5057), .Y(n2659) );
  OAI21X1 U1906 ( .A(n4939), .B(n4803), .C(n4185), .Y(n3137) );
  AOI21X1 U1907 ( .A(n5013), .B(n84), .C(n1754), .Y(n3171) );
  XOR2X1 U1910 ( .A(n3138), .B(n5058), .Y(n2660) );
  OAI21X1 U1911 ( .A(n4939), .B(n4766), .C(n4184), .Y(n3138) );
  AOI21X1 U1912 ( .A(b[17]), .B(n84), .C(n1756), .Y(n3172) );
  XOR2X1 U1915 ( .A(n3139), .B(a[20]), .Y(n2661) );
  OAI21X1 U1916 ( .A(n4939), .B(n4773), .C(n4183), .Y(n3139) );
  AOI21X1 U1917 ( .A(n5011), .B(n84), .C(n1758), .Y(n3173) );
  XOR2X1 U1920 ( .A(n3140), .B(n5057), .Y(n2662) );
  OAI21X1 U1921 ( .A(n4939), .B(n4768), .C(n4182), .Y(n3140) );
  AOI21X1 U1922 ( .A(n5009), .B(n84), .C(n1760), .Y(n3174) );
  XOR2X1 U1925 ( .A(n3141), .B(n5057), .Y(n2663) );
  OAI21X1 U1926 ( .A(n4939), .B(n3923), .C(n4181), .Y(n3141) );
  AOI21X1 U1927 ( .A(n5007), .B(n84), .C(n1762), .Y(n3175) );
  XOR2X1 U1930 ( .A(n3142), .B(n5057), .Y(n2664) );
  OAI21X1 U1931 ( .A(n4939), .B(n4783), .C(n4180), .Y(n3142) );
  AOI21X1 U1932 ( .A(n5005), .B(n84), .C(n1764), .Y(n3176) );
  XOR2X1 U1935 ( .A(n3143), .B(n5058), .Y(n2665) );
  OAI21X1 U1936 ( .A(n4939), .B(n3917), .C(n4179), .Y(n3143) );
  AOI21X1 U1937 ( .A(n5003), .B(n84), .C(n1766), .Y(n3177) );
  XOR2X1 U1940 ( .A(n3144), .B(n5058), .Y(n2666) );
  OAI21X1 U1941 ( .A(n4939), .B(n3913), .C(n4178), .Y(n3144) );
  AOI21X1 U1942 ( .A(n5001), .B(n84), .C(n1768), .Y(n3178) );
  XOR2X1 U1945 ( .A(n3145), .B(n5058), .Y(n2667) );
  OAI21X1 U1946 ( .A(n4939), .B(n3918), .C(n4177), .Y(n3145) );
  AOI21X1 U1947 ( .A(n4999), .B(n84), .C(n1770), .Y(n3179) );
  XOR2X1 U1950 ( .A(n3146), .B(n5057), .Y(n2668) );
  OAI21X1 U1951 ( .A(n4939), .B(n4782), .C(n4176), .Y(n3146) );
  AOI21X1 U1952 ( .A(n4997), .B(n84), .C(n1772), .Y(n3180) );
  XOR2X1 U1955 ( .A(n3147), .B(n5057), .Y(n2669) );
  OAI21X1 U1956 ( .A(n4939), .B(n3916), .C(n4175), .Y(n3147) );
  AOI21X1 U1957 ( .A(n4995), .B(n84), .C(n1774), .Y(n3181) );
  XOR2X1 U1960 ( .A(n3148), .B(n5057), .Y(n2670) );
  OAI21X1 U1961 ( .A(n82), .B(n3921), .C(n4174), .Y(n3148) );
  AOI21X1 U1962 ( .A(n4993), .B(n84), .C(n1776), .Y(n3182) );
  XOR2X1 U1965 ( .A(n3149), .B(n5058), .Y(n2671) );
  OAI21X1 U1966 ( .A(n82), .B(n4784), .C(n4173), .Y(n3149) );
  AOI21X1 U1967 ( .A(n4991), .B(n84), .C(n1778), .Y(n3183) );
  XOR2X1 U1970 ( .A(n3150), .B(n5058), .Y(n2672) );
  OAI21X1 U1971 ( .A(n82), .B(n3920), .C(n4172), .Y(n3150) );
  AOI21X1 U1972 ( .A(n4989), .B(n84), .C(n1780), .Y(n3184) );
  XOR2X1 U1975 ( .A(n3151), .B(n5058), .Y(n2673) );
  OAI21X1 U1976 ( .A(n82), .B(n4802), .C(n4171), .Y(n3151) );
  AOI21X1 U1977 ( .A(n4987), .B(n84), .C(n1782), .Y(n3185) );
  XOR2X1 U1980 ( .A(n3152), .B(n5058), .Y(n2674) );
  OAI21X1 U1981 ( .A(n82), .B(n4801), .C(n4170), .Y(n3152) );
  AOI21X1 U1982 ( .A(b[3]), .B(n84), .C(n1784), .Y(n3186) );
  XOR2X1 U1985 ( .A(n3153), .B(n5058), .Y(n2675) );
  OAI21X1 U1986 ( .A(n82), .B(n3922), .C(n4169), .Y(n3153) );
  AOI21X1 U1987 ( .A(n4983), .B(n84), .C(n1786), .Y(n3187) );
  XOR2X1 U1990 ( .A(n3154), .B(n5058), .Y(n2676) );
  OAI21X1 U1991 ( .A(n82), .B(n3919), .C(n4168), .Y(n3154) );
  AOI21X1 U1992 ( .A(b[1]), .B(n84), .C(n1788), .Y(n3188) );
  XOR2X1 U1995 ( .A(n3155), .B(n5058), .Y(n2677) );
  OAI21X1 U1996 ( .A(n82), .B(n4765), .C(n4167), .Y(n3155) );
  AOI21X1 U1997 ( .A(b[0]), .B(n84), .C(n1790), .Y(n3189) );
  XOR2X1 U2000 ( .A(n3156), .B(n5058), .Y(n2678) );
  OAI21X1 U2001 ( .A(n82), .B(n4359), .C(n3973), .Y(n3156) );
  XOR2X1 U2003 ( .A(n3157), .B(n5058), .Y(n2679) );
  OAI21X1 U2004 ( .A(n82), .B(n4982), .C(n3190), .Y(n3157) );
  AND2X1 U2006 ( .A(n4941), .B(n4981), .Y(n1792) );
  XOR2X1 U2008 ( .A(n3191), .B(n5054), .Y(n2681) );
  OAI21X1 U2009 ( .A(n4942), .B(n3593), .C(n4487), .Y(n3191) );
  XOR2X1 U2011 ( .A(n3192), .B(n5054), .Y(n2682) );
  OAI21X1 U2012 ( .A(n4942), .B(n4809), .C(n4706), .Y(n3192) );
  AOI21X1 U2013 ( .A(n5033), .B(n72), .C(n1793), .Y(n3226) );
  AND2X1 U2014 ( .A(n64), .B(n5035), .Y(n1793) );
  XOR2X1 U2015 ( .A(n3193), .B(n5054), .Y(n2683) );
  OAI21X1 U2016 ( .A(n4942), .B(n4779), .C(n4166), .Y(n3193) );
  AOI21X1 U2017 ( .A(n5031), .B(n72), .C(n1795), .Y(n3227) );
  XOR2X1 U2020 ( .A(n3194), .B(n5054), .Y(n2684) );
  OAI21X1 U2021 ( .A(n4942), .B(n4780), .C(n4165), .Y(n3194) );
  AOI21X1 U2022 ( .A(n5029), .B(n72), .C(n1797), .Y(n3228) );
  XOR2X1 U2025 ( .A(n3195), .B(n5054), .Y(n2685) );
  OAI21X1 U2026 ( .A(n4942), .B(n4776), .C(n4164), .Y(n3195) );
  AOI21X1 U2027 ( .A(n5027), .B(n72), .C(n1799), .Y(n3229) );
  XOR2X1 U2030 ( .A(n3196), .B(n5054), .Y(n2686) );
  OAI21X1 U2031 ( .A(n4942), .B(n4769), .C(n4163), .Y(n3196) );
  AOI21X1 U2032 ( .A(n5025), .B(n72), .C(n1801), .Y(n3230) );
  XOR2X1 U2035 ( .A(n3197), .B(n5054), .Y(n2687) );
  OAI21X1 U2036 ( .A(n4942), .B(n4778), .C(n4162), .Y(n3197) );
  AOI21X1 U2037 ( .A(n5023), .B(n72), .C(n1803), .Y(n3231) );
  XOR2X1 U2040 ( .A(n3198), .B(n5055), .Y(n2688) );
  OAI21X1 U2041 ( .A(n4942), .B(n3914), .C(n4161), .Y(n3198) );
  AOI21X1 U2042 ( .A(n5021), .B(n72), .C(n1805), .Y(n3232) );
  XOR2X1 U2045 ( .A(n3199), .B(n5054), .Y(n2689) );
  OAI21X1 U2046 ( .A(n4942), .B(n4767), .C(n4160), .Y(n3199) );
  AOI21X1 U2047 ( .A(n5019), .B(n72), .C(n1807), .Y(n3233) );
  XOR2X1 U2050 ( .A(n3200), .B(n5054), .Y(n2690) );
  OAI21X1 U2051 ( .A(n4942), .B(n4775), .C(n4159), .Y(n3200) );
  AOI21X1 U2052 ( .A(b[22]), .B(n72), .C(n1809), .Y(n3234) );
  XOR2X1 U2055 ( .A(n3201), .B(n5054), .Y(n2691) );
  OAI21X1 U2056 ( .A(n70), .B(n4774), .C(n4158), .Y(n3201) );
  AOI21X1 U2057 ( .A(n5017), .B(n72), .C(n1811), .Y(n3235) );
  XOR2X1 U2060 ( .A(n3202), .B(n5054), .Y(n2692) );
  OAI21X1 U2061 ( .A(n70), .B(n4772), .C(n4157), .Y(n3202) );
  AOI21X1 U2062 ( .A(b[20]), .B(n72), .C(n1813), .Y(n3236) );
  XOR2X1 U2065 ( .A(n3203), .B(n5055), .Y(n2693) );
  OAI21X1 U2066 ( .A(n4942), .B(n4804), .C(n4156), .Y(n3203) );
  AOI21X1 U2067 ( .A(n5015), .B(n72), .C(n1815), .Y(n3237) );
  XOR2X1 U2070 ( .A(n3204), .B(n5055), .Y(n2694) );
  OAI21X1 U2071 ( .A(n4942), .B(n4803), .C(n4155), .Y(n3204) );
  AOI21X1 U2072 ( .A(n5013), .B(n72), .C(n1817), .Y(n3238) );
  XOR2X1 U2075 ( .A(n3205), .B(n5055), .Y(n2695) );
  OAI21X1 U2076 ( .A(n4942), .B(n4766), .C(n4154), .Y(n3205) );
  AOI21X1 U2077 ( .A(b[17]), .B(n72), .C(n1819), .Y(n3239) );
  XOR2X1 U2080 ( .A(n3206), .B(n5054), .Y(n2696) );
  OAI21X1 U2081 ( .A(n4942), .B(n4773), .C(n4153), .Y(n3206) );
  AOI21X1 U2082 ( .A(n5011), .B(n72), .C(n1821), .Y(n3240) );
  XOR2X1 U2085 ( .A(n3207), .B(n5054), .Y(n2697) );
  OAI21X1 U2086 ( .A(n4942), .B(n4768), .C(n4152), .Y(n3207) );
  AOI21X1 U2087 ( .A(n5009), .B(n72), .C(n1823), .Y(n3241) );
  XOR2X1 U2090 ( .A(n3208), .B(n5054), .Y(n2698) );
  OAI21X1 U2091 ( .A(n4942), .B(n3923), .C(n4151), .Y(n3208) );
  AOI21X1 U2092 ( .A(n5007), .B(n72), .C(n1825), .Y(n3242) );
  XOR2X1 U2095 ( .A(n3209), .B(n5054), .Y(n2699) );
  OAI21X1 U2096 ( .A(n4942), .B(n4783), .C(n4150), .Y(n3209) );
  AOI21X1 U2097 ( .A(n5005), .B(n72), .C(n1827), .Y(n3243) );
  XOR2X1 U2100 ( .A(n3210), .B(n5055), .Y(n2700) );
  OAI21X1 U2101 ( .A(n4942), .B(n3917), .C(n4149), .Y(n3210) );
  AOI21X1 U2102 ( .A(n5003), .B(n72), .C(n1829), .Y(n3244) );
  XOR2X1 U2105 ( .A(n3211), .B(n5055), .Y(n2701) );
  OAI21X1 U2106 ( .A(n4942), .B(n3913), .C(n4148), .Y(n3211) );
  AOI21X1 U2107 ( .A(n5001), .B(n72), .C(n1831), .Y(n3245) );
  XOR2X1 U2110 ( .A(n3212), .B(n5055), .Y(n2702) );
  OAI21X1 U2111 ( .A(n4942), .B(n3918), .C(n4147), .Y(n3212) );
  AOI21X1 U2112 ( .A(n4999), .B(n72), .C(n1833), .Y(n3246) );
  XOR2X1 U2115 ( .A(n3213), .B(n5054), .Y(n2703) );
  OAI21X1 U2116 ( .A(n4942), .B(n4782), .C(n4146), .Y(n3213) );
  AOI21X1 U2117 ( .A(n4997), .B(n72), .C(n1835), .Y(n3247) );
  XOR2X1 U2120 ( .A(n3214), .B(n5054), .Y(n2704) );
  OAI21X1 U2121 ( .A(n4942), .B(n3916), .C(n4145), .Y(n3214) );
  AOI21X1 U2122 ( .A(n4995), .B(n72), .C(n1837), .Y(n3248) );
  XOR2X1 U2125 ( .A(n3215), .B(n5054), .Y(n2705) );
  OAI21X1 U2126 ( .A(n70), .B(n3921), .C(n4144), .Y(n3215) );
  AOI21X1 U2127 ( .A(n4993), .B(n72), .C(n1839), .Y(n3249) );
  XOR2X1 U2130 ( .A(n3216), .B(n5055), .Y(n2706) );
  OAI21X1 U2131 ( .A(n70), .B(n4784), .C(n4143), .Y(n3216) );
  AOI21X1 U2132 ( .A(n4991), .B(n72), .C(n1841), .Y(n3250) );
  XOR2X1 U2135 ( .A(n3217), .B(n5055), .Y(n2707) );
  OAI21X1 U2136 ( .A(n70), .B(n3920), .C(n4142), .Y(n3217) );
  AOI21X1 U2137 ( .A(n4989), .B(n72), .C(n1843), .Y(n3251) );
  XOR2X1 U2140 ( .A(n3218), .B(n5055), .Y(n2708) );
  OAI21X1 U2141 ( .A(n70), .B(n4802), .C(n4141), .Y(n3218) );
  AOI21X1 U2142 ( .A(n4987), .B(n72), .C(n1845), .Y(n3252) );
  XOR2X1 U2145 ( .A(n3219), .B(n5055), .Y(n2709) );
  OAI21X1 U2146 ( .A(n70), .B(n4801), .C(n4140), .Y(n3219) );
  AOI21X1 U2147 ( .A(n4985), .B(n72), .C(n1847), .Y(n3253) );
  XOR2X1 U2150 ( .A(n3220), .B(n5055), .Y(n2710) );
  OAI21X1 U2151 ( .A(n70), .B(n3922), .C(n4139), .Y(n3220) );
  AOI21X1 U2152 ( .A(b[2]), .B(n72), .C(n1849), .Y(n3254) );
  XOR2X1 U2155 ( .A(n3221), .B(n5055), .Y(n2711) );
  OAI21X1 U2156 ( .A(n70), .B(n3919), .C(n4138), .Y(n3221) );
  AOI21X1 U2157 ( .A(b[1]), .B(n72), .C(n1851), .Y(n3255) );
  XOR2X1 U2160 ( .A(n3222), .B(n5055), .Y(n2712) );
  OAI21X1 U2161 ( .A(n70), .B(n4765), .C(n4137), .Y(n3222) );
  AOI21X1 U2162 ( .A(b[0]), .B(n72), .C(n1853), .Y(n3256) );
  XOR2X1 U2165 ( .A(n3223), .B(n5055), .Y(n2713) );
  OAI21X1 U2166 ( .A(n70), .B(n4359), .C(n3972), .Y(n3223) );
  XOR2X1 U2168 ( .A(n3224), .B(n5055), .Y(n2714) );
  OAI21X1 U2169 ( .A(n70), .B(n4982), .C(n3257), .Y(n3224) );
  AND2X1 U2171 ( .A(n4944), .B(n4981), .Y(n1855) );
  XOR2X1 U2173 ( .A(n3258), .B(n5051), .Y(n2716) );
  OAI21X1 U2174 ( .A(n4945), .B(n3593), .C(n4466), .Y(n3258) );
  XOR2X1 U2176 ( .A(n3259), .B(n5051), .Y(n2717) );
  OAI21X1 U2177 ( .A(n4945), .B(n4809), .C(n4578), .Y(n3259) );
  AOI21X1 U2178 ( .A(n5033), .B(n60), .C(n1856), .Y(n3293) );
  AND2X1 U2179 ( .A(n52), .B(n5035), .Y(n1856) );
  XOR2X1 U2180 ( .A(n3260), .B(n5051), .Y(n2718) );
  OAI21X1 U2181 ( .A(n4945), .B(n4779), .C(n4136), .Y(n3260) );
  AOI21X1 U2182 ( .A(n5031), .B(n60), .C(n1858), .Y(n3294) );
  XOR2X1 U2185 ( .A(n3261), .B(n5051), .Y(n2719) );
  OAI21X1 U2186 ( .A(n4945), .B(n4780), .C(n4135), .Y(n3261) );
  AOI21X1 U2187 ( .A(n5029), .B(n60), .C(n1860), .Y(n3295) );
  XOR2X1 U2190 ( .A(n3262), .B(n5051), .Y(n2720) );
  OAI21X1 U2191 ( .A(n4945), .B(n4776), .C(n4134), .Y(n3262) );
  AOI21X1 U2192 ( .A(n5027), .B(n60), .C(n1862), .Y(n3296) );
  XOR2X1 U2195 ( .A(n3263), .B(n5051), .Y(n2721) );
  OAI21X1 U2196 ( .A(n4945), .B(n4769), .C(n4133), .Y(n3263) );
  AOI21X1 U2197 ( .A(n5025), .B(n60), .C(n1864), .Y(n3297) );
  XOR2X1 U2200 ( .A(n3264), .B(n5051), .Y(n2722) );
  OAI21X1 U2201 ( .A(n4945), .B(n4778), .C(n4132), .Y(n3264) );
  AOI21X1 U2202 ( .A(n5023), .B(n60), .C(n1866), .Y(n3298) );
  XOR2X1 U2205 ( .A(n3265), .B(n5052), .Y(n2723) );
  OAI21X1 U2206 ( .A(n4945), .B(n3914), .C(n4131), .Y(n3265) );
  AOI21X1 U2207 ( .A(n5021), .B(n60), .C(n1868), .Y(n3299) );
  XOR2X1 U2210 ( .A(n3266), .B(n5051), .Y(n2724) );
  OAI21X1 U2211 ( .A(n4945), .B(n4767), .C(n4130), .Y(n3266) );
  AOI21X1 U2212 ( .A(n5019), .B(n60), .C(n1870), .Y(n3300) );
  XOR2X1 U2215 ( .A(n3267), .B(n5051), .Y(n2725) );
  OAI21X1 U2216 ( .A(n4945), .B(n4775), .C(n4129), .Y(n3267) );
  AOI21X1 U2217 ( .A(b[22]), .B(n60), .C(n1872), .Y(n3301) );
  XOR2X1 U2220 ( .A(n3268), .B(n5051), .Y(n2726) );
  OAI21X1 U2221 ( .A(n58), .B(n4774), .C(n4128), .Y(n3268) );
  AOI21X1 U2222 ( .A(n5017), .B(n60), .C(n1874), .Y(n3302) );
  XOR2X1 U2225 ( .A(n3269), .B(n5052), .Y(n2727) );
  OAI21X1 U2226 ( .A(n58), .B(n4772), .C(n4127), .Y(n3269) );
  AOI21X1 U2227 ( .A(b[20]), .B(n60), .C(n1876), .Y(n3303) );
  XOR2X1 U2230 ( .A(n3270), .B(n5051), .Y(n2728) );
  OAI21X1 U2231 ( .A(n4945), .B(n4804), .C(n4126), .Y(n3270) );
  AOI21X1 U2232 ( .A(n5015), .B(n60), .C(n1878), .Y(n3304) );
  XOR2X1 U2235 ( .A(n3271), .B(n5051), .Y(n2729) );
  OAI21X1 U2236 ( .A(n4945), .B(n4803), .C(n4125), .Y(n3271) );
  AOI21X1 U2237 ( .A(n5013), .B(n60), .C(n1880), .Y(n3305) );
  XOR2X1 U2240 ( .A(n3272), .B(n5051), .Y(n2730) );
  OAI21X1 U2241 ( .A(n4945), .B(n4766), .C(n4124), .Y(n3272) );
  AOI21X1 U2242 ( .A(b[17]), .B(n60), .C(n1882), .Y(n3306) );
  XOR2X1 U2245 ( .A(n3273), .B(a[14]), .Y(n2731) );
  OAI21X1 U2246 ( .A(n4945), .B(n4773), .C(n4123), .Y(n3273) );
  AOI21X1 U2247 ( .A(n5011), .B(n60), .C(n1884), .Y(n3307) );
  XOR2X1 U2250 ( .A(n3274), .B(a[14]), .Y(n2732) );
  OAI21X1 U2251 ( .A(n4945), .B(n4768), .C(n4122), .Y(n3274) );
  AOI21X1 U2252 ( .A(n5009), .B(n60), .C(n1886), .Y(n3308) );
  XOR2X1 U2255 ( .A(n3275), .B(n5051), .Y(n2733) );
  OAI21X1 U2256 ( .A(n4945), .B(n3923), .C(n4121), .Y(n3275) );
  AOI21X1 U2257 ( .A(n5007), .B(n60), .C(n1888), .Y(n3309) );
  XOR2X1 U2260 ( .A(n3276), .B(a[14]), .Y(n2734) );
  OAI21X1 U2261 ( .A(n4945), .B(n4783), .C(n4120), .Y(n3276) );
  AOI21X1 U2262 ( .A(n5005), .B(n60), .C(n1890), .Y(n3310) );
  XOR2X1 U2265 ( .A(n3277), .B(n5052), .Y(n2735) );
  OAI21X1 U2266 ( .A(n4945), .B(n3917), .C(n4119), .Y(n3277) );
  AOI21X1 U2267 ( .A(n5003), .B(n60), .C(n1892), .Y(n3311) );
  XOR2X1 U2270 ( .A(n3278), .B(n5052), .Y(n2736) );
  OAI21X1 U2271 ( .A(n4945), .B(n3913), .C(n4118), .Y(n3278) );
  AOI21X1 U2272 ( .A(n5001), .B(n60), .C(n1894), .Y(n3312) );
  XOR2X1 U2275 ( .A(n3279), .B(n5052), .Y(n2737) );
  OAI21X1 U2276 ( .A(n4945), .B(n3918), .C(n4117), .Y(n3279) );
  AOI21X1 U2277 ( .A(n4999), .B(n60), .C(n1896), .Y(n3313) );
  XOR2X1 U2280 ( .A(n3280), .B(n5051), .Y(n2738) );
  OAI21X1 U2281 ( .A(n4945), .B(n4782), .C(n4116), .Y(n3280) );
  AOI21X1 U2282 ( .A(n4997), .B(n60), .C(n1898), .Y(n3314) );
  XOR2X1 U2285 ( .A(n3281), .B(n5051), .Y(n2739) );
  OAI21X1 U2286 ( .A(n4945), .B(n3916), .C(n4115), .Y(n3281) );
  AOI21X1 U2287 ( .A(n4995), .B(n60), .C(n1900), .Y(n3315) );
  XOR2X1 U2290 ( .A(n3282), .B(n5051), .Y(n2740) );
  OAI21X1 U2291 ( .A(n58), .B(n3921), .C(n4114), .Y(n3282) );
  AOI21X1 U2292 ( .A(n4993), .B(n60), .C(n1902), .Y(n3316) );
  XOR2X1 U2295 ( .A(n3283), .B(n5052), .Y(n2741) );
  OAI21X1 U2296 ( .A(n58), .B(n4784), .C(n4113), .Y(n3283) );
  AOI21X1 U2297 ( .A(n4991), .B(n60), .C(n1904), .Y(n3317) );
  XOR2X1 U2300 ( .A(n3284), .B(n5052), .Y(n2742) );
  OAI21X1 U2301 ( .A(n58), .B(n3920), .C(n4112), .Y(n3284) );
  AOI21X1 U2302 ( .A(n4989), .B(n60), .C(n1906), .Y(n3318) );
  XOR2X1 U2305 ( .A(n3285), .B(n5052), .Y(n2743) );
  OAI21X1 U2306 ( .A(n4945), .B(n4802), .C(n4111), .Y(n3285) );
  AOI21X1 U2307 ( .A(n4987), .B(n60), .C(n1908), .Y(n3319) );
  XOR2X1 U2310 ( .A(n3286), .B(n5052), .Y(n2744) );
  OAI21X1 U2311 ( .A(n4945), .B(n4801), .C(n4110), .Y(n3286) );
  AOI21X1 U2312 ( .A(n4985), .B(n60), .C(n1910), .Y(n3320) );
  XOR2X1 U2315 ( .A(n3287), .B(n5052), .Y(n2745) );
  OAI21X1 U2316 ( .A(n4945), .B(n3922), .C(n4109), .Y(n3287) );
  AOI21X1 U2317 ( .A(n4983), .B(n60), .C(n1912), .Y(n3321) );
  XOR2X1 U2320 ( .A(n3288), .B(n5052), .Y(n2746) );
  OAI21X1 U2321 ( .A(n58), .B(n3919), .C(n4108), .Y(n3288) );
  AOI21X1 U2322 ( .A(b[1]), .B(n60), .C(n1914), .Y(n3322) );
  XOR2X1 U2325 ( .A(n3289), .B(n5052), .Y(n2747) );
  OAI21X1 U2326 ( .A(n58), .B(n4765), .C(n4107), .Y(n3289) );
  AOI21X1 U2327 ( .A(b[0]), .B(n60), .C(n1916), .Y(n3323) );
  XOR2X1 U2330 ( .A(n3290), .B(n5052), .Y(n2748) );
  OAI21X1 U2331 ( .A(n58), .B(n4359), .C(n3971), .Y(n3290) );
  XOR2X1 U2333 ( .A(n3291), .B(n5052), .Y(n2749) );
  OAI21X1 U2334 ( .A(n58), .B(n4982), .C(n3324), .Y(n3291) );
  AND2X1 U2336 ( .A(n4948), .B(b[0]), .Y(n1918) );
  XOR2X1 U2338 ( .A(n3325), .B(n5048), .Y(n2751) );
  OAI21X1 U2339 ( .A(n4951), .B(n3593), .C(n4577), .Y(n3325) );
  XOR2X1 U2341 ( .A(n3326), .B(n5048), .Y(n2752) );
  OAI21X1 U2342 ( .A(n4951), .B(n4809), .C(n4640), .Y(n3326) );
  AOI21X1 U2343 ( .A(n5033), .B(n48), .C(n1919), .Y(n3360) );
  AND2X1 U2344 ( .A(n40), .B(n5036), .Y(n1919) );
  XOR2X1 U2345 ( .A(n3327), .B(n5048), .Y(n2753) );
  OAI21X1 U2346 ( .A(n4951), .B(n4779), .C(n4106), .Y(n3327) );
  AOI21X1 U2347 ( .A(n5031), .B(n48), .C(n1921), .Y(n3361) );
  XOR2X1 U2350 ( .A(n3328), .B(n5048), .Y(n2754) );
  OAI21X1 U2351 ( .A(n4951), .B(n4780), .C(n4105), .Y(n3328) );
  AOI21X1 U2352 ( .A(n5029), .B(n48), .C(n1923), .Y(n3362) );
  XOR2X1 U2355 ( .A(n3329), .B(n5048), .Y(n2755) );
  OAI21X1 U2356 ( .A(n4951), .B(n4776), .C(n4104), .Y(n3329) );
  AOI21X1 U2357 ( .A(n5027), .B(n48), .C(n1925), .Y(n3363) );
  XOR2X1 U2360 ( .A(n3330), .B(n5048), .Y(n2756) );
  OAI21X1 U2361 ( .A(n4951), .B(n4769), .C(n4103), .Y(n3330) );
  AOI21X1 U2362 ( .A(n5025), .B(n48), .C(n1927), .Y(n3364) );
  XOR2X1 U2365 ( .A(n3331), .B(n5048), .Y(n2757) );
  OAI21X1 U2366 ( .A(n4951), .B(n4778), .C(n4102), .Y(n3331) );
  AOI21X1 U2367 ( .A(n5023), .B(n4949), .C(n1929), .Y(n3365) );
  XOR2X1 U2370 ( .A(n3332), .B(n5049), .Y(n2758) );
  OAI21X1 U2371 ( .A(n4951), .B(n3914), .C(n4101), .Y(n3332) );
  AOI21X1 U2372 ( .A(n5021), .B(n4949), .C(n1931), .Y(n3366) );
  XOR2X1 U2375 ( .A(n3333), .B(n5048), .Y(n2759) );
  OAI21X1 U2376 ( .A(n4951), .B(n4767), .C(n4100), .Y(n3333) );
  AOI21X1 U2377 ( .A(n5019), .B(n4949), .C(n1933), .Y(n3367) );
  XOR2X1 U2380 ( .A(n3334), .B(n5048), .Y(n2760) );
  OAI21X1 U2381 ( .A(n4951), .B(n4775), .C(n4099), .Y(n3334) );
  AOI21X1 U2382 ( .A(b[22]), .B(n4949), .C(n1935), .Y(n3368) );
  XOR2X1 U2385 ( .A(n3335), .B(n5048), .Y(n2761) );
  OAI21X1 U2386 ( .A(n46), .B(n4774), .C(n4098), .Y(n3335) );
  AOI21X1 U2387 ( .A(n5017), .B(n4949), .C(n1937), .Y(n3369) );
  XOR2X1 U2390 ( .A(n3336), .B(n5048), .Y(n2762) );
  OAI21X1 U2391 ( .A(n4951), .B(n4772), .C(n4097), .Y(n3336) );
  AOI21X1 U2392 ( .A(b[20]), .B(n4949), .C(n1939), .Y(n3370) );
  XOR2X1 U2395 ( .A(n3337), .B(n5048), .Y(n2763) );
  OAI21X1 U2396 ( .A(n4951), .B(n4804), .C(n4096), .Y(n3337) );
  AOI21X1 U2397 ( .A(n5015), .B(n4949), .C(n1941), .Y(n3371) );
  XOR2X1 U2400 ( .A(n3338), .B(n5048), .Y(n2764) );
  OAI21X1 U2401 ( .A(n4951), .B(n4803), .C(n4095), .Y(n3338) );
  AOI21X1 U2402 ( .A(n5013), .B(n4949), .C(n1943), .Y(n3372) );
  XOR2X1 U2405 ( .A(n3339), .B(n5048), .Y(n2765) );
  OAI21X1 U2406 ( .A(n4951), .B(n4766), .C(n4094), .Y(n3339) );
  AOI21X1 U2407 ( .A(b[17]), .B(n4949), .C(n1945), .Y(n3373) );
  XOR2X1 U2410 ( .A(n3340), .B(n5049), .Y(n2766) );
  OAI21X1 U2411 ( .A(n4951), .B(n4773), .C(n4093), .Y(n3340) );
  AOI21X1 U2412 ( .A(n5011), .B(n4949), .C(n1947), .Y(n3374) );
  XOR2X1 U2415 ( .A(n3341), .B(n5049), .Y(n2767) );
  OAI21X1 U2416 ( .A(n4951), .B(n4768), .C(n4092), .Y(n3341) );
  AOI21X1 U2417 ( .A(n5009), .B(n48), .C(n1949), .Y(n3375) );
  XOR2X1 U2420 ( .A(n3342), .B(n5048), .Y(n2768) );
  OAI21X1 U2421 ( .A(n4951), .B(n3923), .C(n4091), .Y(n3342) );
  AOI21X1 U2422 ( .A(n5007), .B(n48), .C(n1951), .Y(n3376) );
  XOR2X1 U2425 ( .A(n3343), .B(n5048), .Y(n2769) );
  OAI21X1 U2426 ( .A(n4951), .B(n4783), .C(n4090), .Y(n3343) );
  AOI21X1 U2427 ( .A(n5005), .B(n48), .C(n1953), .Y(n3377) );
  XOR2X1 U2430 ( .A(n3344), .B(n5049), .Y(n2770) );
  OAI21X1 U2431 ( .A(n4951), .B(n3917), .C(n4089), .Y(n3344) );
  AOI21X1 U2432 ( .A(n5003), .B(n48), .C(n1955), .Y(n3378) );
  XOR2X1 U2435 ( .A(n3345), .B(n5049), .Y(n2771) );
  OAI21X1 U2436 ( .A(n4951), .B(n3913), .C(n4088), .Y(n3345) );
  AOI21X1 U2437 ( .A(n5001), .B(n48), .C(n1957), .Y(n3379) );
  XOR2X1 U2440 ( .A(n3346), .B(n5049), .Y(n2772) );
  OAI21X1 U2441 ( .A(n4951), .B(n3918), .C(n4087), .Y(n3346) );
  AOI21X1 U2442 ( .A(n4999), .B(n48), .C(n1959), .Y(n3380) );
  XOR2X1 U2445 ( .A(n3347), .B(n5048), .Y(n2773) );
  OAI21X1 U2446 ( .A(n4951), .B(n4782), .C(n4086), .Y(n3347) );
  AOI21X1 U2447 ( .A(n4997), .B(n48), .C(n1961), .Y(n3381) );
  XOR2X1 U2450 ( .A(n3348), .B(n5048), .Y(n2774) );
  OAI21X1 U2451 ( .A(n4951), .B(n3916), .C(n4085), .Y(n3348) );
  AOI21X1 U2452 ( .A(n4995), .B(n48), .C(n1963), .Y(n3382) );
  XOR2X1 U2455 ( .A(n3349), .B(n5048), .Y(n2775) );
  OAI21X1 U2456 ( .A(n4951), .B(n3921), .C(n4084), .Y(n3349) );
  AOI21X1 U2457 ( .A(n4993), .B(n48), .C(n1965), .Y(n3383) );
  XOR2X1 U2460 ( .A(n3350), .B(n5049), .Y(n2776) );
  OAI21X1 U2461 ( .A(n4951), .B(n4784), .C(n4083), .Y(n3350) );
  AOI21X1 U2462 ( .A(n4991), .B(n48), .C(n1967), .Y(n3384) );
  XOR2X1 U2465 ( .A(n3351), .B(n5049), .Y(n2777) );
  OAI21X1 U2466 ( .A(n4951), .B(n3920), .C(n4082), .Y(n3351) );
  AOI21X1 U2467 ( .A(n4989), .B(n48), .C(n1969), .Y(n3385) );
  XOR2X1 U2470 ( .A(n3352), .B(n5049), .Y(n2778) );
  OAI21X1 U2471 ( .A(n46), .B(n4802), .C(n4081), .Y(n3352) );
  AOI21X1 U2472 ( .A(n4987), .B(n48), .C(n1971), .Y(n3386) );
  XOR2X1 U2475 ( .A(n3353), .B(n5049), .Y(n2779) );
  OAI21X1 U2476 ( .A(n46), .B(n4801), .C(n4080), .Y(n3353) );
  AOI21X1 U2477 ( .A(n4985), .B(n48), .C(n1973), .Y(n3387) );
  XOR2X1 U2480 ( .A(n3354), .B(n5049), .Y(n2780) );
  OAI21X1 U2481 ( .A(n46), .B(n3922), .C(n4079), .Y(n3354) );
  AOI21X1 U2482 ( .A(b[2]), .B(n4949), .C(n1975), .Y(n3388) );
  XOR2X1 U2485 ( .A(n3355), .B(n5049), .Y(n2781) );
  OAI21X1 U2486 ( .A(n46), .B(n3919), .C(n4078), .Y(n3355) );
  AOI21X1 U2487 ( .A(b[1]), .B(n4949), .C(n1977), .Y(n3389) );
  XOR2X1 U2490 ( .A(n3356), .B(n5049), .Y(n2782) );
  OAI21X1 U2491 ( .A(n46), .B(n4765), .C(n4077), .Y(n3356) );
  AOI21X1 U2492 ( .A(b[0]), .B(n4949), .C(n1979), .Y(n3390) );
  XOR2X1 U2495 ( .A(n3357), .B(n5049), .Y(n2783) );
  OAI21X1 U2496 ( .A(n46), .B(n4359), .C(n3970), .Y(n3357) );
  XOR2X1 U2498 ( .A(n3358), .B(n5049), .Y(n2784) );
  OAI21X1 U2499 ( .A(n46), .B(n4982), .C(n3391), .Y(n3358) );
  AND2X1 U2501 ( .A(n4955), .B(n4981), .Y(n1981) );
  XOR2X1 U2503 ( .A(n3392), .B(n5045), .Y(n2786) );
  OAI21X1 U2504 ( .A(n4959), .B(n3593), .C(n4448), .Y(n3392) );
  XOR2X1 U2506 ( .A(n3393), .B(n5045), .Y(n2787) );
  OAI21X1 U2507 ( .A(n4959), .B(n4809), .C(n4454), .Y(n3393) );
  AOI21X1 U2508 ( .A(n5033), .B(n4956), .C(n1982), .Y(n3427) );
  AND2X1 U2509 ( .A(n4961), .B(n5036), .Y(n1982) );
  XOR2X1 U2510 ( .A(n3394), .B(n5045), .Y(n2788) );
  OAI21X1 U2511 ( .A(n4959), .B(n4779), .C(n4076), .Y(n3394) );
  AOI21X1 U2512 ( .A(n5031), .B(n4956), .C(n1984), .Y(n3428) );
  XOR2X1 U2515 ( .A(n3395), .B(n5045), .Y(n2789) );
  OAI21X1 U2516 ( .A(n4959), .B(n4780), .C(n4075), .Y(n3395) );
  AOI21X1 U2517 ( .A(n5029), .B(n4956), .C(n1986), .Y(n3429) );
  XOR2X1 U2520 ( .A(n3396), .B(n5045), .Y(n2790) );
  OAI21X1 U2521 ( .A(n4959), .B(n4776), .C(n4074), .Y(n3396) );
  AOI21X1 U2522 ( .A(n5027), .B(n4956), .C(n1988), .Y(n3430) );
  XOR2X1 U2525 ( .A(n3397), .B(n5045), .Y(n2791) );
  OAI21X1 U2526 ( .A(n4959), .B(n4769), .C(n4073), .Y(n3397) );
  AOI21X1 U2527 ( .A(n5025), .B(n4956), .C(n1990), .Y(n3431) );
  XOR2X1 U2530 ( .A(n3398), .B(n5045), .Y(n2792) );
  OAI21X1 U2531 ( .A(n4959), .B(n4778), .C(n4072), .Y(n3398) );
  AOI21X1 U2532 ( .A(n5023), .B(n4957), .C(n1992), .Y(n3432) );
  XOR2X1 U2535 ( .A(n3399), .B(n5046), .Y(n2793) );
  OAI21X1 U2536 ( .A(n4959), .B(n3914), .C(n4071), .Y(n3399) );
  AOI21X1 U2537 ( .A(n5021), .B(n4957), .C(n1994), .Y(n3433) );
  XOR2X1 U2540 ( .A(n3400), .B(n5045), .Y(n2794) );
  OAI21X1 U2541 ( .A(n4959), .B(n4767), .C(n4070), .Y(n3400) );
  AOI21X1 U2542 ( .A(n5019), .B(n4957), .C(n1996), .Y(n3434) );
  XOR2X1 U2545 ( .A(n3401), .B(n5045), .Y(n2795) );
  OAI21X1 U2546 ( .A(n4959), .B(n4775), .C(n4069), .Y(n3401) );
  AOI21X1 U2547 ( .A(b[22]), .B(n4957), .C(n1998), .Y(n3435) );
  XOR2X1 U2550 ( .A(n3402), .B(n5045), .Y(n2796) );
  OAI21X1 U2551 ( .A(n34), .B(n4774), .C(n4068), .Y(n3402) );
  AOI21X1 U2552 ( .A(n5017), .B(n4957), .C(n2000), .Y(n3436) );
  XOR2X1 U2555 ( .A(n3403), .B(n5045), .Y(n2797) );
  OAI21X1 U2556 ( .A(n34), .B(n4772), .C(n4067), .Y(n3403) );
  AOI21X1 U2557 ( .A(b[20]), .B(n4957), .C(n2002), .Y(n3437) );
  XOR2X1 U2560 ( .A(n3404), .B(n5045), .Y(n2798) );
  OAI21X1 U2561 ( .A(n4959), .B(n4804), .C(n4066), .Y(n3404) );
  AOI21X1 U2562 ( .A(n5015), .B(n4957), .C(n2004), .Y(n3438) );
  XOR2X1 U2565 ( .A(n3405), .B(a[8]), .Y(n2799) );
  OAI21X1 U2566 ( .A(n4959), .B(n4803), .C(n4065), .Y(n3405) );
  AOI21X1 U2567 ( .A(n5013), .B(n4957), .C(n2006), .Y(n3439) );
  XOR2X1 U2570 ( .A(n3406), .B(n5045), .Y(n2800) );
  OAI21X1 U2571 ( .A(n4959), .B(n4766), .C(n4064), .Y(n3406) );
  AOI21X1 U2572 ( .A(b[17]), .B(n4957), .C(n2008), .Y(n3440) );
  XOR2X1 U2575 ( .A(n3407), .B(n5046), .Y(n2801) );
  OAI21X1 U2576 ( .A(n4959), .B(n4773), .C(n4063), .Y(n3407) );
  AOI21X1 U2577 ( .A(n5011), .B(n4957), .C(n2010), .Y(n3441) );
  XOR2X1 U2580 ( .A(n3408), .B(n5045), .Y(n2802) );
  OAI21X1 U2581 ( .A(n4959), .B(n4768), .C(n4062), .Y(n3408) );
  AOI21X1 U2582 ( .A(n5009), .B(n4956), .C(n2012), .Y(n3442) );
  XOR2X1 U2585 ( .A(n3409), .B(n5045), .Y(n2803) );
  OAI21X1 U2586 ( .A(n4959), .B(n3923), .C(n4061), .Y(n3409) );
  AOI21X1 U2587 ( .A(n5007), .B(n4956), .C(n2014), .Y(n3443) );
  XOR2X1 U2590 ( .A(n3410), .B(a[8]), .Y(n2804) );
  OAI21X1 U2591 ( .A(n4959), .B(n4783), .C(n4060), .Y(n3410) );
  AOI21X1 U2592 ( .A(n5005), .B(n4956), .C(n2016), .Y(n3444) );
  XOR2X1 U2595 ( .A(n3411), .B(n5046), .Y(n2805) );
  OAI21X1 U2596 ( .A(n4959), .B(n3917), .C(n4059), .Y(n3411) );
  AOI21X1 U2597 ( .A(n5003), .B(n4956), .C(n2018), .Y(n3445) );
  XOR2X1 U2600 ( .A(n3412), .B(n5046), .Y(n2806) );
  OAI21X1 U2601 ( .A(n4959), .B(n3913), .C(n4058), .Y(n3412) );
  AOI21X1 U2602 ( .A(n5001), .B(n4956), .C(n2020), .Y(n3446) );
  XOR2X1 U2605 ( .A(n3413), .B(n5046), .Y(n2807) );
  OAI21X1 U2606 ( .A(n4959), .B(n3918), .C(n4057), .Y(n3413) );
  AOI21X1 U2607 ( .A(n4999), .B(n4956), .C(n2022), .Y(n3447) );
  XOR2X1 U2610 ( .A(n3414), .B(n5045), .Y(n2808) );
  OAI21X1 U2611 ( .A(n4959), .B(n4782), .C(n4056), .Y(n3414) );
  AOI21X1 U2612 ( .A(n4997), .B(n4956), .C(n2024), .Y(n3448) );
  XOR2X1 U2615 ( .A(n3415), .B(n5045), .Y(n2809) );
  OAI21X1 U2616 ( .A(n4959), .B(n3916), .C(n4055), .Y(n3415) );
  AOI21X1 U2617 ( .A(n4995), .B(n4956), .C(n2026), .Y(n3449) );
  XOR2X1 U2620 ( .A(n3416), .B(n5045), .Y(n2810) );
  OAI21X1 U2621 ( .A(n34), .B(n3921), .C(n4054), .Y(n3416) );
  AOI21X1 U2622 ( .A(n4993), .B(n4956), .C(n2028), .Y(n3450) );
  XOR2X1 U2625 ( .A(n3417), .B(n5046), .Y(n2811) );
  OAI21X1 U2626 ( .A(n34), .B(n4784), .C(n4053), .Y(n3417) );
  AOI21X1 U2627 ( .A(n4991), .B(n4956), .C(n2030), .Y(n3451) );
  XOR2X1 U2630 ( .A(n3418), .B(n5046), .Y(n2812) );
  OAI21X1 U2631 ( .A(n4959), .B(n3920), .C(n4052), .Y(n3418) );
  AOI21X1 U2632 ( .A(n4989), .B(n4956), .C(n2032), .Y(n3452) );
  XOR2X1 U2635 ( .A(n3419), .B(n5046), .Y(n2813) );
  OAI21X1 U2636 ( .A(n4959), .B(n4802), .C(n4051), .Y(n3419) );
  AOI21X1 U2637 ( .A(n4987), .B(n4956), .C(n2034), .Y(n3453) );
  XOR2X1 U2640 ( .A(n3420), .B(n5046), .Y(n2814) );
  OAI21X1 U2641 ( .A(n34), .B(n4801), .C(n4050), .Y(n3420) );
  AOI21X1 U2642 ( .A(b[3]), .B(n4956), .C(n2036), .Y(n3454) );
  XOR2X1 U2645 ( .A(n3421), .B(n5046), .Y(n2815) );
  OAI21X1 U2646 ( .A(n34), .B(n3922), .C(n4049), .Y(n3421) );
  AOI21X1 U2647 ( .A(n4983), .B(n4957), .C(n2038), .Y(n3455) );
  XOR2X1 U2650 ( .A(n3422), .B(n5046), .Y(n2816) );
  OAI21X1 U2651 ( .A(n34), .B(n3919), .C(n4048), .Y(n3422) );
  AOI21X1 U2652 ( .A(b[1]), .B(n4957), .C(n2040), .Y(n3456) );
  XOR2X1 U2655 ( .A(n3423), .B(n5046), .Y(n2817) );
  OAI21X1 U2656 ( .A(n34), .B(n4765), .C(n4047), .Y(n3423) );
  AOI21X1 U2657 ( .A(n4981), .B(n4957), .C(n2042), .Y(n3457) );
  XOR2X1 U2660 ( .A(n3424), .B(n5046), .Y(n2818) );
  OAI21X1 U2661 ( .A(n34), .B(n4359), .C(n3968), .Y(n3424) );
  XOR2X1 U2663 ( .A(n3425), .B(n5046), .Y(n2819) );
  OAI21X1 U2664 ( .A(n34), .B(n4982), .C(n3458), .Y(n3425) );
  AND2X1 U2666 ( .A(n4963), .B(b[0]), .Y(n2044) );
  XOR2X1 U2668 ( .A(n3459), .B(n5042), .Y(n2821) );
  OAI21X1 U2669 ( .A(n4968), .B(n3593), .C(n4705), .Y(n3459) );
  XOR2X1 U2671 ( .A(n3460), .B(n5042), .Y(n2822) );
  OAI21X1 U2672 ( .A(n4968), .B(n4809), .C(n4467), .Y(n3460) );
  AOI21X1 U2673 ( .A(n5033), .B(n4965), .C(n2045), .Y(n3494) );
  AND2X1 U2674 ( .A(n4970), .B(n5036), .Y(n2045) );
  XOR2X1 U2675 ( .A(n3461), .B(n5042), .Y(n2823) );
  OAI21X1 U2676 ( .A(n4968), .B(n4779), .C(n4046), .Y(n3461) );
  AOI21X1 U2677 ( .A(n5031), .B(n4965), .C(n2047), .Y(n3495) );
  XOR2X1 U2680 ( .A(n3462), .B(n5042), .Y(n2824) );
  OAI21X1 U2681 ( .A(n4968), .B(n4780), .C(n4045), .Y(n3462) );
  AOI21X1 U2682 ( .A(n5029), .B(n4965), .C(n2049), .Y(n3496) );
  XOR2X1 U2685 ( .A(n3463), .B(n5042), .Y(n2825) );
  OAI21X1 U2686 ( .A(n4968), .B(n4776), .C(n4044), .Y(n3463) );
  AOI21X1 U2687 ( .A(n5027), .B(n4965), .C(n2051), .Y(n3497) );
  XOR2X1 U2690 ( .A(n3464), .B(n5042), .Y(n2826) );
  OAI21X1 U2691 ( .A(n4968), .B(n4769), .C(n4043), .Y(n3464) );
  AOI21X1 U2692 ( .A(n5025), .B(n4965), .C(n2053), .Y(n3498) );
  XOR2X1 U2695 ( .A(n3465), .B(n5042), .Y(n2827) );
  OAI21X1 U2696 ( .A(n4968), .B(n4778), .C(n4042), .Y(n3465) );
  AOI21X1 U2697 ( .A(n5023), .B(n4966), .C(n2055), .Y(n3499) );
  XOR2X1 U2700 ( .A(n3466), .B(n5043), .Y(n2828) );
  OAI21X1 U2701 ( .A(n4968), .B(n3914), .C(n4041), .Y(n3466) );
  AOI21X1 U2702 ( .A(n5021), .B(n4966), .C(n2057), .Y(n3500) );
  XOR2X1 U2705 ( .A(n3467), .B(n5042), .Y(n2829) );
  OAI21X1 U2706 ( .A(n4968), .B(n4767), .C(n4040), .Y(n3467) );
  AOI21X1 U2707 ( .A(n5019), .B(n4966), .C(n2059), .Y(n3501) );
  XOR2X1 U2710 ( .A(n3468), .B(n5042), .Y(n2830) );
  OAI21X1 U2711 ( .A(n4968), .B(n4775), .C(n4039), .Y(n3468) );
  AOI21X1 U2712 ( .A(b[22]), .B(n4966), .C(n2061), .Y(n3502) );
  XOR2X1 U2715 ( .A(n3469), .B(n5042), .Y(n2831) );
  OAI21X1 U2716 ( .A(n22), .B(n4774), .C(n4038), .Y(n3469) );
  AOI21X1 U2717 ( .A(n5017), .B(n4966), .C(n2063), .Y(n3503) );
  XOR2X1 U2720 ( .A(n3470), .B(a[5]), .Y(n2832) );
  OAI21X1 U2721 ( .A(n22), .B(n4772), .C(n4037), .Y(n3470) );
  AOI21X1 U2722 ( .A(b[20]), .B(n4966), .C(n2065), .Y(n3504) );
  XOR2X1 U2725 ( .A(n3471), .B(n5042), .Y(n2833) );
  OAI21X1 U2726 ( .A(n4968), .B(n4804), .C(n4036), .Y(n3471) );
  AOI21X1 U2727 ( .A(n5015), .B(n4966), .C(n2067), .Y(n3505) );
  XOR2X1 U2730 ( .A(n3472), .B(n5043), .Y(n2834) );
  OAI21X1 U2731 ( .A(n4968), .B(n4803), .C(n4035), .Y(n3472) );
  AOI21X1 U2732 ( .A(n5013), .B(n4966), .C(n2069), .Y(n3506) );
  XOR2X1 U2735 ( .A(n3473), .B(a[5]), .Y(n2835) );
  OAI21X1 U2736 ( .A(n4968), .B(n4766), .C(n4034), .Y(n3473) );
  AOI21X1 U2737 ( .A(b[17]), .B(n4966), .C(n2071), .Y(n3507) );
  XOR2X1 U2740 ( .A(n3474), .B(a[5]), .Y(n2836) );
  OAI21X1 U2741 ( .A(n4968), .B(n4773), .C(n4033), .Y(n3474) );
  AOI21X1 U2742 ( .A(n5011), .B(n4966), .C(n2073), .Y(n3508) );
  XOR2X1 U2745 ( .A(n3475), .B(n5042), .Y(n2837) );
  OAI21X1 U2746 ( .A(n4968), .B(n4768), .C(n4032), .Y(n3475) );
  AOI21X1 U2747 ( .A(n5009), .B(n4965), .C(n2075), .Y(n3509) );
  XOR2X1 U2750 ( .A(n3476), .B(n5042), .Y(n2838) );
  OAI21X1 U2751 ( .A(n4968), .B(n3923), .C(n4031), .Y(n3476) );
  AOI21X1 U2752 ( .A(n5007), .B(n4965), .C(n2077), .Y(n3510) );
  XOR2X1 U2755 ( .A(n3477), .B(n5043), .Y(n2839) );
  OAI21X1 U2756 ( .A(n4968), .B(n4783), .C(n4030), .Y(n3477) );
  AOI21X1 U2757 ( .A(n5005), .B(n4965), .C(n2079), .Y(n3511) );
  XOR2X1 U2760 ( .A(n3478), .B(n5043), .Y(n2840) );
  OAI21X1 U2761 ( .A(n4968), .B(n3917), .C(n4029), .Y(n3478) );
  AOI21X1 U2762 ( .A(n5003), .B(n4965), .C(n2081), .Y(n3512) );
  XOR2X1 U2765 ( .A(n3479), .B(n5043), .Y(n2841) );
  OAI21X1 U2766 ( .A(n4968), .B(n3913), .C(n4028), .Y(n3479) );
  AOI21X1 U2767 ( .A(n5001), .B(n4965), .C(n2083), .Y(n3513) );
  XOR2X1 U2770 ( .A(n3480), .B(n5043), .Y(n2842) );
  OAI21X1 U2771 ( .A(n4968), .B(n3918), .C(n4027), .Y(n3480) );
  AOI21X1 U2772 ( .A(n4999), .B(n4965), .C(n2085), .Y(n3514) );
  XOR2X1 U2775 ( .A(n3481), .B(n5042), .Y(n2843) );
  OAI21X1 U2776 ( .A(n4968), .B(n4782), .C(n4026), .Y(n3481) );
  AOI21X1 U2777 ( .A(n4997), .B(n4965), .C(n2087), .Y(n3515) );
  XOR2X1 U2780 ( .A(n3482), .B(n5042), .Y(n2844) );
  OAI21X1 U2781 ( .A(n4968), .B(n3916), .C(n4025), .Y(n3482) );
  AOI21X1 U2782 ( .A(n4995), .B(n4965), .C(n2089), .Y(n3516) );
  XOR2X1 U2785 ( .A(n3483), .B(n5042), .Y(n2845) );
  OAI21X1 U2786 ( .A(n22), .B(n3921), .C(n4024), .Y(n3483) );
  AOI21X1 U2787 ( .A(n4993), .B(n4965), .C(n2091), .Y(n3517) );
  XOR2X1 U2790 ( .A(n3484), .B(n5043), .Y(n2846) );
  OAI21X1 U2791 ( .A(n4968), .B(n4784), .C(n4023), .Y(n3484) );
  AOI21X1 U2792 ( .A(n4991), .B(n4965), .C(n2093), .Y(n3518) );
  XOR2X1 U2795 ( .A(n3485), .B(n5043), .Y(n2847) );
  OAI21X1 U2796 ( .A(n22), .B(n3920), .C(n4022), .Y(n3485) );
  AOI21X1 U2797 ( .A(n4989), .B(n4965), .C(n2095), .Y(n3519) );
  XOR2X1 U2800 ( .A(n3486), .B(n5043), .Y(n2848) );
  OAI21X1 U2801 ( .A(n22), .B(n4802), .C(n4021), .Y(n3486) );
  AOI21X1 U2802 ( .A(n4987), .B(n4965), .C(n2097), .Y(n3520) );
  XOR2X1 U2805 ( .A(n3487), .B(n5043), .Y(n2849) );
  OAI21X1 U2806 ( .A(n22), .B(n4801), .C(n4020), .Y(n3487) );
  AOI21X1 U2807 ( .A(b[3]), .B(n4965), .C(n2099), .Y(n3521) );
  XOR2X1 U2810 ( .A(n3488), .B(n5043), .Y(n2850) );
  OAI21X1 U2811 ( .A(n22), .B(n3922), .C(n4019), .Y(n3488) );
  AOI21X1 U2812 ( .A(b[2]), .B(n4966), .C(n2101), .Y(n3522) );
  XOR2X1 U2815 ( .A(n3489), .B(n5043), .Y(n2851) );
  OAI21X1 U2816 ( .A(n22), .B(n3919), .C(n4018), .Y(n3489) );
  AOI21X1 U2817 ( .A(b[1]), .B(n4966), .C(n2103), .Y(n3523) );
  XOR2X1 U2820 ( .A(n3490), .B(n5043), .Y(n2852) );
  OAI21X1 U2821 ( .A(n22), .B(n4765), .C(n4017), .Y(n3490) );
  AOI21X1 U2822 ( .A(b[0]), .B(n4966), .C(n2105), .Y(n3524) );
  XOR2X1 U2825 ( .A(n3491), .B(n5043), .Y(n2853) );
  OAI21X1 U2826 ( .A(n22), .B(n4359), .C(n3967), .Y(n3491) );
  XOR2X1 U2828 ( .A(n3492), .B(n5043), .Y(n2854) );
  OAI21X1 U2829 ( .A(n22), .B(n4982), .C(n3525), .Y(n3492) );
  AND2X1 U2831 ( .A(n4973), .B(b[0]), .Y(n2107) );
  XOR2X1 U2833 ( .A(n3526), .B(n5038), .Y(n2856) );
  OAI21X1 U2834 ( .A(n4977), .B(n3593), .C(n4639), .Y(n3526) );
  XOR2X1 U2836 ( .A(n3527), .B(n5038), .Y(n2857) );
  OAI21X1 U2837 ( .A(n4977), .B(n4809), .C(n4449), .Y(n3527) );
  AOI21X1 U2838 ( .A(n5033), .B(n4974), .C(n2108), .Y(n3561) );
  AND2X1 U2839 ( .A(n4), .B(n5036), .Y(n2108) );
  XOR2X1 U2840 ( .A(n3528), .B(n5038), .Y(n2858) );
  OAI21X1 U2841 ( .A(n4977), .B(n4779), .C(n4016), .Y(n3528) );
  AOI21X1 U2842 ( .A(n5031), .B(n4974), .C(n2110), .Y(n3562) );
  XOR2X1 U2845 ( .A(n3529), .B(n5038), .Y(n2859) );
  OAI21X1 U2846 ( .A(n4977), .B(n4780), .C(n4015), .Y(n3529) );
  AOI21X1 U2847 ( .A(n5029), .B(n4974), .C(n2112), .Y(n3563) );
  XOR2X1 U2850 ( .A(n3530), .B(n5038), .Y(n2860) );
  OAI21X1 U2851 ( .A(n4977), .B(n4776), .C(n4014), .Y(n3530) );
  AOI21X1 U2852 ( .A(n5027), .B(n4974), .C(n2114), .Y(n3564) );
  XOR2X1 U2855 ( .A(n3531), .B(n5038), .Y(n2861) );
  OAI21X1 U2856 ( .A(n4977), .B(n4769), .C(n4013), .Y(n3531) );
  AOI21X1 U2857 ( .A(n5025), .B(n4974), .C(n2116), .Y(n3565) );
  XOR2X1 U2860 ( .A(n3532), .B(n5038), .Y(n2862) );
  OAI21X1 U2861 ( .A(n4977), .B(n4778), .C(n4012), .Y(n3532) );
  AOI21X1 U2862 ( .A(n5023), .B(n4975), .C(n2118), .Y(n3566) );
  XOR2X1 U2865 ( .A(n3533), .B(n5038), .Y(n2863) );
  OAI21X1 U2866 ( .A(n4977), .B(n3914), .C(n4011), .Y(n3533) );
  AOI21X1 U2867 ( .A(n5021), .B(n4975), .C(n2120), .Y(n3567) );
  XOR2X1 U2870 ( .A(n3534), .B(n5038), .Y(n2864) );
  OAI21X1 U2871 ( .A(n4977), .B(n4767), .C(n4010), .Y(n3534) );
  AOI21X1 U2872 ( .A(n5019), .B(n4975), .C(n2122), .Y(n3568) );
  XOR2X1 U2875 ( .A(n3535), .B(n5039), .Y(n2865) );
  OAI21X1 U2876 ( .A(n4977), .B(n4775), .C(n4009), .Y(n3535) );
  AOI21X1 U2877 ( .A(b[22]), .B(n4975), .C(n2124), .Y(n3569) );
  XOR2X1 U2880 ( .A(n3536), .B(n5039), .Y(n2866) );
  OAI21X1 U2881 ( .A(n9), .B(n4774), .C(n4008), .Y(n3536) );
  AOI21X1 U2882 ( .A(n5017), .B(n4975), .C(n2126), .Y(n3570) );
  XOR2X1 U2885 ( .A(n3537), .B(n5039), .Y(n2867) );
  OAI21X1 U2886 ( .A(n9), .B(n4772), .C(n4007), .Y(n3537) );
  AOI21X1 U2887 ( .A(b[20]), .B(n4975), .C(n2128), .Y(n3571) );
  XOR2X1 U2890 ( .A(n3538), .B(n5039), .Y(n2868) );
  OAI21X1 U2891 ( .A(n4977), .B(n4804), .C(n4006), .Y(n3538) );
  AOI21X1 U2892 ( .A(n5015), .B(n4975), .C(n2130), .Y(n3572) );
  XOR2X1 U2895 ( .A(n3539), .B(n5039), .Y(n2869) );
  OAI21X1 U2896 ( .A(n4977), .B(n4803), .C(n4005), .Y(n3539) );
  AOI21X1 U2897 ( .A(n5013), .B(n4975), .C(n2132), .Y(n3573) );
  XOR2X1 U2900 ( .A(n3540), .B(n5039), .Y(n2870) );
  OAI21X1 U2901 ( .A(n4977), .B(n4766), .C(n4004), .Y(n3540) );
  AOI21X1 U2902 ( .A(b[17]), .B(n4975), .C(n2134), .Y(n3574) );
  XOR2X1 U2905 ( .A(n3541), .B(n5039), .Y(n2871) );
  OAI21X1 U2906 ( .A(n4977), .B(n4773), .C(n4003), .Y(n3541) );
  AOI21X1 U2907 ( .A(n5011), .B(n4975), .C(n2136), .Y(n3575) );
  XOR2X1 U2910 ( .A(n3542), .B(n5039), .Y(n2872) );
  OAI21X1 U2911 ( .A(n4977), .B(n4768), .C(n4002), .Y(n3542) );
  AOI21X1 U2912 ( .A(n5009), .B(n4974), .C(n2138), .Y(n3576) );
  XOR2X1 U2915 ( .A(n3543), .B(n5039), .Y(n2873) );
  OAI21X1 U2916 ( .A(n4977), .B(n3923), .C(n4001), .Y(n3543) );
  AOI21X1 U2917 ( .A(n5007), .B(n4974), .C(n2140), .Y(n3577) );
  XOR2X1 U2920 ( .A(n3544), .B(n5039), .Y(n2874) );
  OAI21X1 U2921 ( .A(n4977), .B(n4783), .C(n4000), .Y(n3544) );
  AOI21X1 U2922 ( .A(n5005), .B(n4974), .C(n2142), .Y(n3578) );
  XOR2X1 U2925 ( .A(n3545), .B(n5039), .Y(n2875) );
  OAI21X1 U2926 ( .A(n4977), .B(n3917), .C(n3999), .Y(n3545) );
  AOI21X1 U2927 ( .A(n5003), .B(n4974), .C(n2144), .Y(n3579) );
  XOR2X1 U2930 ( .A(n3546), .B(n5039), .Y(n2876) );
  OAI21X1 U2931 ( .A(n4977), .B(n3913), .C(n3998), .Y(n3546) );
  AOI21X1 U2932 ( .A(n5001), .B(n4974), .C(n2146), .Y(n3580) );
  XOR2X1 U2935 ( .A(n3547), .B(n5039), .Y(n2877) );
  OAI21X1 U2936 ( .A(n4977), .B(n3918), .C(n3997), .Y(n3547) );
  AOI21X1 U2937 ( .A(n4999), .B(n4974), .C(n2148), .Y(n3581) );
  XOR2X1 U2940 ( .A(n3548), .B(n5038), .Y(n2878) );
  OAI21X1 U2941 ( .A(n4977), .B(n4782), .C(n3996), .Y(n3548) );
  AOI21X1 U2942 ( .A(n4997), .B(n4974), .C(n2150), .Y(n3582) );
  XOR2X1 U2945 ( .A(n3549), .B(n5038), .Y(n2879) );
  OAI21X1 U2946 ( .A(n4977), .B(n3916), .C(n3995), .Y(n3549) );
  AOI21X1 U2947 ( .A(n4995), .B(n4974), .C(n2152), .Y(n3583) );
  XOR2X1 U2950 ( .A(n3550), .B(n5038), .Y(n2880) );
  OAI21X1 U2951 ( .A(n4977), .B(n3921), .C(n3994), .Y(n3550) );
  AOI21X1 U2952 ( .A(n4993), .B(n4974), .C(n2154), .Y(n3584) );
  XOR2X1 U2955 ( .A(n3551), .B(n5038), .Y(n2881) );
  OAI21X1 U2956 ( .A(n4977), .B(n4784), .C(n3993), .Y(n3551) );
  AOI21X1 U2957 ( .A(n4991), .B(n4974), .C(n2156), .Y(n3585) );
  XOR2X1 U2960 ( .A(n3552), .B(n5038), .Y(n2882) );
  OAI21X1 U2961 ( .A(n4977), .B(n3920), .C(n3992), .Y(n3552) );
  AOI21X1 U2962 ( .A(n4989), .B(n4974), .C(n2158), .Y(n3586) );
  XOR2X1 U2965 ( .A(n3553), .B(n5038), .Y(n2883) );
  OAI21X1 U2966 ( .A(n4977), .B(n4802), .C(n3991), .Y(n3553) );
  AOI21X1 U2967 ( .A(n4987), .B(n4974), .C(n2160), .Y(n3587) );
  XOR2X1 U2970 ( .A(n3554), .B(n5038), .Y(n2884) );
  OAI21X1 U2971 ( .A(n4977), .B(n4801), .C(n3990), .Y(n3554) );
  AOI21X1 U2972 ( .A(b[3]), .B(n4974), .C(n2162), .Y(n3588) );
  XOR2X1 U2975 ( .A(n3555), .B(n5038), .Y(n2885) );
  OAI21X1 U2976 ( .A(n9), .B(n3922), .C(n3989), .Y(n3555) );
  AOI21X1 U2977 ( .A(n4983), .B(n4975), .C(n2164), .Y(n3589) );
  XOR2X1 U2980 ( .A(n3556), .B(n5038), .Y(n2886) );
  OAI21X1 U2981 ( .A(n9), .B(n3919), .C(n3988), .Y(n3556) );
  AOI21X1 U2982 ( .A(b[1]), .B(n4975), .C(n2166), .Y(n3590) );
  OAI21X1 U2986 ( .A(n9), .B(n4765), .C(n3987), .Y(n3557) );
  AOI21X1 U2987 ( .A(b[0]), .B(n4975), .C(n2168), .Y(n3591) );
  XOR2X1 U2990 ( .A(n3558), .B(n5038), .Y(n754) );
  OAI21X1 U2991 ( .A(n9), .B(n4359), .C(n3966), .Y(n3558) );
  XOR2X1 U2993 ( .A(n3559), .B(n5038), .Y(n2889) );
  OAI21X1 U2994 ( .A(n9), .B(n4982), .C(n3592), .Y(n3559) );
  AND2X1 U2996 ( .A(n4979), .B(n4981), .Y(n2170) );
  AND2X1 U3073 ( .A(a[31]), .B(n2171), .Y(n129) );
  OR2X1 U3075 ( .A(n3692), .B(n2172), .Y(n127) );
  AND2X1 U3077 ( .A(n3692), .B(n2173), .Y(n124) );
  XNOR2X1 U3080 ( .A(a[30]), .B(a[31]), .Y(n3703) );
  XNOR2X1 U3081 ( .A(a[29]), .B(a[30]), .Y(n3692) );
  OR2X1 U3084 ( .A(n3693), .B(n2175), .Y(n118) );
  XNOR2X1 U3089 ( .A(a[27]), .B(a[28]), .Y(n3704) );
  XNOR2X1 U3090 ( .A(a[26]), .B(a[27]), .Y(n3693) );
  XOR2X1 U3091 ( .A(a[29]), .B(a[28]), .Y(n3715) );
  AND2X1 U3092 ( .A(n3705), .B(n2177), .Y(n108) );
  OR2X1 U3094 ( .A(n3694), .B(n2178), .Y(n106) );
  AND2X1 U3096 ( .A(n3694), .B(n2179), .Y(n100) );
  XNOR2X1 U3099 ( .A(a[25]), .B(a[24]), .Y(n3705) );
  XNOR2X1 U3100 ( .A(a[23]), .B(a[24]), .Y(n3694) );
  XOR2X1 U3101 ( .A(a[26]), .B(a[25]), .Y(n3716) );
  AND2X1 U3102 ( .A(n3706), .B(n2180), .Y(n96) );
  OR2X1 U3104 ( .A(n3695), .B(n2181), .Y(n94) );
  AND2X1 U3106 ( .A(n3695), .B(n2182), .Y(n88) );
  XNOR2X1 U3109 ( .A(a[22]), .B(a[21]), .Y(n3706) );
  XNOR2X1 U3110 ( .A(a[20]), .B(a[21]), .Y(n3695) );
  XOR2X1 U3111 ( .A(a[23]), .B(a[22]), .Y(n3717) );
  AND2X1 U3112 ( .A(n3707), .B(n2183), .Y(n84) );
  OR2X1 U3114 ( .A(n3696), .B(n2184), .Y(n82) );
  AND2X1 U3116 ( .A(n3696), .B(n2185), .Y(n76) );
  XNOR2X1 U3119 ( .A(a[19]), .B(a[18]), .Y(n3707) );
  XNOR2X1 U3120 ( .A(a[17]), .B(a[18]), .Y(n3696) );
  XOR2X1 U3121 ( .A(a[20]), .B(a[19]), .Y(n3718) );
  AND2X1 U3122 ( .A(n3708), .B(n2186), .Y(n72) );
  OR2X1 U3124 ( .A(n3697), .B(n2187), .Y(n70) );
  XNOR2X1 U3129 ( .A(a[15]), .B(a[16]), .Y(n3708) );
  XNOR2X1 U3130 ( .A(a[14]), .B(a[15]), .Y(n3697) );
  XOR2X1 U3131 ( .A(a[17]), .B(a[16]), .Y(n3719) );
  OR2X1 U3134 ( .A(n3698), .B(n2190), .Y(n58) );
  XNOR2X1 U3139 ( .A(a[13]), .B(a[12]), .Y(n3709) );
  XNOR2X1 U3140 ( .A(a[11]), .B(a[12]), .Y(n3698) );
  XOR2X1 U3141 ( .A(a[14]), .B(a[13]), .Y(n3720) );
  AND2X1 U3142 ( .A(n3710), .B(n2192), .Y(n48) );
  OR2X1 U3144 ( .A(n3699), .B(n2193), .Y(n46) );
  AND2X1 U3146 ( .A(n3699), .B(n2194), .Y(n40) );
  XNOR2X1 U3149 ( .A(a[9]), .B(a[10]), .Y(n3710) );
  XNOR2X1 U3150 ( .A(a[8]), .B(a[9]), .Y(n3699) );
  XOR2X1 U3151 ( .A(a[11]), .B(a[10]), .Y(n3721) );
  AND2X1 U3152 ( .A(n3711), .B(n2195), .Y(n36) );
  OR2X1 U3154 ( .A(n3700), .B(n2196), .Y(n34) );
  AND2X1 U3156 ( .A(n3700), .B(n2197), .Y(n28) );
  XNOR2X1 U3159 ( .A(a[7]), .B(a[6]), .Y(n3711) );
  XNOR2X1 U3160 ( .A(a[5]), .B(a[6]), .Y(n3700) );
  XOR2X1 U3161 ( .A(a[8]), .B(a[7]), .Y(n3722) );
  AND2X1 U3162 ( .A(n3712), .B(n2198), .Y(n24) );
  OR2X1 U3164 ( .A(n3701), .B(n2199), .Y(n22) );
  AND2X1 U3166 ( .A(n3701), .B(n2200), .Y(n16) );
  XNOR2X1 U3169 ( .A(a[4]), .B(a[3]), .Y(n3712) );
  XNOR2X1 U3170 ( .A(n5039), .B(a[3]), .Y(n3701) );
  XOR2X1 U3171 ( .A(a[5]), .B(a[4]), .Y(n3723) );
  AND2X1 U3172 ( .A(n3702), .B(n4342), .Y(n12) );
  OR2X1 U3174 ( .A(n3702), .B(n2202), .Y(n9) );
  XOR2X1 U3181 ( .A(n5039), .B(a[1]), .Y(n3724) );
  OAI21X1 U3188 ( .A(n3956), .B(n3955), .C(n3947), .Y(n2238) );
  AOI21X1 U3190 ( .A(n2326), .B(n4407), .C(n2242), .Y(n2240) );
  OAI21X1 U3192 ( .A(n4411), .B(n4428), .C(n3986), .Y(n2242) );
  AOI21X1 U3194 ( .A(n2266), .B(n4515), .C(n2246), .Y(n2244) );
  OAI21X1 U3196 ( .A(n4683), .B(n4622), .C(n4544), .Y(n2246) );
  AOI21X1 U3202 ( .A(n2396), .B(n4350), .C(n2251), .Y(n2249) );
  OAI21X1 U3204 ( .A(n3944), .B(n2328), .C(n3985), .Y(n2251) );
  AOI21X1 U3206 ( .A(n4427), .B(n4554), .C(n2255), .Y(n2253) );
  OAI21X1 U3208 ( .A(n4756), .B(n2268), .C(n4683), .Y(n2255) );
  AOI21X1 U3216 ( .A(n2396), .B(n3950), .C(n2262), .Y(n2260) );
  OAI21X1 U3218 ( .A(n4416), .B(n2328), .C(n3984), .Y(n2262) );
  AOI21X1 U3220 ( .A(n4427), .B(n4687), .C(n2266), .Y(n2264) );
  OAI21X1 U3226 ( .A(n4561), .B(n4626), .C(n4510), .Y(n2266) );
  AOI21X1 U3232 ( .A(n2396), .B(n3943), .C(n2275), .Y(n2273) );
  OAI21X1 U3234 ( .A(n4415), .B(n2328), .C(n3983), .Y(n2275) );
  AOI21X1 U3236 ( .A(n4427), .B(n2280), .C(n2281), .Y(n2277) );
  AOI21X1 U3244 ( .A(n2396), .B(n4349), .C(n2284), .Y(n2282) );
  OAI21X1 U3246 ( .A(n4442), .B(n2328), .C(n4428), .Y(n2284) );
  AOI21X1 U3252 ( .A(n2310), .B(n3962), .C(n2292), .Y(n2286) );
  OAI21X1 U3254 ( .A(n4674), .B(n4745), .C(n4603), .Y(n2292) );
  AOI21X1 U3260 ( .A(n2396), .B(n4348), .C(n2297), .Y(n2295) );
  OAI21X1 U3262 ( .A(n4414), .B(n2328), .C(n3982), .Y(n2297) );
  AOI21X1 U3264 ( .A(n2310), .B(n2302), .C(n2303), .Y(n2299) );
  AOI21X1 U3272 ( .A(n2396), .B(n4347), .C(n2306), .Y(n2304) );
  OAI21X1 U3274 ( .A(n2309), .B(n2328), .C(n2308), .Y(n2306) );
  OAI21X1 U3282 ( .A(n4682), .B(n4627), .C(n4543), .Y(n2310) );
  AOI21X1 U3288 ( .A(n2396), .B(n4346), .C(n2319), .Y(n2317) );
  OAI21X1 U3290 ( .A(n4755), .B(n2328), .C(n4682), .Y(n2319) );
  AOI21X1 U3298 ( .A(n2396), .B(n4424), .C(n2326), .Y(n2324) );
  OAI21X1 U3304 ( .A(n4412), .B(n4439), .C(n3981), .Y(n2326) );
  AOI21X1 U3306 ( .A(n2352), .B(n4404), .C(n2334), .Y(n2332) );
  OAI21X1 U3308 ( .A(n4436), .B(n4429), .C(n4398), .Y(n2334) );
  AOI21X1 U3314 ( .A(n2396), .B(n4345), .C(n2339), .Y(n2337) );
  OAI21X1 U3316 ( .A(n4441), .B(n4400), .C(n4436), .Y(n2339) );
  AOI21X1 U3324 ( .A(n2396), .B(n2347), .C(n4399), .Y(n2344) );
  AOI21X1 U3328 ( .A(n4438), .B(n4437), .C(n2352), .Y(n2348) );
  OAI21X1 U3332 ( .A(n4435), .B(n4431), .C(n4397), .Y(n2352) );
  AOI21X1 U3338 ( .A(n2396), .B(n4344), .C(n2357), .Y(n2355) );
  OAI21X1 U3340 ( .A(n4754), .B(n4439), .C(n4435), .Y(n2357) );
  AOI21X1 U3348 ( .A(n2396), .B(n2365), .C(n4438), .Y(n2362) );
  AOI21X1 U3356 ( .A(n2384), .B(n4406), .C(n2372), .Y(n2366) );
  OAI21X1 U3358 ( .A(n4434), .B(n4432), .C(n4396), .Y(n2372) );
  AOI21X1 U3364 ( .A(n2396), .B(n4343), .C(n2377), .Y(n2375) );
  OAI21X1 U3366 ( .A(n4440), .B(n2386), .C(n4434), .Y(n2377) );
  AOI21X1 U3374 ( .A(n2396), .B(n4423), .C(n2384), .Y(n2382) );
  OAI21X1 U3380 ( .A(n4673), .B(n4747), .C(n4600), .Y(n2384) );
  AOI21X1 U3386 ( .A(n2396), .B(n2394), .C(n2395), .Y(n2391) );
  AOI21X1 U3395 ( .A(n2452), .B(n3949), .C(n2399), .Y(n2397) );
  OAI21X1 U3397 ( .A(n4410), .B(n4426), .C(n3980), .Y(n2399) );
  AOI21X1 U3399 ( .A(n2417), .B(n4403), .C(n2403), .Y(n2401) );
  OAI21X1 U3401 ( .A(n4675), .B(n4741), .C(n4604), .Y(n2403) );
  AOI21X1 U3407 ( .A(n2411), .B(n2409), .C(n2410), .Y(n2406) );
  OAI21X1 U3415 ( .A(n4353), .B(n2451), .C(n3979), .Y(n2411) );
  AOI21X1 U3417 ( .A(n4425), .B(n4686), .C(n2417), .Y(n2413) );
  OAI21X1 U3421 ( .A(n4672), .B(n4748), .C(n4601), .Y(n2417) );
  AOI21X1 U3427 ( .A(n2425), .B(n2423), .C(n2424), .Y(n2420) );
  OAI21X1 U3435 ( .A(n4430), .B(n2451), .C(n4426), .Y(n2425) );
  AOI21X1 U3441 ( .A(n2445), .B(n3963), .C(n2433), .Y(n2427) );
  OAI21X1 U3443 ( .A(n4676), .B(n4750), .C(n4605), .Y(n2433) );
  AOI21X1 U3449 ( .A(n2441), .B(n2439), .C(n2440), .Y(n2436) );
  OAI21X1 U3457 ( .A(n2444), .B(n2451), .C(n2443), .Y(n2441) );
  OAI21X1 U3461 ( .A(n4684), .B(n4749), .C(n4548), .Y(n2445) );
  OAI21X1 U3467 ( .A(n4620), .B(n2451), .C(n4684), .Y(n2448) );
  OAI21X1 U3474 ( .A(n4352), .B(n4513), .C(n3978), .Y(n2452) );
  AOI21X1 U3476 ( .A(n2464), .B(n4408), .C(n2456), .Y(n2454) );
  OAI21X1 U3478 ( .A(n4433), .B(n4744), .C(n4395), .Y(n2456) );
  OAI21X1 U3484 ( .A(n4679), .B(n4421), .C(n4433), .Y(n2459) );
  AOI21X1 U3490 ( .A(n2472), .B(n4405), .C(n2464), .Y(n2462) );
  OAI21X1 U3492 ( .A(n4671), .B(n4746), .C(n4602), .Y(n2464) );
  AOI21X1 U3498 ( .A(n2472), .B(n2470), .C(n2471), .Y(n2467) );
  AOI21X1 U3507 ( .A(n4514), .B(n2481), .C(n2475), .Y(n2473) );
  OAI21X1 U3509 ( .A(n4685), .B(n4562), .C(n4481), .Y(n2475) );
  OAI21X1 U3515 ( .A(n4624), .B(n4757), .C(n4685), .Y(n2478) );
  DFFPOSX1 clk_r_REG11_S1 ( .D(n4821), .CLK(ALU1ALU_MUL32_CLK), .Q(n4919) );
  DFFPOSX1 clk_r_REG48_S1 ( .D(n4787), .CLK(ALU1ALU_MUL32_CLK), .Q(n4918) );
  DFFPOSX1 clk_r_REG46_S1 ( .D(n4800), .CLK(ALU1ALU_MUL32_CLK), .Q(n4917) );
  DFFPOSX1 clk_r_REG44_S1 ( .D(n4799), .CLK(ALU1ALU_MUL32_CLK), .Q(n4916) );
  DFFPOSX1 clk_r_REG42_S1 ( .D(n4786), .CLK(ALU1ALU_MUL32_CLK), .Q(n4915) );
  DFFPOSX1 clk_r_REG32_S1 ( .D(n4785), .CLK(ALU1ALU_MUL32_CLK), .Q(n4914) );
  DFFPOSX1 clk_r_REG30_S1 ( .D(n4798), .CLK(ALU1ALU_MUL32_CLK), .Q(n4913) );
  DFFPOSX1 clk_r_REG28_S1 ( .D(n4797), .CLK(ALU1ALU_MUL32_CLK), .Q(n4912) );
  DFFPOSX1 clk_r_REG26_S1 ( .D(n4796), .CLK(ALU1ALU_MUL32_CLK), .Q(n4911) );
  DFFPOSX1 clk_r_REG38_S1 ( .D(n4795), .CLK(ALU1ALU_MUL32_CLK), .Q(n4910) );
  DFFPOSX1 clk_r_REG36_S1 ( .D(n4794), .CLK(ALU1ALU_MUL32_CLK), .Q(n4909) );
  DFFPOSX1 clk_r_REG70_S1 ( .D(n4793), .CLK(ALU1ALU_MUL32_CLK), .Q(n4908) );
  DFFPOSX1 clk_r_REG72_S1 ( .D(n4792), .CLK(ALU1ALU_MUL32_CLK), .Q(n4907) );
  DFFPOSX1 clk_r_REG74_S1 ( .D(n4791), .CLK(ALU1ALU_MUL32_CLK), .Q(n4906) );
  DFFPOSX1 clk_r_REG76_S1 ( .D(n4790), .CLK(ALU1ALU_MUL32_CLK), .Q(n4905) );
  DFFPOSX1 clk_r_REG78_S1 ( .D(n4789), .CLK(ALU1ALU_MUL32_CLK), .Q(n4904) );
  DFFPOSX1 clk_r_REG82_S1 ( .D(n4788), .CLK(ALU1ALU_MUL32_CLK), .Q(n4903) );
  DFFPOSX1 clk_r_REG68_S1 ( .D(n232), .CLK(ALU1ALU_MUL32_CLK), .Q(n4902) );
  DFFPOSX1 clk_r_REG10_S1 ( .D(n4690), .CLK(ALU1ALU_MUL32_CLK), .Q(n4901) );
  DFFPOSX1 clk_r_REG9_S1 ( .D(n4564), .CLK(ALU1ALU_MUL32_CLK), .Q(n4900) );
  DFFPOSX1 clk_r_REG8_S1 ( .D(n4517), .CLK(ALU1ALU_MUL32_CLK), .Q(n4899) );
  DFFPOSX1 clk_r_REG7_S1 ( .D(n4629), .CLK(ALU1ALU_MUL32_CLK), .Q(n4898) );
  DFFPOSX1 clk_r_REG6_S1 ( .D(n4465), .CLK(ALU1ALU_MUL32_CLK), .Q(n4897) );
  DFFPOSX1 clk_r_REG5_S1 ( .D(n4518), .CLK(ALU1ALU_MUL32_CLK), .Q(n4896) );
  DFFPOSX1 clk_r_REG4_S1 ( .D(n4691), .CLK(ALU1ALU_MUL32_CLK), .Q(n4895) );
  DFFPOSX1 clk_r_REG3_S1 ( .D(n4630), .CLK(ALU1ALU_MUL32_CLK), .Q(n4894) );
  DFFPOSX1 clk_r_REG2_S1 ( .D(n4563), .CLK(ALU1ALU_MUL32_CLK), .Q(n4893) );
  DFFPOSX1 clk_r_REG1_S1 ( .D(n4519), .CLK(ALU1ALU_MUL32_CLK), .Q(n4892) );
  DFFPOSX1 clk_r_REG0_S1 ( .D(n4483), .CLK(ALU1ALU_MUL32_CLK), .Q(n4891) );
  DFFPOSX1 clk_r_REG50_S1 ( .D(n4692), .CLK(ALU1ALU_MUL32_CLK), .Q(n4890) );
  DFFPOSX1 clk_r_REG49_S1 ( .D(n4565), .CLK(ALU1ALU_MUL32_CLK), .Q(n4889) );
  DFFPOSX1 clk_r_REG47_S1 ( .D(n4631), .CLK(ALU1ALU_MUL32_CLK), .Q(n4888) );
  DFFPOSX1 clk_r_REG45_S1 ( .D(n4694), .CLK(ALU1ALU_MUL32_CLK), .Q(n4887) );
  DFFPOSX1 clk_r_REG43_S1 ( .D(n4566), .CLK(ALU1ALU_MUL32_CLK), .Q(n4886) );
  DFFPOSX1 clk_r_REG41_S1 ( .D(n4632), .CLK(ALU1ALU_MUL32_CLK), .Q(n4885) );
  DFFPOSX1 clk_r_REG40_S1 ( .D(n4569), .CLK(ALU1ALU_MUL32_CLK), .Q(n4884) );
  DFFPOSX1 clk_r_REG39_S1 ( .D(n4697), .CLK(ALU1ALU_MUL32_CLK), .Q(n4883) );
  DFFPOSX1 clk_r_REG34_S1 ( .D(n4635), .CLK(ALU1ALU_MUL32_CLK), .Q(n4882) );
  DFFPOSX1 clk_r_REG33_S1 ( .D(n4522), .CLK(ALU1ALU_MUL32_CLK), .Q(n4881) );
  DFFPOSX1 clk_r_REG31_S1 ( .D(n4702), .CLK(ALU1ALU_MUL32_CLK), .Q(n4880) );
  DFFPOSX1 clk_r_REG29_S1 ( .D(n4523), .CLK(ALU1ALU_MUL32_CLK), .Q(n4879) );
  DFFPOSX1 clk_r_REG27_S1 ( .D(n4696), .CLK(ALU1ALU_MUL32_CLK), .Q(n4878) );
  DFFPOSX1 clk_r_REG25_S1 ( .D(n4568), .CLK(ALU1ALU_MUL32_CLK), .Q(n4877) );
  DFFPOSX1 clk_r_REG37_S1 ( .D(n4693), .CLK(ALU1ALU_MUL32_CLK), .Q(n4876) );
  DFFPOSX1 clk_r_REG35_S1 ( .D(n4521), .CLK(ALU1ALU_MUL32_CLK), .Q(n4875) );
  DFFPOSX1 clk_r_REG67_S1 ( .D(n4699), .CLK(ALU1ALU_MUL32_CLK), .Q(n4874) );
  DFFPOSX1 clk_r_REG66_S1 ( .D(n4571), .CLK(ALU1ALU_MUL32_CLK), .Q(n4873) );
  DFFPOSX1 clk_r_REG23_S1 ( .D(n4700), .CLK(ALU1ALU_MUL32_CLK), .Q(n4872) );
  DFFPOSX1 clk_r_REG22_S1 ( .D(n4572), .CLK(ALU1ALU_MUL32_CLK), .Q(n4871) );
  DFFPOSX1 clk_r_REG19_S1 ( .D(n4524), .CLK(ALU1ALU_MUL32_CLK), .Q(n4870) );
  DFFPOSX1 clk_r_REG18_S1 ( .D(n4576), .CLK(ALU1ALU_MUL32_CLK), .Q(n4869) );
  DFFPOSX1 clk_r_REG17_S1 ( .D(n4638), .CLK(ALU1ALU_MUL32_CLK), .Q(n4868) );
  DFFPOSX1 clk_r_REG16_S1 ( .D(n4703), .CLK(ALU1ALU_MUL32_CLK), .Q(n4867) );
  DFFPOSX1 clk_r_REG15_S1 ( .D(n4525), .CLK(ALU1ALU_MUL32_CLK), .Q(n4866) );
  DFFPOSX1 clk_r_REG14_S1 ( .D(n4575), .CLK(ALU1ALU_MUL32_CLK), .Q(n4865) );
  DFFPOSX1 clk_r_REG13_S1 ( .D(n4637), .CLK(ALU1ALU_MUL32_CLK), .Q(n4864) );
  DFFPOSX1 clk_r_REG12_S1 ( .D(n4485), .CLK(ALU1ALU_MUL32_CLK), .Q(n4863) );
  DFFPOSX1 clk_r_REG69_S1 ( .D(n4574), .CLK(ALU1ALU_MUL32_CLK), .Q(n4862) );
  DFFPOSX1 clk_r_REG71_S1 ( .D(n4636), .CLK(ALU1ALU_MUL32_CLK), .Q(n4861) );
  DFFPOSX1 clk_r_REG73_S1 ( .D(n4701), .CLK(ALU1ALU_MUL32_CLK), .Q(n4860) );
  DFFPOSX1 clk_r_REG75_S1 ( .D(n4573), .CLK(ALU1ALU_MUL32_CLK), .Q(n4859) );
  DFFPOSX1 clk_r_REG77_S1 ( .D(n4634), .CLK(ALU1ALU_MUL32_CLK), .Q(n4858) );
  DFFPOSX1 clk_r_REG80_S1 ( .D(n4698), .CLK(ALU1ALU_MUL32_CLK), .Q(n4857) );
  DFFPOSX1 clk_r_REG79_S1 ( .D(n4570), .CLK(ALU1ALU_MUL32_CLK), .Q(n4856) );
  DFFPOSX1 clk_r_REG81_S1 ( .D(n4520), .CLK(ALU1ALU_MUL32_CLK), .Q(n4855) );
  DFFPOSX1 clk_r_REG84_S1 ( .D(n4484), .CLK(ALU1ALU_MUL32_CLK), .Q(n4854) );
  DFFPOSX1 clk_r_REG83_S1 ( .D(n4567), .CLK(ALU1ALU_MUL32_CLK), .Q(n4853) );
  DFFPOSX1 clk_r_REG86_S1 ( .D(n4633), .CLK(ALU1ALU_MUL32_CLK), .Q(n4852) );
  DFFPOSX1 clk_r_REG85_S1 ( .D(n4695), .CLK(ALU1ALU_MUL32_CLK), .Q(n4851) );
  DFFPOSX1 clk_r_REG87_S1 ( .D(n3965), .CLK(ALU1ALU_MUL32_CLK), .Q(n4850) );
  DFFPOSX1 clk_r_REG88_S1 ( .D(n3964), .CLK(ALU1ALU_MUL32_CLK), .Q(n4849) );
  DFFPOSX1 clk_r_REG90_S1 ( .D(n658), .CLK(ALU1ALU_MUL32_CLK), .Q(n4848) );
  DFFPOSX1 clk_r_REG65_S1 ( .D(n982), .CLK(ALU1ALU_MUL32_CLK), .Q(n4847) );
  DFFPOSX1 clk_r_REG63_S1 ( .D(n997), .CLK(ALU1ALU_MUL32_CLK), .Q(n4846) );
  DFFPOSX1 clk_r_REG64_S1 ( .D(n998), .CLK(ALU1ALU_MUL32_CLK), .Q(n4845) );
  DFFPOSX1 clk_r_REG61_S1 ( .D(n1013), .CLK(ALU1ALU_MUL32_CLK), .Q(n4844) );
  DFFPOSX1 clk_r_REG62_S1 ( .D(n1014), .CLK(ALU1ALU_MUL32_CLK), .Q(n4843) );
  DFFPOSX1 clk_r_REG58_S1 ( .D(n1029), .CLK(ALU1ALU_MUL32_CLK), .Q(n4842) );
  DFFPOSX1 clk_r_REG59_S1 ( .D(n1030), .CLK(ALU1ALU_MUL32_CLK), .Q(n4841) );
  DFFPOSX1 clk_r_REG57_S1 ( .D(n1050), .CLK(ALU1ALU_MUL32_CLK), .Q(n4840) );
  DFFPOSX1 clk_r_REG60_S1 ( .D(n1052), .CLK(ALU1ALU_MUL32_CLK), .Q(n4839) );
  DFFPOSX1 clk_r_REG54_S1 ( .D(n1066), .CLK(ALU1ALU_MUL32_CLK), .Q(n4838) );
  DFFPOSX1 clk_r_REG55_S1 ( .D(n1067), .CLK(ALU1ALU_MUL32_CLK), .Q(n4837) );
  DFFPOSX1 clk_r_REG56_S1 ( .D(n1069), .CLK(ALU1ALU_MUL32_CLK), .Q(n4836) );
  DFFPOSX1 clk_r_REG51_S1 ( .D(n1082), .CLK(ALU1ALU_MUL32_CLK), .Q(n4835) );
  DFFPOSX1 clk_r_REG52_S1 ( .D(n1083), .CLK(ALU1ALU_MUL32_CLK), .Q(n4834) );
  DFFPOSX1 clk_r_REG53_S1 ( .D(n1084), .CLK(ALU1ALU_MUL32_CLK), .Q(n4833) );
  DFFPOSX1 clk_r_REG24_S1 ( .D(n1100), .CLK(ALU1ALU_MUL32_CLK), .Q(n4832) );
  DFFPOSX1 clk_r_REG21_S1 ( .D(n1119), .CLK(ALU1ALU_MUL32_CLK), .Q(n4831) );
  DFFPOSX1 clk_r_REG20_S1 ( .D(n1136), .CLK(ALU1ALU_MUL32_CLK), .Q(n4830) );
  AND2X2 U3530 ( .A(n3697), .B(n2188), .Y(n64) );
  OR2X2 U3531 ( .A(n5036), .B(b[30]), .Y(n2247) );
  AND2X2 U3532 ( .A(n5036), .B(n2238), .Y(n4771) );
  INVX2 U3533 ( .A(n5037), .Y(n5036) );
  AND2X2 U3534 ( .A(n533), .B(n528), .Y(n3925) );
  AND2X2 U3535 ( .A(n3704), .B(n2174), .Y(n120) );
  INVX2 U3536 ( .A(n3956), .Y(n2396) );
  INVX2 U3537 ( .A(n5041), .Y(n5039) );
  AND2X2 U3538 ( .A(n3702), .B(n3924), .Y(n4) );
  INVX2 U3539 ( .A(n4813), .Y(n4944) );
  OR2X2 U3540 ( .A(n3719), .B(n3697), .Y(n4813) );
  AND2X2 U3541 ( .A(n3698), .B(n2191), .Y(n52) );
  AND2X2 U3542 ( .A(n765), .B(n4560), .Y(n357) );
  AND2X2 U3543 ( .A(n3709), .B(n2189), .Y(n60) );
  AND2X2 U3544 ( .A(n3698), .B(n3720), .Y(n2189) );
  AND2X1 U3545 ( .A(n4914), .B(n4731), .Y(n424) );
  OR2X1 U3546 ( .A(n4540), .B(n4614), .Y(n475) );
  OR2X1 U3547 ( .A(n4896), .B(n4894), .Y(n330) );
  OR2X1 U3548 ( .A(n4394), .B(n4900), .Y(n308) );
  AND2X1 U3549 ( .A(n4503), .B(n4553), .Y(n550) );
  OR2X1 U3550 ( .A(n4506), .B(n4750), .Y(n2432) );
  OR2X1 U3551 ( .A(n4868), .B(n4866), .Y(n579) );
  AND2X1 U3552 ( .A(n1047), .B(n4841), .Y(n534) );
  AND2X1 U3553 ( .A(n400), .B(n4688), .Y(n396) );
  AND2X1 U3554 ( .A(n4628), .B(n4688), .Y(n368) );
  AND2X1 U3555 ( .A(n763), .B(n3961), .Y(n335) );
  AND2X1 U3556 ( .A(n4686), .B(n2426), .Y(n2412) );
  OR2X1 U3557 ( .A(n4754), .B(n4431), .Y(n2349) );
  AND2X1 U3558 ( .A(n2280), .B(n2285), .Y(n2276) );
  AND2X1 U3559 ( .A(n4853), .B(n799), .Y(n273) );
  AND2X1 U3560 ( .A(n4855), .B(n4903), .Y(n272) );
  AND2X1 U3561 ( .A(n4860), .B(n4906), .Y(n268) );
  AND2X1 U3562 ( .A(n4862), .B(n4908), .Y(n266) );
  OR2X1 U3563 ( .A(n4508), .B(n4864), .Y(n587) );
  AND2X1 U3564 ( .A(n4830), .B(n4831), .Y(n571) );
  AND2X1 U3565 ( .A(n4832), .B(n4834), .Y(n559) );
  AND2X1 U3566 ( .A(n326), .B(n4560), .Y(n324) );
  AND2X1 U3567 ( .A(b[24]), .B(b[25]), .Y(n2316) );
  AND2X1 U3568 ( .A(n4687), .B(n2285), .Y(n2263) );
  AND2X1 U3569 ( .A(n4686), .B(n4403), .Y(n2400) );
  OR2X1 U3570 ( .A(n4410), .B(n4430), .Y(n2398) );
  AND2X1 U3571 ( .A(b[24]), .B(b[23]), .Y(n2323) );
  OR2X1 U3572 ( .A(n2325), .B(n4442), .Y(n2283) );
  AND2X1 U3573 ( .A(n2285), .B(n4554), .Y(n2252) );
  INVX1 U3574 ( .A(n2326), .Y(n2328) );
  AND2X1 U3575 ( .A(n4851), .B(n800), .Y(n274) );
  AND2X1 U3576 ( .A(n4859), .B(n4905), .Y(n269) );
  AND2X1 U3577 ( .A(n4599), .B(n570), .Y(n261) );
  AND2X1 U3578 ( .A(n4606), .B(n558), .Y(n259) );
  AND2X1 U3579 ( .A(n4739), .B(n3935), .Y(n258) );
  AND2X1 U3580 ( .A(n4549), .B(n783), .Y(n257) );
  INVX1 U3581 ( .A(n5010), .Y(n5009) );
  AND2X1 U3582 ( .A(n3693), .B(n2176), .Y(n112) );
  AND2X1 U3583 ( .A(n4424), .B(n4407), .Y(n2239) );
  AND2X1 U3584 ( .A(n4867), .B(n789), .Y(n263) );
  AND2X1 U3585 ( .A(n4805), .B(n4808), .Y(n663) );
  OR2X1 U3586 ( .A(n4740), .B(n4613), .Y(n676) );
  INVX2 U3587 ( .A(n4771), .Y(n3593) );
  AND2X1 U3588 ( .A(n5039), .B(n2889), .Y(n758) );
  OR2X1 U3589 ( .A(n4827), .B(n4616), .Y(n751) );
  AND2X1 U3590 ( .A(n1244), .B(n1227), .Y(n604) );
  AND2X1 U3591 ( .A(n1226), .B(n1209), .Y(n599) );
  AND2X1 U3592 ( .A(n1208), .B(n1191), .Y(n590) );
  OR2X1 U3593 ( .A(n1191), .B(n1208), .Y(n589) );
  AND2X1 U3594 ( .A(n1190), .B(n1173), .Y(n585) );
  OR2X1 U3595 ( .A(n1173), .B(n1190), .Y(n584) );
  OR2X1 U3596 ( .A(n1155), .B(n1172), .Y(n581) );
  AND2X1 U3597 ( .A(n1154), .B(n1137), .Y(n574) );
  OR2X1 U3598 ( .A(n1137), .B(n1154), .Y(n573) );
  AND2X1 U3599 ( .A(n1118), .B(n1101), .Y(n564) );
  AND2X1 U3600 ( .A(n981), .B(n968), .Y(n503) );
  AND2X1 U3601 ( .A(n967), .B(n955), .Y(n498) );
  AND2X1 U3602 ( .A(n940), .B(n929), .Y(n482) );
  AND2X1 U3603 ( .A(n917), .B(n906), .Y(n462) );
  AND2X1 U3604 ( .A(n4594), .B(n4807), .Y(n282) );
  AND2X1 U3605 ( .A(n4598), .B(n4806), .Y(n280) );
  AND2X1 U3606 ( .A(n4661), .B(n678), .Y(n279) );
  AND2X1 U3607 ( .A(n4595), .B(n4805), .Y(n278) );
  AND2X1 U3608 ( .A(n4539), .B(n4808), .Y(n277) );
  BUFX2 U3609 ( .A(n4781), .Y(n3913) );
  BUFX2 U3610 ( .A(n4777), .Y(n3914) );
  AND2X2 U3611 ( .A(n524), .B(n550), .Y(n3938) );
  INVX2 U3612 ( .A(n469), .Y(n4689) );
  BUFX2 U3613 ( .A(n4852), .Y(n3915) );
  INVX2 U3614 ( .A(n4921), .Y(n4763) );
  INVX1 U3615 ( .A(n576), .Y(n575) );
  OR2X1 U3616 ( .A(n4412), .B(n3942), .Y(n2325) );
  AND2X1 U3617 ( .A(n4422), .B(n3962), .Y(n2285) );
  OR2X1 U3618 ( .A(b[25]), .B(b[26]), .Y(n2302) );
  OR2X1 U3619 ( .A(n4393), .B(n4747), .Y(n2383) );
  AND2X1 U3620 ( .A(n3941), .B(n3963), .Y(n2426) );
  OR2X1 U3621 ( .A(n4620), .B(n4749), .Y(n2444) );
  XOR2X1 U3622 ( .A(n2441), .B(n4459), .Y(n3916) );
  XOR2X1 U3623 ( .A(n2411), .B(n4377), .Y(n3917) );
  XOR2X1 U3624 ( .A(n2425), .B(n4375), .Y(n3918) );
  XOR2X1 U3625 ( .A(n2478), .B(n4461), .Y(n3919) );
  XOR2X1 U3626 ( .A(n2459), .B(n4374), .Y(n3920) );
  XOR2X1 U3627 ( .A(n2448), .B(n4496), .Y(n3921) );
  XOR2X1 U3628 ( .A(n2472), .B(n4473), .Y(n3922) );
  XOR2X1 U3629 ( .A(n2396), .B(n4378), .Y(n3923) );
  XOR2X1 U3630 ( .A(a[1]), .B(a[0]), .Y(n3924) );
  INVX1 U3631 ( .A(b[11]), .Y(n5002) );
  INVX1 U3632 ( .A(b[21]), .Y(n5018) );
  INVX1 U3633 ( .A(b[9]), .Y(n4998) );
  INVX1 U3634 ( .A(b[18]), .Y(n5014) );
  AND2X1 U3635 ( .A(b[26]), .B(b[25]), .Y(n2303) );
  OR2X1 U3636 ( .A(n4755), .B(n4627), .Y(n2309) );
  OR2X1 U3637 ( .A(n4411), .B(n4442), .Y(n2241) );
  INVX1 U3638 ( .A(n518), .Y(n3937) );
  OR2X1 U3639 ( .A(n4742), .B(n4870), .Y(n568) );
  AND2X1 U3640 ( .A(n4423), .B(n4406), .Y(n2365) );
  AND2X1 U3641 ( .A(n4909), .B(n778), .Y(n493) );
  OR2X1 U3642 ( .A(n4689), .B(n4413), .Y(n366) );
  OR2X1 U3643 ( .A(n4507), .B(n4736), .Y(n370) );
  OR2X1 U3644 ( .A(n4480), .B(n4626), .Y(n2265) );
  OR2X1 U3645 ( .A(b[11]), .B(b[10]), .Y(n2434) );
  INVX1 U3646 ( .A(n2446), .Y(n4749) );
  OR2X1 U3647 ( .A(b[9]), .B(b[8]), .Y(n2446) );
  AND2X1 U3648 ( .A(n4557), .B(n4688), .Y(n306) );
  OR2X1 U3649 ( .A(b[23]), .B(b[24]), .Y(n2320) );
  INVX1 U3650 ( .A(n558), .Y(n4743) );
  OR2X1 U3651 ( .A(n4743), .B(n4872), .Y(n556) );
  OR2X1 U3652 ( .A(n4420), .B(n4689), .Y(n304) );
  AND2X1 U3653 ( .A(n4516), .B(n4482), .Y(n469) );
  AND2X1 U3654 ( .A(n4907), .B(n4908), .Y(n594) );
  XOR2X1 U3655 ( .A(n583), .B(n263), .Y(product[32]) );
  OR2X2 U3656 ( .A(n2325), .B(n3944), .Y(n2250) );
  XOR2X1 U3657 ( .A(n3926), .B(n247), .Y(product[48]) );
  INVX1 U3658 ( .A(n463), .Y(n3926) );
  INVX1 U3659 ( .A(n3933), .Y(n3927) );
  INVX1 U3660 ( .A(n3927), .Y(n3928) );
  INVX1 U3661 ( .A(n4923), .Y(n520) );
  BUFX2 U3662 ( .A(n533), .Y(n3929) );
  AND2X2 U3663 ( .A(n4409), .B(n4628), .Y(n317) );
  INVX1 U3664 ( .A(n468), .Y(n3930) );
  INVX1 U3665 ( .A(n3930), .Y(n3931) );
  XNOR2X1 U3666 ( .A(n3936), .B(n4390), .Y(product[42]) );
  AND2X2 U3667 ( .A(n4762), .B(n547), .Y(n3932) );
  INVX2 U3668 ( .A(n576), .Y(n3933) );
  OAI21X1 U3669 ( .A(n3933), .B(n4358), .C(n4320), .Y(n3934) );
  XOR2X1 U3670 ( .A(n520), .B(n254), .Y(product[41]) );
  BUFX2 U3671 ( .A(n547), .Y(n3935) );
  OAI21X1 U3672 ( .A(n4923), .B(n3937), .C(n4678), .Y(n3936) );
  AND2X2 U3673 ( .A(n4556), .B(n4688), .Y(n346) );
  BUFX2 U3674 ( .A(n643), .Y(n3939) );
  AND2X2 U3675 ( .A(n4764), .B(n552), .Y(n536) );
  INVX1 U3676 ( .A(n4921), .Y(n3940) );
  INVX2 U3677 ( .A(n4921), .Y(n4923) );
  INVX1 U3678 ( .A(n4921), .Y(n4922) );
  OR2X2 U3679 ( .A(n1377), .B(n1388), .Y(n4808) );
  INVX1 U3680 ( .A(n2444), .Y(n3941) );
  INVX1 U3681 ( .A(n2365), .Y(n3942) );
  OR2X2 U3682 ( .A(n2325), .B(n4415), .Y(n2274) );
  INVX1 U3683 ( .A(n2274), .Y(n3943) );
  INVX1 U3684 ( .A(n2252), .Y(n3944) );
  INVX1 U3685 ( .A(n676), .Y(n3945) );
  AND2X2 U3686 ( .A(n3932), .B(n3925), .Y(n524) );
  INVX1 U3687 ( .A(n357), .Y(n3946) );
  BUFX2 U3688 ( .A(n2240), .Y(n3947) );
  BUFX2 U3689 ( .A(n296), .Y(n3948) );
  INVX1 U3690 ( .A(n2398), .Y(n3949) );
  OR2X2 U3691 ( .A(n2325), .B(n4416), .Y(n2261) );
  INVX1 U3692 ( .A(n2261), .Y(n3950) );
  AND2X2 U3693 ( .A(n4917), .B(n4391), .Y(n383) );
  INVX1 U3694 ( .A(n383), .Y(n3951) );
  INVX1 U3695 ( .A(n335), .Y(n3952) );
  INVX1 U3696 ( .A(n324), .Y(n3953) );
  AND2X2 U3697 ( .A(n4919), .B(n3957), .Y(n295) );
  INVX1 U3698 ( .A(n295), .Y(n3954) );
  INVX1 U3699 ( .A(n2239), .Y(n3955) );
  BUFX2 U3700 ( .A(n2397), .Y(n3956) );
  INVX1 U3701 ( .A(n304), .Y(n3957) );
  AND2X2 U3702 ( .A(n4732), .B(n4658), .Y(n328) );
  INVX1 U3703 ( .A(n328), .Y(n3958) );
  BUFX2 U3704 ( .A(n2273), .Y(n3959) );
  BUFX2 U3705 ( .A(n530), .Y(n3960) );
  INVX4 U3706 ( .A(n231), .Y(n4688) );
  OR2X2 U3707 ( .A(n4689), .B(n4419), .Y(n344) );
  INVX1 U3708 ( .A(n344), .Y(n3961) );
  OR2X2 U3709 ( .A(n4505), .B(n4745), .Y(n2291) );
  INVX1 U3710 ( .A(n2291), .Y(n3962) );
  INVX1 U3711 ( .A(n2432), .Y(n3963) );
  BUFX2 U3712 ( .A(n653), .Y(n3964) );
  AND2X1 U3713 ( .A(n4546), .B(n656), .Y(n275) );
  INVX1 U3714 ( .A(n275), .Y(n3965) );
  BUFX2 U3715 ( .A(n2169), .Y(n3966) );
  BUFX2 U3716 ( .A(n2106), .Y(n3967) );
  BUFX2 U3717 ( .A(n2043), .Y(n3968) );
  INVX1 U3718 ( .A(n1980), .Y(n3969) );
  INVX1 U3719 ( .A(n3969), .Y(n3970) );
  BUFX2 U3720 ( .A(n1917), .Y(n3971) );
  BUFX2 U3721 ( .A(n1854), .Y(n3972) );
  BUFX2 U3722 ( .A(n1791), .Y(n3973) );
  BUFX2 U3723 ( .A(n1728), .Y(n3974) );
  BUFX2 U3724 ( .A(n1665), .Y(n3975) );
  BUFX2 U3725 ( .A(n1602), .Y(n3976) );
  BUFX2 U3726 ( .A(n1539), .Y(n3977) );
  BUFX2 U3727 ( .A(n2454), .Y(n3978) );
  BUFX2 U3728 ( .A(n2413), .Y(n3979) );
  BUFX2 U3729 ( .A(n2401), .Y(n3980) );
  BUFX2 U3730 ( .A(n2332), .Y(n3981) );
  BUFX2 U3731 ( .A(n2299), .Y(n3982) );
  BUFX2 U3732 ( .A(n2277), .Y(n3983) );
  BUFX2 U3733 ( .A(n2264), .Y(n3984) );
  BUFX2 U3734 ( .A(n2253), .Y(n3985) );
  BUFX2 U3735 ( .A(n2244), .Y(n3986) );
  BUFX2 U3736 ( .A(n3591), .Y(n3987) );
  BUFX2 U3737 ( .A(n3590), .Y(n3988) );
  BUFX2 U3738 ( .A(n3589), .Y(n3989) );
  BUFX2 U3739 ( .A(n3588), .Y(n3990) );
  BUFX2 U3740 ( .A(n3587), .Y(n3991) );
  BUFX2 U3741 ( .A(n3586), .Y(n3992) );
  BUFX2 U3742 ( .A(n3585), .Y(n3993) );
  BUFX2 U3743 ( .A(n3584), .Y(n3994) );
  BUFX2 U3744 ( .A(n3583), .Y(n3995) );
  BUFX2 U3745 ( .A(n3582), .Y(n3996) );
  BUFX2 U3746 ( .A(n3581), .Y(n3997) );
  BUFX2 U3747 ( .A(n3580), .Y(n3998) );
  BUFX2 U3748 ( .A(n3579), .Y(n3999) );
  BUFX2 U3749 ( .A(n3578), .Y(n4000) );
  BUFX2 U3750 ( .A(n3577), .Y(n4001) );
  BUFX2 U3751 ( .A(n3576), .Y(n4002) );
  BUFX2 U3752 ( .A(n3575), .Y(n4003) );
  BUFX2 U3753 ( .A(n3574), .Y(n4004) );
  BUFX2 U3754 ( .A(n3573), .Y(n4005) );
  BUFX2 U3755 ( .A(n3572), .Y(n4006) );
  BUFX2 U3756 ( .A(n3571), .Y(n4007) );
  BUFX2 U3757 ( .A(n3570), .Y(n4008) );
  BUFX2 U3758 ( .A(n3569), .Y(n4009) );
  BUFX2 U3759 ( .A(n3568), .Y(n4010) );
  BUFX2 U3760 ( .A(n3567), .Y(n4011) );
  BUFX2 U3761 ( .A(n3566), .Y(n4012) );
  BUFX2 U3762 ( .A(n3565), .Y(n4013) );
  BUFX2 U3763 ( .A(n3564), .Y(n4014) );
  BUFX2 U3764 ( .A(n3563), .Y(n4015) );
  BUFX2 U3765 ( .A(n3562), .Y(n4016) );
  BUFX2 U3766 ( .A(n3524), .Y(n4017) );
  BUFX2 U3767 ( .A(n3523), .Y(n4018) );
  BUFX2 U3768 ( .A(n3522), .Y(n4019) );
  BUFX2 U3769 ( .A(n3521), .Y(n4020) );
  BUFX2 U3770 ( .A(n3520), .Y(n4021) );
  BUFX2 U3771 ( .A(n3519), .Y(n4022) );
  BUFX2 U3772 ( .A(n3518), .Y(n4023) );
  BUFX2 U3773 ( .A(n3517), .Y(n4024) );
  BUFX2 U3774 ( .A(n3516), .Y(n4025) );
  BUFX2 U3775 ( .A(n3515), .Y(n4026) );
  BUFX2 U3776 ( .A(n3514), .Y(n4027) );
  BUFX2 U3777 ( .A(n3513), .Y(n4028) );
  BUFX2 U3778 ( .A(n3512), .Y(n4029) );
  BUFX2 U3779 ( .A(n3511), .Y(n4030) );
  BUFX2 U3780 ( .A(n3510), .Y(n4031) );
  BUFX2 U3781 ( .A(n3509), .Y(n4032) );
  BUFX2 U3782 ( .A(n3508), .Y(n4033) );
  BUFX2 U3783 ( .A(n3507), .Y(n4034) );
  BUFX2 U3784 ( .A(n3506), .Y(n4035) );
  BUFX2 U3785 ( .A(n3505), .Y(n4036) );
  BUFX2 U3786 ( .A(n3504), .Y(n4037) );
  BUFX2 U3787 ( .A(n3503), .Y(n4038) );
  BUFX2 U3788 ( .A(n3502), .Y(n4039) );
  BUFX2 U3789 ( .A(n3501), .Y(n4040) );
  BUFX2 U3790 ( .A(n3500), .Y(n4041) );
  BUFX2 U3791 ( .A(n3499), .Y(n4042) );
  BUFX2 U3792 ( .A(n3498), .Y(n4043) );
  BUFX2 U3793 ( .A(n3497), .Y(n4044) );
  BUFX2 U3794 ( .A(n3496), .Y(n4045) );
  BUFX2 U3795 ( .A(n3495), .Y(n4046) );
  BUFX2 U3796 ( .A(n3457), .Y(n4047) );
  BUFX2 U3797 ( .A(n3456), .Y(n4048) );
  BUFX2 U3798 ( .A(n3455), .Y(n4049) );
  BUFX2 U3799 ( .A(n3454), .Y(n4050) );
  BUFX2 U3800 ( .A(n3453), .Y(n4051) );
  BUFX2 U3801 ( .A(n3452), .Y(n4052) );
  BUFX2 U3802 ( .A(n3451), .Y(n4053) );
  BUFX2 U3803 ( .A(n3450), .Y(n4054) );
  BUFX2 U3804 ( .A(n3449), .Y(n4055) );
  BUFX2 U3805 ( .A(n3448), .Y(n4056) );
  BUFX2 U3806 ( .A(n3447), .Y(n4057) );
  BUFX2 U3807 ( .A(n3446), .Y(n4058) );
  BUFX2 U3808 ( .A(n3445), .Y(n4059) );
  BUFX2 U3809 ( .A(n3444), .Y(n4060) );
  BUFX2 U3810 ( .A(n3443), .Y(n4061) );
  BUFX2 U3811 ( .A(n3442), .Y(n4062) );
  BUFX2 U3812 ( .A(n3441), .Y(n4063) );
  BUFX2 U3813 ( .A(n3440), .Y(n4064) );
  BUFX2 U3814 ( .A(n3439), .Y(n4065) );
  BUFX2 U3815 ( .A(n3438), .Y(n4066) );
  BUFX2 U3816 ( .A(n3437), .Y(n4067) );
  BUFX2 U3817 ( .A(n3436), .Y(n4068) );
  BUFX2 U3818 ( .A(n3435), .Y(n4069) );
  BUFX2 U3819 ( .A(n3434), .Y(n4070) );
  BUFX2 U3820 ( .A(n3433), .Y(n4071) );
  BUFX2 U3821 ( .A(n3432), .Y(n4072) );
  BUFX2 U3822 ( .A(n3431), .Y(n4073) );
  BUFX2 U3823 ( .A(n3430), .Y(n4074) );
  BUFX2 U3824 ( .A(n3429), .Y(n4075) );
  BUFX2 U3825 ( .A(n3428), .Y(n4076) );
  BUFX2 U3826 ( .A(n3390), .Y(n4077) );
  BUFX2 U3827 ( .A(n3389), .Y(n4078) );
  BUFX2 U3828 ( .A(n3388), .Y(n4079) );
  BUFX2 U3829 ( .A(n3387), .Y(n4080) );
  BUFX2 U3830 ( .A(n3386), .Y(n4081) );
  BUFX2 U3831 ( .A(n3385), .Y(n4082) );
  BUFX2 U3832 ( .A(n3384), .Y(n4083) );
  BUFX2 U3833 ( .A(n3383), .Y(n4084) );
  BUFX2 U3834 ( .A(n3382), .Y(n4085) );
  BUFX2 U3835 ( .A(n3381), .Y(n4086) );
  BUFX2 U3836 ( .A(n3380), .Y(n4087) );
  BUFX2 U3837 ( .A(n3379), .Y(n4088) );
  BUFX2 U3838 ( .A(n3378), .Y(n4089) );
  BUFX2 U3839 ( .A(n3377), .Y(n4090) );
  BUFX2 U3840 ( .A(n3376), .Y(n4091) );
  BUFX2 U3841 ( .A(n3375), .Y(n4092) );
  BUFX2 U3842 ( .A(n3374), .Y(n4093) );
  BUFX2 U3843 ( .A(n3373), .Y(n4094) );
  BUFX2 U3844 ( .A(n3372), .Y(n4095) );
  BUFX2 U3845 ( .A(n3371), .Y(n4096) );
  BUFX2 U3846 ( .A(n3370), .Y(n4097) );
  BUFX2 U3847 ( .A(n3369), .Y(n4098) );
  BUFX2 U3848 ( .A(n3368), .Y(n4099) );
  BUFX2 U3849 ( .A(n3367), .Y(n4100) );
  BUFX2 U3850 ( .A(n3366), .Y(n4101) );
  BUFX2 U3851 ( .A(n3365), .Y(n4102) );
  BUFX2 U3852 ( .A(n3364), .Y(n4103) );
  BUFX2 U3853 ( .A(n3363), .Y(n4104) );
  BUFX2 U3854 ( .A(n3362), .Y(n4105) );
  BUFX2 U3855 ( .A(n3361), .Y(n4106) );
  BUFX2 U3856 ( .A(n3323), .Y(n4107) );
  BUFX2 U3857 ( .A(n3322), .Y(n4108) );
  BUFX2 U3858 ( .A(n3321), .Y(n4109) );
  BUFX2 U3859 ( .A(n3320), .Y(n4110) );
  BUFX2 U3860 ( .A(n3319), .Y(n4111) );
  BUFX2 U3861 ( .A(n3318), .Y(n4112) );
  BUFX2 U3862 ( .A(n3317), .Y(n4113) );
  BUFX2 U3863 ( .A(n3316), .Y(n4114) );
  BUFX2 U3864 ( .A(n3315), .Y(n4115) );
  BUFX2 U3865 ( .A(n3314), .Y(n4116) );
  BUFX2 U3866 ( .A(n3313), .Y(n4117) );
  BUFX2 U3867 ( .A(n3312), .Y(n4118) );
  BUFX2 U3868 ( .A(n3311), .Y(n4119) );
  BUFX2 U3869 ( .A(n3310), .Y(n4120) );
  BUFX2 U3870 ( .A(n3309), .Y(n4121) );
  BUFX2 U3871 ( .A(n3308), .Y(n4122) );
  BUFX2 U3872 ( .A(n3307), .Y(n4123) );
  BUFX2 U3873 ( .A(n3306), .Y(n4124) );
  BUFX2 U3874 ( .A(n3305), .Y(n4125) );
  BUFX2 U3875 ( .A(n3304), .Y(n4126) );
  BUFX2 U3876 ( .A(n3303), .Y(n4127) );
  BUFX2 U3877 ( .A(n3302), .Y(n4128) );
  BUFX2 U3878 ( .A(n3301), .Y(n4129) );
  BUFX2 U3879 ( .A(n3300), .Y(n4130) );
  BUFX2 U3880 ( .A(n3299), .Y(n4131) );
  BUFX2 U3881 ( .A(n3298), .Y(n4132) );
  BUFX2 U3882 ( .A(n3297), .Y(n4133) );
  BUFX2 U3883 ( .A(n3296), .Y(n4134) );
  BUFX2 U3884 ( .A(n3295), .Y(n4135) );
  BUFX2 U3885 ( .A(n3294), .Y(n4136) );
  BUFX2 U3886 ( .A(n3256), .Y(n4137) );
  BUFX2 U3887 ( .A(n3255), .Y(n4138) );
  BUFX2 U3888 ( .A(n3254), .Y(n4139) );
  BUFX2 U3889 ( .A(n3253), .Y(n4140) );
  BUFX2 U3890 ( .A(n3252), .Y(n4141) );
  BUFX2 U3891 ( .A(n3251), .Y(n4142) );
  BUFX2 U3892 ( .A(n3250), .Y(n4143) );
  BUFX2 U3893 ( .A(n3249), .Y(n4144) );
  BUFX2 U3894 ( .A(n3248), .Y(n4145) );
  BUFX2 U3895 ( .A(n3247), .Y(n4146) );
  BUFX2 U3896 ( .A(n3246), .Y(n4147) );
  BUFX2 U3897 ( .A(n3245), .Y(n4148) );
  BUFX2 U3898 ( .A(n3244), .Y(n4149) );
  BUFX2 U3899 ( .A(n3243), .Y(n4150) );
  BUFX2 U3900 ( .A(n3242), .Y(n4151) );
  BUFX2 U3901 ( .A(n3241), .Y(n4152) );
  BUFX2 U3902 ( .A(n3240), .Y(n4153) );
  BUFX2 U3903 ( .A(n3239), .Y(n4154) );
  BUFX2 U3904 ( .A(n3238), .Y(n4155) );
  BUFX2 U3905 ( .A(n3237), .Y(n4156) );
  BUFX2 U3906 ( .A(n3236), .Y(n4157) );
  BUFX2 U3907 ( .A(n3235), .Y(n4158) );
  BUFX2 U3908 ( .A(n3234), .Y(n4159) );
  BUFX2 U3909 ( .A(n3233), .Y(n4160) );
  BUFX2 U3910 ( .A(n3232), .Y(n4161) );
  BUFX2 U3911 ( .A(n3231), .Y(n4162) );
  BUFX2 U3912 ( .A(n3230), .Y(n4163) );
  BUFX2 U3913 ( .A(n3229), .Y(n4164) );
  BUFX2 U3914 ( .A(n3228), .Y(n4165) );
  BUFX2 U3915 ( .A(n3227), .Y(n4166) );
  BUFX2 U3916 ( .A(n3189), .Y(n4167) );
  BUFX2 U3917 ( .A(n3188), .Y(n4168) );
  BUFX2 U3918 ( .A(n3187), .Y(n4169) );
  BUFX2 U3919 ( .A(n3186), .Y(n4170) );
  BUFX2 U3920 ( .A(n3185), .Y(n4171) );
  BUFX2 U3921 ( .A(n3184), .Y(n4172) );
  BUFX2 U3922 ( .A(n3183), .Y(n4173) );
  BUFX2 U3923 ( .A(n3182), .Y(n4174) );
  BUFX2 U3924 ( .A(n3181), .Y(n4175) );
  BUFX2 U3925 ( .A(n3180), .Y(n4176) );
  BUFX2 U3926 ( .A(n3179), .Y(n4177) );
  BUFX2 U3927 ( .A(n3178), .Y(n4178) );
  BUFX2 U3928 ( .A(n3177), .Y(n4179) );
  BUFX2 U3929 ( .A(n3176), .Y(n4180) );
  BUFX2 U3930 ( .A(n3175), .Y(n4181) );
  BUFX2 U3931 ( .A(n3174), .Y(n4182) );
  BUFX2 U3932 ( .A(n3173), .Y(n4183) );
  BUFX2 U3933 ( .A(n3172), .Y(n4184) );
  BUFX2 U3934 ( .A(n3171), .Y(n4185) );
  BUFX2 U3935 ( .A(n3170), .Y(n4186) );
  BUFX2 U3936 ( .A(n3169), .Y(n4187) );
  BUFX2 U3937 ( .A(n3168), .Y(n4188) );
  BUFX2 U3938 ( .A(n3167), .Y(n4189) );
  BUFX2 U3939 ( .A(n3166), .Y(n4190) );
  BUFX2 U3940 ( .A(n3165), .Y(n4191) );
  BUFX2 U3941 ( .A(n3164), .Y(n4192) );
  BUFX2 U3942 ( .A(n3163), .Y(n4193) );
  BUFX2 U3943 ( .A(n3162), .Y(n4194) );
  BUFX2 U3944 ( .A(n3161), .Y(n4195) );
  BUFX2 U3945 ( .A(n3160), .Y(n4196) );
  BUFX2 U3946 ( .A(n3122), .Y(n4197) );
  BUFX2 U3947 ( .A(n3121), .Y(n4198) );
  BUFX2 U3948 ( .A(n3120), .Y(n4199) );
  BUFX2 U3949 ( .A(n3119), .Y(n4200) );
  BUFX2 U3950 ( .A(n3118), .Y(n4201) );
  BUFX2 U3951 ( .A(n3117), .Y(n4202) );
  BUFX2 U3952 ( .A(n3116), .Y(n4203) );
  BUFX2 U3953 ( .A(n3115), .Y(n4204) );
  BUFX2 U3954 ( .A(n3114), .Y(n4205) );
  BUFX2 U3955 ( .A(n3113), .Y(n4206) );
  BUFX2 U3956 ( .A(n3112), .Y(n4207) );
  BUFX2 U3957 ( .A(n3111), .Y(n4208) );
  BUFX2 U3958 ( .A(n3110), .Y(n4209) );
  BUFX2 U3959 ( .A(n3109), .Y(n4210) );
  BUFX2 U3960 ( .A(n3108), .Y(n4211) );
  BUFX2 U3961 ( .A(n3107), .Y(n4212) );
  BUFX2 U3962 ( .A(n3106), .Y(n4213) );
  BUFX2 U3963 ( .A(n3105), .Y(n4214) );
  BUFX2 U3964 ( .A(n3104), .Y(n4215) );
  BUFX2 U3965 ( .A(n3103), .Y(n4216) );
  BUFX2 U3966 ( .A(n3102), .Y(n4217) );
  BUFX2 U3967 ( .A(n3101), .Y(n4218) );
  BUFX2 U3968 ( .A(n3100), .Y(n4219) );
  BUFX2 U3969 ( .A(n3099), .Y(n4220) );
  BUFX2 U3970 ( .A(n3098), .Y(n4221) );
  BUFX2 U3971 ( .A(n3097), .Y(n4222) );
  BUFX2 U3972 ( .A(n3096), .Y(n4223) );
  BUFX2 U3973 ( .A(n3095), .Y(n4224) );
  BUFX2 U3974 ( .A(n3094), .Y(n4225) );
  BUFX2 U3975 ( .A(n3093), .Y(n4226) );
  BUFX2 U3976 ( .A(n3055), .Y(n4227) );
  BUFX2 U3977 ( .A(n3054), .Y(n4228) );
  BUFX2 U3978 ( .A(n3053), .Y(n4229) );
  BUFX2 U3979 ( .A(n3052), .Y(n4230) );
  BUFX2 U3980 ( .A(n3051), .Y(n4231) );
  BUFX2 U3981 ( .A(n3050), .Y(n4232) );
  BUFX2 U3982 ( .A(n3049), .Y(n4233) );
  BUFX2 U3983 ( .A(n3048), .Y(n4234) );
  BUFX2 U3984 ( .A(n3047), .Y(n4235) );
  BUFX2 U3985 ( .A(n3046), .Y(n4236) );
  BUFX2 U3986 ( .A(n3045), .Y(n4237) );
  BUFX2 U3987 ( .A(n3044), .Y(n4238) );
  BUFX2 U3988 ( .A(n3043), .Y(n4239) );
  BUFX2 U3989 ( .A(n3042), .Y(n4240) );
  BUFX2 U3990 ( .A(n3041), .Y(n4241) );
  BUFX2 U3991 ( .A(n3040), .Y(n4242) );
  BUFX2 U3992 ( .A(n3039), .Y(n4243) );
  BUFX2 U3993 ( .A(n3038), .Y(n4244) );
  BUFX2 U3994 ( .A(n3037), .Y(n4245) );
  BUFX2 U3995 ( .A(n3036), .Y(n4246) );
  BUFX2 U3996 ( .A(n3035), .Y(n4247) );
  BUFX2 U3997 ( .A(n3034), .Y(n4248) );
  BUFX2 U3998 ( .A(n3033), .Y(n4249) );
  BUFX2 U3999 ( .A(n3032), .Y(n4250) );
  BUFX2 U4000 ( .A(n3031), .Y(n4251) );
  BUFX2 U4001 ( .A(n3030), .Y(n4252) );
  BUFX2 U4002 ( .A(n3029), .Y(n4253) );
  BUFX2 U4003 ( .A(n3028), .Y(n4254) );
  BUFX2 U4004 ( .A(n3027), .Y(n4255) );
  BUFX2 U4005 ( .A(n3026), .Y(n4256) );
  BUFX2 U4006 ( .A(n3025), .Y(n4257) );
  BUFX2 U4007 ( .A(n2988), .Y(n4258) );
  BUFX2 U4008 ( .A(n2987), .Y(n4259) );
  BUFX2 U4009 ( .A(n2986), .Y(n4260) );
  BUFX2 U4010 ( .A(n2985), .Y(n4261) );
  BUFX2 U4011 ( .A(n2984), .Y(n4262) );
  BUFX2 U4012 ( .A(n2983), .Y(n4263) );
  BUFX2 U4013 ( .A(n2982), .Y(n4264) );
  BUFX2 U4014 ( .A(n2981), .Y(n4265) );
  BUFX2 U4015 ( .A(n2980), .Y(n4266) );
  BUFX2 U4016 ( .A(n2979), .Y(n4267) );
  BUFX2 U4017 ( .A(n2978), .Y(n4268) );
  BUFX2 U4018 ( .A(n2977), .Y(n4269) );
  BUFX2 U4019 ( .A(n2976), .Y(n4270) );
  BUFX2 U4020 ( .A(n2975), .Y(n4271) );
  BUFX2 U4021 ( .A(n2974), .Y(n4272) );
  BUFX2 U4022 ( .A(n2973), .Y(n4273) );
  BUFX2 U4023 ( .A(n2972), .Y(n4274) );
  BUFX2 U4024 ( .A(n2971), .Y(n4275) );
  BUFX2 U4025 ( .A(n2970), .Y(n4276) );
  BUFX2 U4026 ( .A(n2969), .Y(n4277) );
  BUFX2 U4027 ( .A(n2968), .Y(n4278) );
  BUFX2 U4028 ( .A(n2967), .Y(n4279) );
  BUFX2 U4029 ( .A(n2966), .Y(n4280) );
  BUFX2 U4030 ( .A(n2965), .Y(n4281) );
  BUFX2 U4031 ( .A(n2964), .Y(n4282) );
  BUFX2 U4032 ( .A(n2963), .Y(n4283) );
  BUFX2 U4033 ( .A(n2962), .Y(n4284) );
  BUFX2 U4034 ( .A(n2961), .Y(n4285) );
  BUFX2 U4035 ( .A(n2960), .Y(n4286) );
  BUFX2 U4036 ( .A(n2959), .Y(n4287) );
  BUFX2 U4037 ( .A(n2921), .Y(n4288) );
  BUFX2 U4038 ( .A(n2920), .Y(n4289) );
  BUFX2 U4039 ( .A(n2919), .Y(n4290) );
  BUFX2 U4040 ( .A(n2918), .Y(n4291) );
  BUFX2 U4041 ( .A(n2917), .Y(n4292) );
  BUFX2 U4042 ( .A(n2916), .Y(n4293) );
  BUFX2 U4043 ( .A(n2915), .Y(n4294) );
  BUFX2 U4044 ( .A(n2914), .Y(n4295) );
  BUFX2 U4045 ( .A(n2913), .Y(n4296) );
  BUFX2 U4046 ( .A(n2912), .Y(n4297) );
  BUFX2 U4047 ( .A(n2911), .Y(n4298) );
  BUFX2 U4048 ( .A(n2910), .Y(n4299) );
  BUFX2 U4049 ( .A(n2909), .Y(n4300) );
  BUFX2 U4050 ( .A(n2908), .Y(n4301) );
  BUFX2 U4051 ( .A(n2907), .Y(n4302) );
  BUFX2 U4052 ( .A(n2906), .Y(n4303) );
  BUFX2 U4053 ( .A(n2905), .Y(n4304) );
  BUFX2 U4054 ( .A(n2904), .Y(n4305) );
  BUFX2 U4055 ( .A(n2903), .Y(n4306) );
  BUFX2 U4056 ( .A(n2902), .Y(n4307) );
  BUFX2 U4057 ( .A(n2901), .Y(n4308) );
  BUFX2 U4058 ( .A(n2900), .Y(n4309) );
  BUFX2 U4059 ( .A(n2899), .Y(n4310) );
  BUFX2 U4060 ( .A(n2898), .Y(n4311) );
  BUFX2 U4061 ( .A(n2897), .Y(n4312) );
  BUFX2 U4062 ( .A(n2896), .Y(n4313) );
  BUFX2 U4063 ( .A(n2895), .Y(n4314) );
  BUFX2 U4064 ( .A(n2894), .Y(n4315) );
  BUFX2 U4065 ( .A(n2893), .Y(n4316) );
  BUFX2 U4066 ( .A(n2892), .Y(n4317) );
  BUFX2 U4067 ( .A(n697), .Y(n4318) );
  BUFX2 U4068 ( .A(n664), .Y(n4319) );
  BUFX2 U4069 ( .A(n537), .Y(n4320) );
  INVX1 U4070 ( .A(n525), .Y(n4321) );
  INVX1 U4071 ( .A(n4321), .Y(n4322) );
  BUFX2 U4072 ( .A(n452), .Y(n4323) );
  BUFX2 U4073 ( .A(n443), .Y(n4324) );
  BUFX2 U4074 ( .A(n432), .Y(n4325) );
  BUFX2 U4075 ( .A(n425), .Y(n4326) );
  BUFX2 U4076 ( .A(n408), .Y(n4327) );
  BUFX2 U4077 ( .A(n397), .Y(n4328) );
  INVX1 U4078 ( .A(n384), .Y(n4329) );
  INVX1 U4079 ( .A(n4329), .Y(n4330) );
  BUFX2 U4080 ( .A(n377), .Y(n4331) );
  BUFX2 U4081 ( .A(n369), .Y(n4332) );
  INVX1 U4082 ( .A(n358), .Y(n4333) );
  INVX1 U4083 ( .A(n4333), .Y(n4334) );
  BUFX2 U4084 ( .A(n347), .Y(n4335) );
  INVX1 U4085 ( .A(n336), .Y(n4336) );
  INVX1 U4086 ( .A(n4336), .Y(n4337) );
  INVX1 U4087 ( .A(n325), .Y(n4338) );
  INVX1 U4088 ( .A(n4338), .Y(n4339) );
  BUFX2 U4089 ( .A(n314), .Y(n4340) );
  BUFX2 U4090 ( .A(n307), .Y(n4341) );
  OR2X1 U4091 ( .A(n3924), .B(n2202), .Y(n2201) );
  INVX1 U4092 ( .A(n2201), .Y(n4342) );
  OR2X1 U4093 ( .A(n2383), .B(n4440), .Y(n2376) );
  INVX1 U4094 ( .A(n2376), .Y(n4343) );
  OR2X1 U4095 ( .A(n3942), .B(n4754), .Y(n2356) );
  INVX1 U4096 ( .A(n2356), .Y(n4344) );
  OR2X1 U4097 ( .A(n4392), .B(n4441), .Y(n2338) );
  INVX1 U4098 ( .A(n2338), .Y(n4345) );
  OR2X1 U4099 ( .A(n2325), .B(n4755), .Y(n2318) );
  INVX1 U4100 ( .A(n2318), .Y(n4346) );
  OR2X1 U4101 ( .A(n2325), .B(n2309), .Y(n2305) );
  INVX1 U4102 ( .A(n2305), .Y(n4347) );
  OR2X1 U4103 ( .A(n2325), .B(n4414), .Y(n2296) );
  INVX1 U4104 ( .A(n2296), .Y(n4348) );
  INVX1 U4105 ( .A(n2283), .Y(n4349) );
  INVX1 U4106 ( .A(n2250), .Y(n4350) );
  OR2X1 U4107 ( .A(n4623), .B(n4680), .Y(n654) );
  INVX1 U4108 ( .A(n654), .Y(n4351) );
  AND2X1 U4109 ( .A(n4408), .B(n4405), .Y(n2453) );
  INVX1 U4110 ( .A(n2453), .Y(n4352) );
  INVX1 U4111 ( .A(n2412), .Y(n4353) );
  AND2X1 U4112 ( .A(n4816), .B(n4807), .Y(n696) );
  INVX1 U4113 ( .A(n696), .Y(n4354) );
  INVX1 U4114 ( .A(n663), .Y(n4355) );
  AND2X1 U4115 ( .A(n771), .B(n4464), .Y(n431) );
  INVX1 U4116 ( .A(n431), .Y(n4356) );
  AND2X1 U4117 ( .A(n317), .B(n4618), .Y(n313) );
  INVX1 U4118 ( .A(n313), .Y(n4357) );
  INVX1 U4119 ( .A(n536), .Y(n4358) );
  AND2X1 U4120 ( .A(n4757), .B(n4770), .Y(n3625) );
  INVX1 U4121 ( .A(n3625), .Y(n4359) );
  BUFX2 U4122 ( .A(n2420), .Y(n4360) );
  INVX1 U4123 ( .A(n2382), .Y(n4361) );
  INVX1 U4124 ( .A(n4361), .Y(n4362) );
  INVX1 U4125 ( .A(n2375), .Y(n4363) );
  INVX1 U4126 ( .A(n4363), .Y(n4364) );
  INVX1 U4127 ( .A(n2362), .Y(n4365) );
  INVX1 U4128 ( .A(n4365), .Y(n4366) );
  BUFX2 U4129 ( .A(n2355), .Y(n4367) );
  INVX1 U4130 ( .A(n2344), .Y(n4368) );
  INVX1 U4131 ( .A(n4368), .Y(n4369) );
  BUFX2 U4132 ( .A(n2337), .Y(n4370) );
  BUFX2 U4133 ( .A(n2324), .Y(n4371) );
  BUFX2 U4134 ( .A(n2282), .Y(n4372) );
  AND2X1 U4135 ( .A(n4433), .B(n2460), .Y(n2229) );
  INVX1 U4136 ( .A(n2229), .Y(n4373) );
  AND2X1 U4137 ( .A(n4395), .B(n2457), .Y(n2228) );
  INVX1 U4138 ( .A(n2228), .Y(n4374) );
  AND2X1 U4139 ( .A(n4672), .B(n2423), .Y(n2223) );
  INVX1 U4140 ( .A(n2223), .Y(n4375) );
  AND2X1 U4141 ( .A(n4601), .B(n2418), .Y(n2222) );
  INVX1 U4142 ( .A(n2222), .Y(n4376) );
  AND2X1 U4143 ( .A(n4675), .B(n2409), .Y(n2221) );
  INVX1 U4144 ( .A(n2221), .Y(n4377) );
  AND2X1 U4145 ( .A(n4673), .B(n2394), .Y(n2219) );
  INVX1 U4146 ( .A(n2219), .Y(n4378) );
  AND2X1 U4147 ( .A(n4434), .B(n2378), .Y(n2217) );
  INVX1 U4148 ( .A(n2217), .Y(n4379) );
  AND2X1 U4149 ( .A(n4396), .B(n2373), .Y(n2216) );
  INVX1 U4150 ( .A(n2216), .Y(n4380) );
  AND2X1 U4151 ( .A(n4435), .B(n2358), .Y(n2215) );
  INVX1 U4152 ( .A(n2215), .Y(n4381) );
  AND2X1 U4153 ( .A(n4397), .B(n2353), .Y(n2214) );
  INVX1 U4154 ( .A(n2214), .Y(n4382) );
  AND2X1 U4155 ( .A(n4436), .B(n2340), .Y(n2213) );
  INVX1 U4156 ( .A(n2213), .Y(n4383) );
  AND2X1 U4157 ( .A(n4398), .B(n2335), .Y(n2212) );
  INVX1 U4158 ( .A(n2212), .Y(n4384) );
  AND2X1 U4159 ( .A(n4682), .B(n2320), .Y(n2211) );
  INVX1 U4160 ( .A(n2211), .Y(n4385) );
  AND2X1 U4161 ( .A(n4561), .B(n2280), .Y(n2207) );
  INVX1 U4162 ( .A(n2207), .Y(n4386) );
  AND2X1 U4163 ( .A(n4510), .B(n2271), .Y(n2206) );
  INVX1 U4164 ( .A(n2206), .Y(n4387) );
  AND2X1 U4165 ( .A(n4677), .B(n3929), .Y(n256) );
  INVX1 U4166 ( .A(n256), .Y(n4388) );
  AND2X1 U4167 ( .A(n4607), .B(n528), .Y(n255) );
  INVX1 U4168 ( .A(n255), .Y(n4389) );
  AND2X1 U4169 ( .A(n4550), .B(n513), .Y(n253) );
  INVX1 U4170 ( .A(n253), .Y(n4390) );
  OR2X1 U4171 ( .A(n4689), .B(n4418), .Y(n394) );
  INVX1 U4172 ( .A(n394), .Y(n4391) );
  AND2X1 U4173 ( .A(n4437), .B(n2365), .Y(n2347) );
  INVX1 U4174 ( .A(n2347), .Y(n4392) );
  OR2X1 U4175 ( .A(b[15]), .B(b[16]), .Y(n2394) );
  INVX1 U4176 ( .A(n2394), .Y(n4393) );
  INVX1 U4177 ( .A(n317), .Y(n4394) );
  AND2X1 U4178 ( .A(b[6]), .B(b[7]), .Y(n2458) );
  INVX1 U4179 ( .A(n2458), .Y(n4395) );
  AND2X1 U4180 ( .A(b[18]), .B(b[19]), .Y(n2374) );
  INVX1 U4181 ( .A(n2374), .Y(n4396) );
  AND2X1 U4182 ( .A(b[20]), .B(b[21]), .Y(n2354) );
  INVX1 U4183 ( .A(n2354), .Y(n4397) );
  AND2X1 U4184 ( .A(b[22]), .B(b[23]), .Y(n2336) );
  INVX1 U4185 ( .A(n2336), .Y(n4398) );
  INVX1 U4186 ( .A(n4400), .Y(n4399) );
  BUFX2 U4187 ( .A(n2348), .Y(n4400) );
  INVX1 U4188 ( .A(n675), .Y(n4401) );
  INVX1 U4189 ( .A(n4401), .Y(n4402) );
  OR2X2 U4190 ( .A(n4741), .B(n4542), .Y(n2402) );
  INVX1 U4191 ( .A(n2402), .Y(n4403) );
  OR2X1 U4192 ( .A(n4429), .B(n4441), .Y(n2333) );
  INVX1 U4193 ( .A(n2333), .Y(n4404) );
  OR2X1 U4194 ( .A(n4504), .B(n4746), .Y(n2463) );
  INVX1 U4195 ( .A(n2463), .Y(n4405) );
  OR2X1 U4196 ( .A(n4440), .B(n4432), .Y(n2371) );
  INVX1 U4197 ( .A(n2371), .Y(n4406) );
  INVX1 U4198 ( .A(n2241), .Y(n4407) );
  OR2X1 U4199 ( .A(n4679), .B(n4744), .Y(n2455) );
  INVX1 U4200 ( .A(n2455), .Y(n4408) );
  INVX1 U4201 ( .A(n319), .Y(n4409) );
  OR2X2 U4202 ( .A(n3958), .B(n4898), .Y(n319) );
  INVX1 U4203 ( .A(n2400), .Y(n4410) );
  AND2X1 U4204 ( .A(n4687), .B(n4515), .Y(n2243) );
  INVX1 U4205 ( .A(n2243), .Y(n4411) );
  AND2X2 U4206 ( .A(n4437), .B(n4404), .Y(n2331) );
  INVX1 U4207 ( .A(n2331), .Y(n4412) );
  INVX1 U4208 ( .A(n368), .Y(n4413) );
  AND2X1 U4209 ( .A(n2302), .B(n4422), .Y(n2298) );
  INVX1 U4210 ( .A(n2298), .Y(n4414) );
  INVX1 U4211 ( .A(n2276), .Y(n4415) );
  INVX1 U4212 ( .A(n2263), .Y(n4416) );
  INVX1 U4213 ( .A(n524), .Y(n4417) );
  INVX1 U4214 ( .A(n396), .Y(n4418) );
  INVX1 U4215 ( .A(n346), .Y(n4419) );
  INVX1 U4216 ( .A(n306), .Y(n4420) );
  BUFX2 U4217 ( .A(n2462), .Y(n4421) );
  INVX1 U4218 ( .A(n2309), .Y(n4422) );
  INVX1 U4219 ( .A(n2383), .Y(n4423) );
  INVX1 U4220 ( .A(n2325), .Y(n4424) );
  INVX1 U4221 ( .A(n2427), .Y(n4425) );
  INVX1 U4222 ( .A(n4425), .Y(n4426) );
  INVX1 U4223 ( .A(n2286), .Y(n4427) );
  INVX1 U4224 ( .A(n4427), .Y(n4428) );
  INVX1 U4225 ( .A(n2335), .Y(n4429) );
  OR2X1 U4226 ( .A(b[23]), .B(b[22]), .Y(n2335) );
  INVX1 U4227 ( .A(n2426), .Y(n4430) );
  INVX1 U4228 ( .A(n2353), .Y(n4431) );
  OR2X1 U4229 ( .A(b[21]), .B(b[20]), .Y(n2353) );
  INVX1 U4230 ( .A(n2373), .Y(n4432) );
  OR2X1 U4231 ( .A(b[19]), .B(b[18]), .Y(n2373) );
  AND2X1 U4232 ( .A(b[6]), .B(b[5]), .Y(n2461) );
  INVX1 U4233 ( .A(n2461), .Y(n4433) );
  AND2X1 U4234 ( .A(b[18]), .B(b[17]), .Y(n2381) );
  INVX1 U4235 ( .A(n2381), .Y(n4434) );
  AND2X1 U4236 ( .A(b[20]), .B(b[19]), .Y(n2361) );
  INVX1 U4237 ( .A(n2361), .Y(n4435) );
  AND2X1 U4238 ( .A(b[21]), .B(b[22]), .Y(n2343) );
  INVX1 U4239 ( .A(n2343), .Y(n4436) );
  INVX1 U4240 ( .A(n2349), .Y(n4437) );
  INVX1 U4241 ( .A(n2366), .Y(n4438) );
  INVX1 U4242 ( .A(n4438), .Y(n4439) );
  INVX1 U4243 ( .A(n2378), .Y(n4440) );
  OR2X1 U4244 ( .A(b[17]), .B(b[18]), .Y(n2378) );
  INVX1 U4245 ( .A(n2340), .Y(n4441) );
  OR2X1 U4246 ( .A(b[22]), .B(b[21]), .Y(n2340) );
  INVX1 U4247 ( .A(n2285), .Y(n4442) );
  AND2X1 U4248 ( .A(n5036), .B(n129), .Y(n2890) );
  INVX1 U4249 ( .A(n2890), .Y(n4443) );
  AND2X1 U4250 ( .A(n5036), .B(n96), .Y(n3091) );
  INVX1 U4251 ( .A(n3091), .Y(n4444) );
  BUFX2 U4252 ( .A(n3159), .Y(n4445) );
  AND2X1 U4253 ( .A(n5036), .B(n84), .Y(n3158) );
  INVX1 U4254 ( .A(n3158), .Y(n4446) );
  BUFX2 U4255 ( .A(n2958), .Y(n4447) );
  AND2X1 U4256 ( .A(n5035), .B(n4956), .Y(n3426) );
  INVX1 U4257 ( .A(n3426), .Y(n4448) );
  BUFX2 U4258 ( .A(n3561), .Y(n4449) );
  AND2X1 U4259 ( .A(n493), .B(n4516), .Y(n489) );
  INVX1 U4260 ( .A(n489), .Y(n4450) );
  BUFX2 U4261 ( .A(n490), .Y(n4451) );
  AND2X1 U4262 ( .A(n4544), .B(n2247), .Y(n2204) );
  INVX1 U4263 ( .A(n2204), .Y(n4452) );
  BUFX2 U4264 ( .A(n2249), .Y(n4453) );
  BUFX2 U4265 ( .A(n3427), .Y(n4454) );
  AND2X1 U4266 ( .A(n457), .B(n469), .Y(n451) );
  INVX1 U4267 ( .A(n451), .Y(n4455) );
  BUFX2 U4268 ( .A(n719), .Y(n4456) );
  AND2X1 U4269 ( .A(n4815), .B(n4817), .Y(n718) );
  INVX1 U4270 ( .A(n718), .Y(n4457) );
  BUFX2 U4271 ( .A(n483), .Y(n4458) );
  AND2X1 U4272 ( .A(n4676), .B(n2439), .Y(n2225) );
  INVX1 U4273 ( .A(n2225), .Y(n4459) );
  INVX1 U4274 ( .A(n279), .Y(n4460) );
  AND2X1 U4275 ( .A(n4481), .B(n2476), .Y(n2232) );
  INVX1 U4276 ( .A(n2232), .Y(n4461) );
  AND2X1 U4277 ( .A(n4683), .B(n2256), .Y(n2205) );
  INVX1 U4278 ( .A(n2205), .Y(n4462) );
  BUFX2 U4279 ( .A(n2260), .Y(n4463) );
  OR2X1 U4280 ( .A(n4689), .B(n4559), .Y(n440) );
  INVX1 U4281 ( .A(n440), .Y(n4464) );
  AND2X1 U4282 ( .A(n826), .B(n829), .Y(n322) );
  INVX1 U4283 ( .A(n322), .Y(n4465) );
  AND2X1 U4284 ( .A(n5035), .B(n60), .Y(n3292) );
  INVX1 U4285 ( .A(n3292), .Y(n4466) );
  BUFX2 U4286 ( .A(n3494), .Y(n4467) );
  BUFX2 U4287 ( .A(n610), .Y(n4468) );
  AND2X2 U4288 ( .A(n4915), .B(n4618), .Y(n407) );
  INVX1 U4289 ( .A(n407), .Y(n4469) );
  BUFX2 U4290 ( .A(n591), .Y(n4470) );
  AND2X1 U4291 ( .A(n4547), .B(n711), .Y(n284) );
  INVX1 U4292 ( .A(n284), .Y(n4471) );
  INVX1 U4293 ( .A(n280), .Y(n4472) );
  OR2X2 U4294 ( .A(n1409), .B(n1418), .Y(n4806) );
  AND2X1 U4295 ( .A(n4671), .B(n2470), .Y(n2231) );
  INVX1 U4296 ( .A(n2231), .Y(n4473) );
  AND2X1 U4297 ( .A(n4543), .B(n2315), .Y(n2210) );
  INVX1 U4298 ( .A(n2210), .Y(n4474) );
  BUFX2 U4299 ( .A(n2317), .Y(n4475) );
  AND2X1 U4300 ( .A(n4605), .B(n2434), .Y(n2224) );
  INVX1 U4301 ( .A(n2224), .Y(n4476) );
  BUFX2 U4302 ( .A(n2436), .Y(n4477) );
  AND2X1 U4303 ( .A(n4876), .B(n4910), .Y(n250) );
  INVX1 U4304 ( .A(n250), .Y(n4478) );
  AND2X1 U4305 ( .A(n4878), .B(n4912), .Y(n248) );
  INVX1 U4306 ( .A(n248), .Y(n4479) );
  OR2X1 U4307 ( .A(b[27]), .B(b[28]), .Y(n2280) );
  INVX1 U4308 ( .A(n2280), .Y(n4480) );
  AND2X1 U4309 ( .A(b[2]), .B(b[3]), .Y(n2477) );
  INVX1 U4310 ( .A(n2477), .Y(n4481) );
  INVX1 U4311 ( .A(n475), .Y(n4482) );
  AND2X1 U4312 ( .A(n837), .B(n842), .Y(n355) );
  INVX1 U4313 ( .A(n355), .Y(n4483) );
  OR2X1 U4314 ( .A(n1325), .B(n1338), .Y(n645) );
  INVX1 U4315 ( .A(n645), .Y(n4484) );
  INVX1 U4316 ( .A(n590), .Y(n4485) );
  AND2X1 U4317 ( .A(n5036), .B(n120), .Y(n2957) );
  INVX1 U4318 ( .A(n2957), .Y(n4486) );
  AND2X1 U4319 ( .A(n5035), .B(n72), .Y(n3225) );
  INVX1 U4320 ( .A(n3225), .Y(n4487) );
  BUFX2 U4321 ( .A(n3092), .Y(n4488) );
  BUFX2 U4322 ( .A(n637), .Y(n4489) );
  AND2X2 U4323 ( .A(n4903), .B(n4579), .Y(n636) );
  INVX1 U4324 ( .A(n636), .Y(n4490) );
  AND2X1 U4325 ( .A(n4597), .B(n4820), .Y(n288) );
  INVX1 U4326 ( .A(n288), .Y(n4491) );
  AND2X1 U4327 ( .A(n4724), .B(n4819), .Y(n290) );
  INVX1 U4328 ( .A(n290), .Y(n4492) );
  AND2X1 U4329 ( .A(n4545), .B(n744), .Y(n291) );
  INVX1 U4330 ( .A(n291), .Y(n4493) );
  AND2X1 U4331 ( .A(n4604), .B(n2404), .Y(n2220) );
  INVX1 U4332 ( .A(n2220), .Y(n4494) );
  BUFX2 U4333 ( .A(n2406), .Y(n4495) );
  AND2X1 U4334 ( .A(n4548), .B(n2446), .Y(n2226) );
  INVX1 U4335 ( .A(n2226), .Y(n4496) );
  AND2X1 U4336 ( .A(n4603), .B(n2293), .Y(n2208) );
  INVX1 U4337 ( .A(n2208), .Y(n4497) );
  BUFX2 U4338 ( .A(n2295), .Y(n4498) );
  AND2X1 U4339 ( .A(n4880), .B(n4914), .Y(n246) );
  INVX1 U4340 ( .A(n246), .Y(n4499) );
  AND2X1 U4341 ( .A(n4738), .B(n688), .Y(n281) );
  INVX1 U4342 ( .A(n281), .Y(n4500) );
  INVX1 U4343 ( .A(n257), .Y(n4501) );
  BUFX2 U4344 ( .A(n544), .Y(n4502) );
  INVX1 U4345 ( .A(n568), .Y(n4503) );
  OR2X1 U4346 ( .A(b[3]), .B(b[4]), .Y(n2470) );
  INVX1 U4347 ( .A(n2470), .Y(n4504) );
  INVX1 U4348 ( .A(n2302), .Y(n4505) );
  OR2X1 U4349 ( .A(b[9]), .B(b[10]), .Y(n2439) );
  INVX1 U4350 ( .A(n2439), .Y(n4506) );
  AND2X1 U4351 ( .A(n4916), .B(n4915), .Y(n400) );
  INVX1 U4352 ( .A(n400), .Y(n4507) );
  INVX1 U4353 ( .A(n594), .Y(n4508) );
  AND2X1 U4354 ( .A(n4913), .B(n4912), .Y(n457) );
  INVX1 U4355 ( .A(n457), .Y(n4509) );
  AND2X1 U4356 ( .A(b[28]), .B(b[29]), .Y(n2272) );
  INVX1 U4357 ( .A(n2272), .Y(n4510) );
  BUFX2 U4358 ( .A(n708), .Y(n4511) );
  OR2X1 U4359 ( .A(n4619), .B(n4681), .Y(n709) );
  INVX1 U4360 ( .A(n709), .Y(n4512) );
  BUFX2 U4361 ( .A(n2473), .Y(n4513) );
  OR2X1 U4362 ( .A(n4562), .B(n4624), .Y(n2474) );
  INVX1 U4363 ( .A(n2474), .Y(n4514) );
  OR2X1 U4364 ( .A(n4622), .B(n4756), .Y(n2245) );
  INVX1 U4365 ( .A(n2245), .Y(n4515) );
  OR2X1 U4366 ( .A(n3937), .B(n4625), .Y(n507) );
  INVX1 U4367 ( .A(n507), .Y(n4516) );
  AND2X1 U4368 ( .A(n824), .B(n825), .Y(n311) );
  INVX1 U4369 ( .A(n311), .Y(n4517) );
  OR2X1 U4370 ( .A(n832), .B(n830), .Y(n332) );
  INVX1 U4371 ( .A(n332), .Y(n4518) );
  OR2X1 U4372 ( .A(n842), .B(n837), .Y(n354) );
  INVX1 U4373 ( .A(n354), .Y(n4519) );
  AND2X1 U4374 ( .A(n1324), .B(n1311), .Y(n641) );
  INVX1 U4375 ( .A(n641), .Y(n4520) );
  INVX1 U4376 ( .A(n498), .Y(n4521) );
  AND2X1 U4377 ( .A(n887), .B(n895), .Y(n436) );
  INVX1 U4378 ( .A(n436), .Y(n4522) );
  INVX1 U4379 ( .A(n462), .Y(n4523) );
  INVX1 U4380 ( .A(n573), .Y(n4524) );
  INVX1 U4381 ( .A(n584), .Y(n4525) );
  BUFX2 U4382 ( .A(n2891), .Y(n4526) );
  AND2X1 U4383 ( .A(n4596), .B(n4818), .Y(n292) );
  INVX1 U4384 ( .A(n292), .Y(n4527) );
  AND2X1 U4385 ( .A(n4685), .B(n2479), .Y(n2233) );
  INVX1 U4386 ( .A(n2233), .Y(n4528) );
  AND2X1 U4387 ( .A(n4660), .B(n736), .Y(n289) );
  INVX1 U4388 ( .A(n289), .Y(n4529) );
  AND2X1 U4389 ( .A(n4602), .B(n2465), .Y(n2230) );
  INVX1 U4390 ( .A(n2230), .Y(n4530) );
  BUFX2 U4391 ( .A(n2467), .Y(n4531) );
  AND2X1 U4392 ( .A(n4600), .B(n2389), .Y(n2218) );
  INVX1 U4393 ( .A(n2218), .Y(n4532) );
  BUFX2 U4394 ( .A(n2391), .Y(n4533) );
  AND2X1 U4395 ( .A(n4684), .B(n2449), .Y(n2227) );
  INVX1 U4396 ( .A(n2227), .Y(n4534) );
  INVX1 U4397 ( .A(n258), .Y(n4535) );
  AND2X1 U4398 ( .A(n4885), .B(n4915), .Y(n243) );
  INVX1 U4399 ( .A(n243), .Y(n4536) );
  INVX1 U4400 ( .A(n259), .Y(n4537) );
  BUFX2 U4401 ( .A(n560), .Y(n4538) );
  AND2X1 U4402 ( .A(n1388), .B(n1377), .Y(n668) );
  INVX1 U4403 ( .A(n668), .Y(n4539) );
  INVX1 U4404 ( .A(n493), .Y(n4540) );
  OR2X2 U4405 ( .A(n1047), .B(n4841), .Y(n533) );
  OR2X1 U4406 ( .A(b[11]), .B(b[12]), .Y(n2423) );
  INVX1 U4407 ( .A(n2423), .Y(n4541) );
  OR2X1 U4408 ( .A(b[14]), .B(b[13]), .Y(n2409) );
  INVX1 U4409 ( .A(n2409), .Y(n4542) );
  INVX1 U4410 ( .A(n2316), .Y(n4543) );
  AND2X1 U4411 ( .A(b[30]), .B(n5035), .Y(n2248) );
  INVX1 U4412 ( .A(n2248), .Y(n4544) );
  AND2X1 U4413 ( .A(n1475), .B(n2885), .Y(n745) );
  INVX1 U4414 ( .A(n745), .Y(n4545) );
  AND2X1 U4415 ( .A(n1364), .B(n1353), .Y(n657) );
  INVX1 U4416 ( .A(n657), .Y(n4546) );
  AND2X1 U4417 ( .A(n1448), .B(n1443), .Y(n712) );
  INVX1 U4418 ( .A(n712), .Y(n4547) );
  AND2X1 U4419 ( .A(b[8]), .B(b[9]), .Y(n2447) );
  INVX1 U4420 ( .A(n2447), .Y(n4548) );
  AND2X2 U4421 ( .A(n1064), .B(n1048), .Y(n543) );
  INVX1 U4422 ( .A(n543), .Y(n4549) );
  AND2X1 U4423 ( .A(n4847), .B(n4846), .Y(n514) );
  INVX1 U4424 ( .A(n514), .Y(n4550) );
  BUFX2 U4425 ( .A(n730), .Y(n4551) );
  INVX1 U4426 ( .A(n587), .Y(n4552) );
  INVX1 U4427 ( .A(n556), .Y(n4553) );
  OR2X1 U4428 ( .A(n2265), .B(n4756), .Y(n2254) );
  INVX1 U4429 ( .A(n2254), .Y(n4554) );
  BUFX2 U4430 ( .A(n622), .Y(n4555) );
  OR2X1 U4431 ( .A(n370), .B(n350), .Y(n348) );
  INVX1 U4432 ( .A(n348), .Y(n4556) );
  INVX1 U4433 ( .A(n308), .Y(n4557) );
  BUFX2 U4434 ( .A(n682), .Y(n4558) );
  AND2X1 U4435 ( .A(n4914), .B(n457), .Y(n442) );
  INVX1 U4436 ( .A(n442), .Y(n4559) );
  INVX1 U4437 ( .A(n366), .Y(n4560) );
  AND2X1 U4438 ( .A(b[28]), .B(b[27]), .Y(n2281) );
  INVX1 U4439 ( .A(n2281), .Y(n4561) );
  OR2X1 U4440 ( .A(b[3]), .B(b[2]), .Y(n2476) );
  INVX1 U4441 ( .A(n2476), .Y(n4562) );
  AND2X1 U4442 ( .A(n833), .B(n836), .Y(n340) );
  INVX1 U4443 ( .A(n340), .Y(n4563) );
  OR2X1 U4444 ( .A(n825), .B(n824), .Y(n310) );
  INVX1 U4445 ( .A(n310), .Y(n4564) );
  AND2X1 U4446 ( .A(n843), .B(n847), .Y(n362) );
  INVX1 U4447 ( .A(n362), .Y(n4565) );
  AND2X1 U4448 ( .A(n868), .B(n862), .Y(n405) );
  INVX1 U4449 ( .A(n405), .Y(n4566) );
  AND2X1 U4450 ( .A(n1338), .B(n1325), .Y(n646) );
  INVX1 U4451 ( .A(n646), .Y(n4567) );
  INVX1 U4452 ( .A(n482), .Y(n4568) );
  OR2X1 U4453 ( .A(n886), .B(n877), .Y(n428) );
  INVX1 U4454 ( .A(n428), .Y(n4569) );
  AND2X1 U4455 ( .A(n1310), .B(n1295), .Y(n629) );
  INVX1 U4456 ( .A(n629), .Y(n4570) );
  INVX1 U4457 ( .A(n503), .Y(n4571) );
  INVX1 U4458 ( .A(n564), .Y(n4572) );
  AND2X1 U4459 ( .A(n1278), .B(n1263), .Y(n619) );
  INVX1 U4460 ( .A(n619), .Y(n4573) );
  INVX1 U4461 ( .A(n599), .Y(n4574) );
  INVX1 U4462 ( .A(n585), .Y(n4575) );
  INVX1 U4463 ( .A(n574), .Y(n4576) );
  AND2X1 U4464 ( .A(n5035), .B(n48), .Y(n3359) );
  INVX1 U4465 ( .A(n3359), .Y(n4577) );
  BUFX2 U4466 ( .A(n3293), .Y(n4578) );
  INVX1 U4467 ( .A(n643), .Y(n4579) );
  BUFX2 U4468 ( .A(n615), .Y(n4580) );
  BUFX2 U4469 ( .A(n600), .Y(n4581) );
  BUFX2 U4470 ( .A(n499), .Y(n4582) );
  INVX1 U4471 ( .A(n274), .Y(n4583) );
  AND2X1 U4472 ( .A(n4727), .B(n4816), .Y(n283) );
  INVX1 U4473 ( .A(n283), .Y(n4584) );
  AND2X1 U4474 ( .A(n4895), .B(n762), .Y(n236) );
  INVX1 U4475 ( .A(n236), .Y(n4585) );
  AND2X1 U4476 ( .A(n4674), .B(n2302), .Y(n2209) );
  INVX1 U4477 ( .A(n2209), .Y(n4586) );
  BUFX2 U4478 ( .A(n2304), .Y(n4587) );
  AND2X1 U4479 ( .A(n4678), .B(n518), .Y(n254) );
  AND2X1 U4480 ( .A(n4887), .B(n4917), .Y(n241) );
  INVX1 U4481 ( .A(n241), .Y(n4588) );
  AND2X1 U4482 ( .A(n4888), .B(n4918), .Y(n240) );
  INVX1 U4483 ( .A(n240), .Y(n4589) );
  AND2X1 U4484 ( .A(n4881), .B(n771), .Y(n245) );
  INVX1 U4485 ( .A(n245), .Y(n4590) );
  BUFX2 U4486 ( .A(n724), .Y(n4591) );
  AND2X1 U4487 ( .A(n4659), .B(n4817), .Y(n286) );
  INVX1 U4488 ( .A(n286), .Y(n4592) );
  AND2X1 U4489 ( .A(n4753), .B(n659), .Y(n276) );
  INVX1 U4490 ( .A(n276), .Y(n4593) );
  AND2X1 U4491 ( .A(n4879), .B(n4913), .Y(n247) );
  AND2X1 U4492 ( .A(n1434), .B(n1427), .Y(n701) );
  INVX1 U4493 ( .A(n701), .Y(n4594) );
  AND2X1 U4494 ( .A(n1398), .B(n1389), .Y(n673) );
  INVX1 U4495 ( .A(n673), .Y(n4595) );
  AND2X1 U4496 ( .A(n1477), .B(n2886), .Y(n750) );
  INVX1 U4497 ( .A(n750), .Y(n4596) );
  AND2X1 U4498 ( .A(n1468), .B(n1465), .Y(n734) );
  INVX1 U4499 ( .A(n734), .Y(n4597) );
  AND2X1 U4500 ( .A(n1418), .B(n1409), .Y(n686) );
  INVX1 U4501 ( .A(n686), .Y(n4598) );
  INVX1 U4502 ( .A(n571), .Y(n4599) );
  AND2X1 U4503 ( .A(b[16]), .B(b[17]), .Y(n2390) );
  INVX1 U4504 ( .A(n2390), .Y(n4600) );
  AND2X1 U4505 ( .A(b[12]), .B(b[13]), .Y(n2419) );
  INVX1 U4506 ( .A(n2419), .Y(n4601) );
  AND2X1 U4507 ( .A(b[4]), .B(b[5]), .Y(n2466) );
  INVX1 U4508 ( .A(n2466), .Y(n4602) );
  AND2X1 U4509 ( .A(b[26]), .B(b[27]), .Y(n2294) );
  INVX1 U4510 ( .A(n2294), .Y(n4603) );
  AND2X1 U4511 ( .A(b[14]), .B(b[15]), .Y(n2405) );
  INVX1 U4512 ( .A(n2405), .Y(n4604) );
  AND2X1 U4513 ( .A(b[10]), .B(b[11]), .Y(n2435) );
  INVX1 U4514 ( .A(n2435), .Y(n4605) );
  INVX1 U4515 ( .A(n559), .Y(n4606) );
  AND2X1 U4516 ( .A(n4843), .B(n4842), .Y(n529) );
  INVX1 U4517 ( .A(n529), .Y(n4607) );
  BUFX2 U4518 ( .A(n318), .Y(n4608) );
  OR2X2 U4519 ( .A(n1048), .B(n1064), .Y(n4762) );
  INVX1 U4520 ( .A(n4762), .Y(n4609) );
  AND2X2 U4521 ( .A(n4612), .B(n4552), .Y(n577) );
  INVX1 U4522 ( .A(n577), .Y(n4610) );
  BUFX2 U4523 ( .A(n578), .Y(n4611) );
  INVX1 U4524 ( .A(n579), .Y(n4612) );
  AND2X1 U4525 ( .A(n688), .B(n4806), .Y(n681) );
  INVX1 U4526 ( .A(n681), .Y(n4613) );
  AND2X1 U4527 ( .A(n4911), .B(n4910), .Y(n477) );
  INVX1 U4528 ( .A(n477), .Y(n4614) );
  INVX1 U4529 ( .A(n424), .Y(n4615) );
  AND2X1 U4530 ( .A(n758), .B(n754), .Y(n753) );
  INVX1 U4531 ( .A(n753), .Y(n4616) );
  BUFX2 U4532 ( .A(n738), .Y(n4617) );
  OR2X1 U4533 ( .A(n4689), .B(n420), .Y(n418) );
  INVX1 U4534 ( .A(n418), .Y(n4618) );
  OR2X1 U4535 ( .A(n1449), .B(n1454), .Y(n714) );
  INVX1 U4536 ( .A(n714), .Y(n4619) );
  OR2X1 U4537 ( .A(b[7]), .B(b[8]), .Y(n2449) );
  INVX1 U4538 ( .A(n2449), .Y(n4620) );
  INVX1 U4539 ( .A(n550), .Y(n4621) );
  INVX1 U4540 ( .A(n2247), .Y(n4622) );
  OR2X1 U4541 ( .A(n1353), .B(n1364), .Y(n656) );
  INVX1 U4542 ( .A(n656), .Y(n4623) );
  OR2X1 U4543 ( .A(b[1]), .B(b[2]), .Y(n2479) );
  INVX1 U4544 ( .A(n2479), .Y(n4624) );
  OR2X1 U4545 ( .A(n4846), .B(n4847), .Y(n513) );
  INVX1 U4546 ( .A(n513), .Y(n4625) );
  OR2X1 U4547 ( .A(b[29]), .B(b[28]), .Y(n2271) );
  INVX1 U4548 ( .A(n2271), .Y(n4626) );
  OR2X1 U4549 ( .A(b[25]), .B(b[24]), .Y(n2315) );
  INVX1 U4550 ( .A(n2315), .Y(n4627) );
  INVX1 U4551 ( .A(n370), .Y(n4628) );
  AND2X1 U4552 ( .A(n4725), .B(n4828), .Y(product[0]) );
  OR2X1 U4553 ( .A(n829), .B(n826), .Y(n321) );
  INVX1 U4554 ( .A(n321), .Y(n4629) );
  OR2X1 U4555 ( .A(n836), .B(n833), .Y(n339) );
  INVX1 U4556 ( .A(n339), .Y(n4630) );
  AND2X1 U4557 ( .A(n848), .B(n853), .Y(n381) );
  INVX1 U4558 ( .A(n381), .Y(n4631) );
  AND2X1 U4559 ( .A(n869), .B(n876), .Y(n414) );
  INVX1 U4560 ( .A(n414), .Y(n4632) );
  OR2X1 U4561 ( .A(n1339), .B(n1352), .Y(n650) );
  INVX1 U4562 ( .A(n650), .Y(n4633) );
  AND2X1 U4563 ( .A(n1294), .B(n1279), .Y(n626) );
  INVX1 U4564 ( .A(n626), .Y(n4634) );
  OR2X1 U4565 ( .A(n895), .B(n887), .Y(n435) );
  INVX1 U4566 ( .A(n435), .Y(n4635) );
  INVX1 U4567 ( .A(n604), .Y(n4636) );
  INVX1 U4568 ( .A(n589), .Y(n4637) );
  INVX1 U4569 ( .A(n581), .Y(n4638) );
  AND2X1 U4570 ( .A(n5035), .B(n4974), .Y(n3560) );
  INVX1 U4571 ( .A(n3560), .Y(n4639) );
  BUFX2 U4572 ( .A(n3360), .Y(n4640) );
  AND2X1 U4573 ( .A(n4752), .B(n714), .Y(n285) );
  INVX1 U4574 ( .A(n285), .Y(n4641) );
  AND2X1 U4575 ( .A(n4726), .B(n4815), .Y(n287) );
  INVX1 U4576 ( .A(n287), .Y(n4642) );
  INVX1 U4577 ( .A(n269), .Y(n4643) );
  AND2X1 U4578 ( .A(n4901), .B(n4919), .Y(n233) );
  INVX1 U4579 ( .A(n233), .Y(n4644) );
  INVX1 U4580 ( .A(n261), .Y(n4645) );
  AND2X1 U4581 ( .A(n4873), .B(n778), .Y(n252) );
  INVX1 U4582 ( .A(n252), .Y(n4646) );
  AND2X1 U4583 ( .A(n4883), .B(n770), .Y(n244) );
  INVX1 U4584 ( .A(n244), .Y(n4647) );
  AND2X1 U4585 ( .A(n4889), .B(n765), .Y(n239) );
  INVX1 U4586 ( .A(n239), .Y(n4648) );
  INVX1 U4587 ( .A(n282), .Y(n4649) );
  BUFX2 U4588 ( .A(n702), .Y(n4650) );
  INVX1 U4589 ( .A(n277), .Y(n4651) );
  BUFX2 U4590 ( .A(n669), .Y(n4652) );
  INVX1 U4591 ( .A(n272), .Y(n4653) );
  BUFX2 U4592 ( .A(n642), .Y(n4654) );
  INVX1 U4593 ( .A(n268), .Y(n4655) );
  AND2X1 U4594 ( .A(n4877), .B(n4911), .Y(n249) );
  INVX1 U4595 ( .A(n249), .Y(n4656) );
  INVX1 U4596 ( .A(n266), .Y(n4657) );
  OR2X1 U4597 ( .A(n4890), .B(n4892), .Y(n352) );
  INVX1 U4598 ( .A(n352), .Y(n4658) );
  AND2X1 U4599 ( .A(n1460), .B(n1455), .Y(n723) );
  INVX1 U4600 ( .A(n723), .Y(n4659) );
  OR2X2 U4601 ( .A(n1065), .B(n4835), .Y(n547) );
  AND2X1 U4602 ( .A(n2883), .B(n1469), .Y(n737) );
  INVX1 U4603 ( .A(n737), .Y(n4660) );
  AND2X1 U4604 ( .A(n1408), .B(n1399), .Y(n679) );
  INVX1 U4605 ( .A(n679), .Y(n4661) );
  OR2X1 U4606 ( .A(n1419), .B(n1426), .Y(n688) );
  INVX1 U4607 ( .A(n688), .Y(n4662) );
  BUFX2 U4608 ( .A(n458), .Y(n4663) );
  BUFX2 U4609 ( .A(n329), .Y(n4664) );
  BUFX2 U4610 ( .A(n494), .Y(n4665) );
  BUFX2 U4611 ( .A(n401), .Y(n4666) );
  AND2X2 U4612 ( .A(n797), .B(n4904), .Y(n621) );
  INVX1 U4613 ( .A(n621), .Y(n4667) );
  BUFX2 U4614 ( .A(n586), .Y(n4668) );
  BUFX2 U4615 ( .A(n746), .Y(n4669) );
  BUFX2 U4616 ( .A(n551), .Y(n4670) );
  AND2X1 U4617 ( .A(b[4]), .B(b[3]), .Y(n2471) );
  INVX1 U4618 ( .A(n2471), .Y(n4671) );
  AND2X1 U4619 ( .A(b[12]), .B(b[11]), .Y(n2424) );
  INVX1 U4620 ( .A(n2424), .Y(n4672) );
  AND2X1 U4621 ( .A(b[16]), .B(b[15]), .Y(n2395) );
  INVX1 U4622 ( .A(n2395), .Y(n4673) );
  INVX1 U4623 ( .A(n2303), .Y(n4674) );
  AND2X1 U4624 ( .A(b[13]), .B(b[14]), .Y(n2410) );
  INVX1 U4625 ( .A(n2410), .Y(n4675) );
  AND2X1 U4626 ( .A(b[10]), .B(b[9]), .Y(n2440) );
  INVX1 U4627 ( .A(n2440), .Y(n4676) );
  INVX1 U4628 ( .A(n534), .Y(n4677) );
  AND2X1 U4629 ( .A(n4845), .B(n4844), .Y(n519) );
  INVX1 U4630 ( .A(n519), .Y(n4678) );
  OR2X1 U4631 ( .A(b[5]), .B(b[6]), .Y(n2460) );
  INVX1 U4632 ( .A(n2460), .Y(n4679) );
  OR2X1 U4633 ( .A(n1365), .B(n1376), .Y(n659) );
  INVX1 U4634 ( .A(n659), .Y(n4680) );
  OR2X1 U4635 ( .A(n1443), .B(n1448), .Y(n711) );
  INVX1 U4636 ( .A(n711), .Y(n4681) );
  INVX1 U4637 ( .A(n2323), .Y(n4682) );
  AND2X1 U4638 ( .A(b[30]), .B(b[29]), .Y(n2259) );
  INVX1 U4639 ( .A(n2259), .Y(n4683) );
  AND2X1 U4640 ( .A(b[8]), .B(b[7]), .Y(n2450) );
  INVX1 U4641 ( .A(n2450), .Y(n4684) );
  AND2X1 U4642 ( .A(b[2]), .B(b[1]), .Y(n2480) );
  INVX1 U4643 ( .A(n2480), .Y(n4685) );
  OR2X2 U4644 ( .A(n4541), .B(n4748), .Y(n2414) );
  INVX1 U4645 ( .A(n2414), .Y(n4686) );
  INVX1 U4646 ( .A(n2265), .Y(n4687) );
  OR2X2 U4647 ( .A(n4615), .B(n4509), .Y(n231) );
  AND2X1 U4648 ( .A(n822), .B(n823), .Y(n300) );
  INVX1 U4649 ( .A(n300), .Y(n4690) );
  AND2X1 U4650 ( .A(n830), .B(n832), .Y(n333) );
  INVX1 U4651 ( .A(n333), .Y(n4691) );
  OR2X1 U4652 ( .A(n847), .B(n843), .Y(n361) );
  INVX1 U4653 ( .A(n361), .Y(n4692) );
  AND2X1 U4654 ( .A(n954), .B(n941), .Y(n487) );
  INVX1 U4655 ( .A(n487), .Y(n4693) );
  AND2X1 U4656 ( .A(n861), .B(n854), .Y(n390) );
  INVX1 U4657 ( .A(n390), .Y(n4694) );
  AND2X1 U4658 ( .A(n1352), .B(n1339), .Y(n651) );
  INVX1 U4659 ( .A(n651), .Y(n4695) );
  AND2X1 U4660 ( .A(n928), .B(n918), .Y(n467) );
  INVX1 U4661 ( .A(n467), .Y(n4696) );
  AND2X1 U4662 ( .A(n877), .B(n886), .Y(n429) );
  INVX1 U4663 ( .A(n429), .Y(n4697) );
  OR2X1 U4664 ( .A(n1295), .B(n1310), .Y(n628) );
  INVX1 U4665 ( .A(n628), .Y(n4698) );
  OR2X1 U4666 ( .A(n968), .B(n981), .Y(n502) );
  INVX1 U4667 ( .A(n502), .Y(n4699) );
  OR2X1 U4668 ( .A(n1101), .B(n1118), .Y(n563) );
  INVX1 U4669 ( .A(n563), .Y(n4700) );
  AND2X1 U4670 ( .A(n1262), .B(n1245), .Y(n614) );
  INVX1 U4671 ( .A(n614), .Y(n4701) );
  AND2X1 U4672 ( .A(n896), .B(n905), .Y(n449) );
  INVX1 U4673 ( .A(n449), .Y(n4702) );
  AND2X1 U4674 ( .A(n1172), .B(n1155), .Y(n582) );
  INVX1 U4675 ( .A(n582), .Y(n4703) );
  AND2X1 U4676 ( .A(n5036), .B(n108), .Y(n3024) );
  INVX1 U4677 ( .A(n3024), .Y(n4704) );
  AND2X1 U4678 ( .A(n5035), .B(n4965), .Y(n3493) );
  INVX1 U4679 ( .A(n3493), .Y(n4705) );
  BUFX2 U4680 ( .A(n3226), .Y(n4706) );
  OR2X2 U4681 ( .A(n4854), .B(n4852), .Y(n643) );
  INVX1 U4682 ( .A(n3939), .Y(n4707) );
  INVX1 U4683 ( .A(n278), .Y(n4708) );
  AND2X1 U4684 ( .A(n4897), .B(n761), .Y(n235) );
  INVX1 U4685 ( .A(n235), .Y(n4709) );
  AND2X1 U4686 ( .A(n4893), .B(n763), .Y(n237) );
  INVX1 U4687 ( .A(n237), .Y(n4710) );
  AND2X1 U4688 ( .A(n4899), .B(n760), .Y(n234) );
  INVX1 U4689 ( .A(n234), .Y(n4711) );
  AND2X1 U4690 ( .A(n4891), .B(n764), .Y(n238) );
  INVX1 U4691 ( .A(n238), .Y(n4712) );
  AND2X2 U4692 ( .A(n4861), .B(n4907), .Y(n267) );
  INVX1 U4693 ( .A(n267), .Y(n4713) );
  AND2X1 U4694 ( .A(n4858), .B(n4904), .Y(n270) );
  INVX1 U4695 ( .A(n270), .Y(n4714) );
  AND2X1 U4696 ( .A(n4886), .B(n4916), .Y(n242) );
  INVX1 U4697 ( .A(n242), .Y(n4715) );
  AND2X1 U4698 ( .A(n4871), .B(n786), .Y(n260) );
  INVX1 U4699 ( .A(n260), .Y(n4716) );
  AND2X1 U4700 ( .A(n4875), .B(n4909), .Y(n251) );
  INVX1 U4701 ( .A(n251), .Y(n4717) );
  BUFX2 U4702 ( .A(n647), .Y(n4718) );
  INVX1 U4703 ( .A(n273), .Y(n4719) );
  AND2X2 U4704 ( .A(n4856), .B(n797), .Y(n271) );
  INVX1 U4705 ( .A(n271), .Y(n4720) );
  AND2X1 U4706 ( .A(n4863), .B(n791), .Y(n265) );
  INVX1 U4707 ( .A(n265), .Y(n4721) );
  AND2X1 U4708 ( .A(n4869), .B(n788), .Y(n262) );
  INVX1 U4709 ( .A(n262), .Y(n4722) );
  AND2X1 U4710 ( .A(n4865), .B(n790), .Y(n264) );
  INVX1 U4711 ( .A(n264), .Y(n4723) );
  AND2X1 U4712 ( .A(n1473), .B(n2884), .Y(n742) );
  INVX1 U4713 ( .A(n742), .Y(n4724) );
  INVX1 U4714 ( .A(n758), .Y(n4725) );
  AND2X1 U4715 ( .A(n1461), .B(n1464), .Y(n728) );
  INVX1 U4716 ( .A(n728), .Y(n4726) );
  AND2X1 U4717 ( .A(n1442), .B(n1435), .Y(n706) );
  INVX1 U4718 ( .A(n706), .Y(n4727) );
  OR2X1 U4719 ( .A(n4844), .B(n4845), .Y(n518) );
  OR2X1 U4720 ( .A(n2885), .B(n1475), .Y(n744) );
  INVX1 U4721 ( .A(n744), .Y(n4728) );
  OR2X1 U4722 ( .A(n1469), .B(n2883), .Y(n736) );
  INVX1 U4723 ( .A(n736), .Y(n4729) );
  BUFX2 U4724 ( .A(n595), .Y(n4730) );
  OR2X1 U4725 ( .A(n4882), .B(n4884), .Y(n426) );
  INVX1 U4726 ( .A(n426), .Y(n4731) );
  INVX1 U4727 ( .A(n330), .Y(n4732) );
  BUFX2 U4728 ( .A(n606), .Y(n4733) );
  OR2X2 U4729 ( .A(n4735), .B(n4667), .Y(n607) );
  INVX1 U4730 ( .A(n607), .Y(n4734) );
  AND2X2 U4731 ( .A(n4905), .B(n4906), .Y(n609) );
  INVX1 U4732 ( .A(n609), .Y(n4735) );
  AND2X1 U4733 ( .A(n4918), .B(n4917), .Y(n376) );
  INVX1 U4734 ( .A(n376), .Y(n4736) );
  INVX1 U4735 ( .A(n751), .Y(n4737) );
  AND2X1 U4736 ( .A(n1426), .B(n1419), .Y(n689) );
  INVX1 U4737 ( .A(n689), .Y(n4738) );
  AND2X2 U4738 ( .A(n4835), .B(n1065), .Y(n548) );
  INVX1 U4739 ( .A(n548), .Y(n4739) );
  OR2X1 U4740 ( .A(n1399), .B(n1408), .Y(n678) );
  INVX1 U4741 ( .A(n678), .Y(n4740) );
  OR2X1 U4742 ( .A(b[15]), .B(b[14]), .Y(n2404) );
  INVX1 U4743 ( .A(n2404), .Y(n4741) );
  OR2X1 U4744 ( .A(n4831), .B(n4830), .Y(n570) );
  INVX1 U4745 ( .A(n570), .Y(n4742) );
  OR2X1 U4746 ( .A(n4834), .B(n4832), .Y(n558) );
  OR2X1 U4747 ( .A(b[7]), .B(b[6]), .Y(n2457) );
  INVX1 U4748 ( .A(n2457), .Y(n4744) );
  OR2X1 U4749 ( .A(b[27]), .B(b[26]), .Y(n2293) );
  INVX1 U4750 ( .A(n2293), .Y(n4745) );
  OR2X1 U4751 ( .A(b[5]), .B(b[4]), .Y(n2465) );
  INVX1 U4752 ( .A(n2465), .Y(n4746) );
  OR2X1 U4753 ( .A(b[17]), .B(b[16]), .Y(n2389) );
  INVX1 U4754 ( .A(n2389), .Y(n4747) );
  OR2X1 U4755 ( .A(b[13]), .B(b[12]), .Y(n2418) );
  INVX1 U4756 ( .A(n2418), .Y(n4748) );
  INVX1 U4757 ( .A(n2434), .Y(n4750) );
  OR2X1 U4758 ( .A(n4842), .B(n4843), .Y(n528) );
  INVX1 U4759 ( .A(n528), .Y(n4751) );
  AND2X1 U4760 ( .A(n1454), .B(n1449), .Y(n715) );
  INVX1 U4761 ( .A(n715), .Y(n4752) );
  AND2X1 U4762 ( .A(n1376), .B(n1365), .Y(n660) );
  INVX1 U4763 ( .A(n660), .Y(n4753) );
  OR2X1 U4764 ( .A(b[19]), .B(b[20]), .Y(n2358) );
  INVX1 U4765 ( .A(n2358), .Y(n4754) );
  INVX1 U4766 ( .A(n2320), .Y(n4755) );
  OR2X1 U4767 ( .A(b[29]), .B(b[30]), .Y(n2256) );
  INVX1 U4768 ( .A(n2256), .Y(n4756) );
  AND2X1 U4769 ( .A(b[0]), .B(b[1]), .Y(n2481) );
  INVX1 U4770 ( .A(n2481), .Y(n4757) );
  BUFX2 U4771 ( .A(n470), .Y(n4758) );
  BUFX2 U4772 ( .A(n478), .Y(n4759) );
  INVX1 U4773 ( .A(n575), .Y(n4760) );
  OAI21X1 U4774 ( .A(n568), .B(n3933), .C(n567), .Y(n4761) );
  INVX1 U4775 ( .A(n4954), .Y(n4953) );
  INVX1 U4776 ( .A(n4812), .Y(n4955) );
  INVX1 U4777 ( .A(n4950), .Y(n4949) );
  INVX1 U4778 ( .A(n4824), .Y(n4964) );
  INVX1 U4779 ( .A(n4958), .Y(n4957) );
  BUFX2 U4780 ( .A(n3932), .Y(n4764) );
  INVX1 U4781 ( .A(n4513), .Y(n2472) );
  INVX1 U4782 ( .A(n2445), .Y(n2443) );
  INVX1 U4783 ( .A(n2310), .Y(n2308) );
  XNOR2X1 U4784 ( .A(n4528), .B(n4757), .Y(n4765) );
  XNOR2X1 U4785 ( .A(n4364), .B(n4380), .Y(n4766) );
  XNOR2X1 U4786 ( .A(n4475), .B(n4474), .Y(n4767) );
  INVX1 U4787 ( .A(n662), .Y(n661) );
  XNOR2X1 U4788 ( .A(n4533), .B(n4532), .Y(n4768) );
  XNOR2X1 U4789 ( .A(n4372), .B(n4386), .Y(n4769) );
  OR2X1 U4790 ( .A(b[1]), .B(b[0]), .Y(n4770) );
  INVX1 U4791 ( .A(n2384), .Y(n2386) );
  INVX1 U4792 ( .A(n2266), .Y(n2268) );
  XNOR2X1 U4793 ( .A(n4369), .B(n4383), .Y(n4772) );
  XNOR2X1 U4794 ( .A(n4362), .B(n4379), .Y(n4773) );
  XNOR2X1 U4795 ( .A(n4370), .B(n4384), .Y(n4774) );
  XNOR2X1 U4796 ( .A(n4371), .B(n4385), .Y(n4775) );
  XNOR2X1 U4797 ( .A(n3959), .B(n4387), .Y(n4776) );
  XNOR2X1 U4798 ( .A(n4587), .B(n4586), .Y(n4777) );
  XNOR2X1 U4799 ( .A(n4498), .B(n4497), .Y(n4778) );
  XNOR2X1 U4800 ( .A(n4453), .B(n4452), .Y(n4779) );
  XNOR2X1 U4801 ( .A(n4463), .B(n4462), .Y(n4780) );
  XNOR2X1 U4802 ( .A(n4360), .B(n4376), .Y(n4781) );
  XNOR2X1 U4803 ( .A(n4477), .B(n4476), .Y(n4782) );
  XNOR2X1 U4804 ( .A(n4495), .B(n4494), .Y(n4783) );
  XNOR2X1 U4805 ( .A(n2451), .B(n4534), .Y(n4784) );
  INVX1 U4806 ( .A(n2452), .Y(n2451) );
  OR2X1 U4807 ( .A(n905), .B(n896), .Y(n4785) );
  OR2X1 U4808 ( .A(n876), .B(n869), .Y(n4786) );
  OR2X1 U4809 ( .A(n853), .B(n848), .Y(n4787) );
  INVX1 U4810 ( .A(n695), .Y(n694) );
  OR2X1 U4811 ( .A(n1311), .B(n1324), .Y(n4788) );
  OR2X1 U4812 ( .A(n1279), .B(n1294), .Y(n4789) );
  OR2X1 U4813 ( .A(n1263), .B(n1278), .Y(n4790) );
  OR2X1 U4814 ( .A(n1245), .B(n1262), .Y(n4791) );
  OR2X1 U4815 ( .A(n1227), .B(n1244), .Y(n4792) );
  OR2X1 U4816 ( .A(n1209), .B(n1226), .Y(n4793) );
  OR2X1 U4817 ( .A(n955), .B(n967), .Y(n4794) );
  OR2X1 U4818 ( .A(n941), .B(n954), .Y(n4795) );
  OR2X1 U4819 ( .A(n929), .B(n940), .Y(n4796) );
  OR2X1 U4820 ( .A(n918), .B(n928), .Y(n4797) );
  OR2X1 U4821 ( .A(n906), .B(n917), .Y(n4798) );
  OR2X1 U4822 ( .A(n862), .B(n868), .Y(n4799) );
  OR2X1 U4823 ( .A(n854), .B(n861), .Y(n4800) );
  INVX1 U4824 ( .A(n717), .Y(n716) );
  INVX1 U4825 ( .A(n1974), .Y(n1975) );
  INVX1 U4826 ( .A(n1848), .Y(n1849) );
  INVX1 U4827 ( .A(n2100), .Y(n2101) );
  INVX1 U4828 ( .A(n1722), .Y(n1723) );
  INVX1 U4829 ( .A(n4511), .Y(n707) );
  INVX1 U4830 ( .A(n4551), .Y(n729) );
  INVX1 U4831 ( .A(n4978), .Y(n4977) );
  INVX1 U4832 ( .A(n1978), .Y(n1979) );
  INVX1 U4833 ( .A(n1976), .Y(n1977) );
  INVX1 U4834 ( .A(n1852), .Y(n1853) );
  INVX1 U4835 ( .A(n1850), .Y(n1851) );
  INVX1 U4836 ( .A(n1726), .Y(n1727) );
  INVX1 U4837 ( .A(n1724), .Y(n1725) );
  INVX1 U4838 ( .A(n2167), .Y(n2168) );
  INVX1 U4839 ( .A(n2104), .Y(n2105) );
  INVX1 U4840 ( .A(n2102), .Y(n2103) );
  INVX1 U4841 ( .A(n1045), .Y(n1063) );
  INVX1 U4842 ( .A(n9), .Y(n4978) );
  INVX1 U4843 ( .A(n2058), .Y(n2059) );
  INVX1 U4844 ( .A(n2147), .Y(n2148) );
  INVX1 U4845 ( .A(n2139), .Y(n2140) );
  INVX1 U4846 ( .A(n2137), .Y(n2138) );
  INVX1 U4847 ( .A(n2145), .Y(n2146) );
  INVX1 U4848 ( .A(n2133), .Y(n2134) );
  INVX1 U4849 ( .A(n1995), .Y(n1996) );
  INVX1 U4850 ( .A(n2052), .Y(n2053) );
  INVX1 U4851 ( .A(n2054), .Y(n2055) );
  INVX1 U4852 ( .A(n2056), .Y(n2057) );
  INVX1 U4853 ( .A(n1997), .Y(n1998) );
  INVX1 U4854 ( .A(n1863), .Y(n1864) );
  INVX1 U4855 ( .A(n1920), .Y(n1921) );
  INVX1 U4856 ( .A(n1804), .Y(n1805) );
  INVX1 U4857 ( .A(n1861), .Y(n1862) );
  INVX1 U4858 ( .A(n1859), .Y(n1860) );
  INVX1 U4859 ( .A(n1802), .Y(n1803) );
  INVX1 U4860 ( .A(n1745), .Y(n1746) );
  INVX1 U4861 ( .A(n1857), .Y(n1858) );
  INVX1 U4862 ( .A(n1800), .Y(n1801) );
  INVX1 U4863 ( .A(n1743), .Y(n1744) );
  INVX1 U4864 ( .A(n1741), .Y(n1742) );
  INVX1 U4865 ( .A(n1798), .Y(n1799) );
  INVX1 U4866 ( .A(n1680), .Y(n1681) );
  INVX1 U4867 ( .A(n1737), .Y(n1738) );
  INVX1 U4868 ( .A(n1794), .Y(n1795) );
  INVX1 U4869 ( .A(n1796), .Y(n1797) );
  INVX1 U4870 ( .A(n1739), .Y(n1740) );
  INVX1 U4871 ( .A(n1930), .Y(n1931) );
  INVX1 U4872 ( .A(n1989), .Y(n1990) );
  INVX1 U4873 ( .A(n2048), .Y(n2049) );
  INVX1 U4874 ( .A(n1991), .Y(n1992) );
  INVX1 U4875 ( .A(n1934), .Y(n1935) );
  INVX1 U4876 ( .A(n2046), .Y(n2047) );
  INVX1 U4877 ( .A(n1924), .Y(n1925) );
  INVX1 U4878 ( .A(n1983), .Y(n1984) );
  INVX1 U4879 ( .A(n1926), .Y(n1927) );
  INVX1 U4880 ( .A(n1869), .Y(n1870) );
  INVX1 U4881 ( .A(n1865), .Y(n1866) );
  INVX1 U4882 ( .A(n1922), .Y(n1923) );
  INVX1 U4883 ( .A(n2050), .Y(n2051) );
  INVX1 U4884 ( .A(n1993), .Y(n1994) );
  INVX1 U4885 ( .A(n1682), .Y(n1683) );
  INVX1 U4886 ( .A(n1735), .Y(n1736) );
  INVX1 U4887 ( .A(n1733), .Y(n1734) );
  INVX1 U4888 ( .A(n1619), .Y(n1620) );
  INVX1 U4889 ( .A(n1617), .Y(n1618) );
  INVX1 U4890 ( .A(n1731), .Y(n1732) );
  INVX1 U4891 ( .A(n1672), .Y(n1673) );
  INVX1 U4892 ( .A(n1613), .Y(n1614) );
  INVX1 U4893 ( .A(n1670), .Y(n1671) );
  INVX1 U4894 ( .A(n1556), .Y(n1557) );
  INVX1 U4895 ( .A(n1554), .Y(n1555) );
  INVX1 U4896 ( .A(n1611), .Y(n1612) );
  INVX1 U4897 ( .A(n1668), .Y(n1669) );
  INVX1 U4898 ( .A(n1987), .Y(n1988) );
  INVX1 U4899 ( .A(n1985), .Y(n1986) );
  INVX1 U4900 ( .A(n1928), .Y(n1929) );
  INVX1 U4901 ( .A(n1871), .Y(n1872) );
  INVX1 U4902 ( .A(n1609), .Y(n1610) );
  INVX1 U4903 ( .A(n1607), .Y(n1608) );
  INVX1 U4904 ( .A(n1605), .Y(n1606) );
  INVX1 U4905 ( .A(n1546), .Y(n1547) );
  INVX1 U4906 ( .A(n2092), .Y(n2093) );
  INVX1 U4907 ( .A(n2090), .Y(n2091) );
  INVX1 U4908 ( .A(n2155), .Y(n2156) );
  INVX1 U4909 ( .A(n2025), .Y(n2026) );
  INVX1 U4910 ( .A(n1966), .Y(n1967) );
  INVX1 U4911 ( .A(n2029), .Y(n2030) );
  INVX1 U4912 ( .A(n2084), .Y(n2085) );
  INVX1 U4913 ( .A(n2027), .Y(n2028) );
  INVX1 U4914 ( .A(n2023), .Y(n2024) );
  INVX1 U4915 ( .A(n2080), .Y(n2081) );
  INVX1 U4916 ( .A(n1598), .Y(n1599) );
  INVX1 U4917 ( .A(n2086), .Y(n2087) );
  INVX1 U4918 ( .A(n1962), .Y(n1963) );
  INVX1 U4919 ( .A(n2021), .Y(n2022) );
  INVX1 U4920 ( .A(n1964), .Y(n1965) );
  INVX1 U4921 ( .A(n2076), .Y(n2077) );
  INVX1 U4922 ( .A(n1840), .Y(n1841) );
  INVX1 U4923 ( .A(n1777), .Y(n1778) );
  INVX1 U4924 ( .A(n1651), .Y(n1652) );
  INVX1 U4925 ( .A(n1824), .Y(n1825) );
  INVX1 U4926 ( .A(n1596), .Y(n1597) );
  INVX1 U4927 ( .A(n1714), .Y(n1715) );
  INVX1 U4928 ( .A(n1769), .Y(n1770) );
  INVX1 U4929 ( .A(n1712), .Y(n1713) );
  INVX1 U4930 ( .A(n1580), .Y(n1581) );
  INVX1 U4931 ( .A(n1706), .Y(n1707) );
  INVX1 U4932 ( .A(n1818), .Y(n1819) );
  INVX1 U4933 ( .A(n1761), .Y(n1762) );
  INVX1 U4934 ( .A(n1647), .Y(n1648) );
  INVX1 U4935 ( .A(n1649), .Y(n1650) );
  INVX1 U4936 ( .A(n1588), .Y(n1589) );
  INVX1 U4937 ( .A(n1698), .Y(n1699) );
  INVX1 U4938 ( .A(n1903), .Y(n1904) );
  INVX1 U4939 ( .A(n1901), .Y(n1902) );
  INVX1 U4940 ( .A(n2070), .Y(n2071) );
  INVX1 U4941 ( .A(n1820), .Y(n1821) );
  INVX1 U4942 ( .A(n1958), .Y(n1959) );
  INVX1 U4943 ( .A(n1956), .Y(n1957) );
  INVX1 U4944 ( .A(n2013), .Y(n2014) );
  INVX1 U4945 ( .A(n2011), .Y(n2012) );
  INVX1 U4946 ( .A(n1954), .Y(n1955) );
  INVX1 U4947 ( .A(n2009), .Y(n2010) );
  INVX1 U4948 ( .A(n2125), .Y(n2126) );
  INVX1 U4949 ( .A(n1895), .Y(n1896) );
  INVX1 U4950 ( .A(n1838), .Y(n1839) );
  INVX1 U4951 ( .A(n2121), .Y(n2122) );
  INVX1 U4952 ( .A(n2007), .Y(n2008) );
  INVX1 U4953 ( .A(n1893), .Y(n1894) );
  INVX1 U4954 ( .A(n1950), .Y(n1951) );
  INVX1 U4955 ( .A(n2062), .Y(n2063) );
  INVX1 U4956 ( .A(n2119), .Y(n2120) );
  INVX1 U4957 ( .A(n1948), .Y(n1949) );
  INVX1 U4958 ( .A(n1891), .Y(n1892) );
  INVX1 U4959 ( .A(n2117), .Y(n2118) );
  INVX1 U4960 ( .A(n1946), .Y(n1947) );
  INVX1 U4961 ( .A(n1775), .Y(n1776) );
  INVX1 U4962 ( .A(n1832), .Y(n1833) );
  INVX1 U4963 ( .A(n2115), .Y(n2116) );
  INVX1 U4964 ( .A(n1944), .Y(n1945) );
  INVX1 U4965 ( .A(n1830), .Y(n1831) );
  INVX1 U4966 ( .A(n1887), .Y(n1888) );
  INVX1 U4967 ( .A(n1936), .Y(n1937) );
  INVX1 U4968 ( .A(n1822), .Y(n1823) );
  INVX1 U4969 ( .A(n1765), .Y(n1766) );
  INVX1 U4970 ( .A(n2109), .Y(n2110) );
  INVX1 U4971 ( .A(n1885), .Y(n1886) );
  INVX1 U4972 ( .A(n1828), .Y(n1829) );
  INVX1 U4973 ( .A(n2111), .Y(n2112) );
  INVX1 U4974 ( .A(n2113), .Y(n2114) );
  INVX1 U4975 ( .A(n1881), .Y(n1882) );
  INVX1 U4976 ( .A(n1767), .Y(n1768) );
  INVX1 U4977 ( .A(n1692), .Y(n1693) );
  INVX1 U4978 ( .A(n1635), .Y(n1636) );
  INVX1 U4979 ( .A(n1633), .Y(n1634) );
  INVX1 U4980 ( .A(n1747), .Y(n1748) );
  INVX1 U4981 ( .A(n1631), .Y(n1632) );
  INVX1 U4982 ( .A(n1574), .Y(n1575) );
  INVX1 U4983 ( .A(n1629), .Y(n1630) );
  INVX1 U4984 ( .A(n1873), .Y(n1874) );
  INVX1 U4985 ( .A(n1704), .Y(n1705) );
  INVX1 U4986 ( .A(n1759), .Y(n1760) );
  INVX1 U4987 ( .A(n1702), .Y(n1703) );
  INVX1 U4988 ( .A(n1643), .Y(n1644) );
  INVX1 U4989 ( .A(n1810), .Y(n1811) );
  INVX1 U4990 ( .A(n1696), .Y(n1697) );
  INVX1 U4991 ( .A(n1755), .Y(n1756) );
  INVX1 U4992 ( .A(n1641), .Y(n1642) );
  INVX1 U4993 ( .A(n1694), .Y(n1695) );
  INVX1 U4994 ( .A(n1582), .Y(n1583) );
  INVX1 U4995 ( .A(n1637), .Y(n1638) );
  INVX1 U4996 ( .A(n2074), .Y(n2075) );
  INVX1 U4997 ( .A(n2017), .Y(n2018) );
  INVX1 U4998 ( .A(n2153), .Y(n2154) );
  INVX1 U4999 ( .A(n1757), .Y(n1758) );
  INVX1 U5000 ( .A(n1700), .Y(n1701) );
  INVX1 U5001 ( .A(n952), .Y(n966) );
  XNOR2X1 U5002 ( .A(n4531), .B(n4530), .Y(n4801) );
  INVX1 U5003 ( .A(n840), .Y(n846) );
  INVX1 U5004 ( .A(n915), .Y(n927) );
  INVX1 U5005 ( .A(n884), .Y(n894) );
  INVX1 U5006 ( .A(n859), .Y(n867) );
  INVX1 U5007 ( .A(n995), .Y(n996) );
  INVX1 U5008 ( .A(n827), .Y(n831) );
  XNOR2X1 U5009 ( .A(n4421), .B(n4373), .Y(n4802) );
  XNOR2X1 U5010 ( .A(n4366), .B(n4381), .Y(n4803) );
  XNOR2X1 U5011 ( .A(n4367), .B(n4382), .Y(n4804) );
  INVX1 U5012 ( .A(n821), .Y(n822) );
  INVX1 U5013 ( .A(n1911), .Y(n1912) );
  INVX1 U5014 ( .A(n1899), .Y(n1900) );
  INVX1 U5015 ( .A(n1897), .Y(n1898) );
  INVX1 U5016 ( .A(n1952), .Y(n1953) );
  INVX1 U5017 ( .A(n1836), .Y(n1837) );
  INVX1 U5018 ( .A(n1834), .Y(n1835) );
  INVX1 U5019 ( .A(n1889), .Y(n1890) );
  INVX1 U5020 ( .A(n1826), .Y(n1827) );
  INVX1 U5021 ( .A(n1883), .Y(n1884) );
  INVX1 U5022 ( .A(n1806), .Y(n1807) );
  INVX1 U5023 ( .A(n1932), .Y(n1933) );
  INVX1 U5024 ( .A(n2037), .Y(n2038) );
  INVX1 U5025 ( .A(n2143), .Y(n2144) );
  INVX1 U5026 ( .A(n2088), .Y(n2089) );
  INVX1 U5027 ( .A(n1710), .Y(n1711) );
  INVX1 U5028 ( .A(n1659), .Y(n1660) );
  INVX1 U5029 ( .A(n1584), .Y(n1585) );
  INVX1 U5030 ( .A(n1785), .Y(n1786) );
  INVX1 U5031 ( .A(n1773), .Y(n1774) );
  INVX1 U5032 ( .A(n1576), .Y(n1577) );
  INVX1 U5033 ( .A(n2072), .Y(n2073) );
  INVX1 U5034 ( .A(n1568), .Y(n1569) );
  INVX1 U5035 ( .A(n1615), .Y(n1616) );
  INVX1 U5036 ( .A(n1552), .Y(n1553) );
  INVX1 U5037 ( .A(n1548), .Y(n1549) );
  INVX1 U5038 ( .A(n2123), .Y(n2124) );
  INVX1 U5039 ( .A(n1999), .Y(n2000) );
  INVX1 U5040 ( .A(n1684), .Y(n1685) );
  INVX1 U5041 ( .A(n1763), .Y(n1764) );
  INVX1 U5042 ( .A(n1558), .Y(n1559) );
  INVX1 U5043 ( .A(n2019), .Y(n2020) );
  INVX1 U5044 ( .A(n1708), .Y(n1709) );
  INVX1 U5045 ( .A(n1771), .Y(n1772) );
  INVX1 U5046 ( .A(n1578), .Y(n1579) );
  INVX1 U5047 ( .A(n1586), .Y(n1587) );
  INVX1 U5048 ( .A(n1566), .Y(n1567) );
  INVX1 U5049 ( .A(n1645), .Y(n1646) );
  INVX1 U5050 ( .A(n1550), .Y(n1551) );
  INVX1 U5051 ( .A(n4967), .Y(n4965) );
  INVX1 U5052 ( .A(n4967), .Y(n4966) );
  INVX1 U5053 ( .A(n4976), .Y(n4974) );
  INVX1 U5054 ( .A(n4976), .Y(n4975) );
  INVX1 U5055 ( .A(n4810), .Y(n4972) );
  INVX1 U5056 ( .A(n4810), .Y(n4973) );
  INVX1 U5057 ( .A(n4811), .Y(n4980) );
  INVX1 U5058 ( .A(n4811), .Y(n4979) );
  INVX1 U5059 ( .A(n4969), .Y(n4968) );
  INVX1 U5060 ( .A(n4937), .Y(n4936) );
  INVX1 U5061 ( .A(n4943), .Y(n4942) );
  INVX1 U5062 ( .A(n4952), .Y(n4951) );
  INVX1 U5063 ( .A(n1663), .Y(n1664) );
  INVX1 U5064 ( .A(n1661), .Y(n1662) );
  INVX1 U5065 ( .A(n2041), .Y(n2042) );
  INVX1 U5066 ( .A(n1915), .Y(n1916) );
  INVX1 U5067 ( .A(n1913), .Y(n1914) );
  INVX1 U5068 ( .A(n1789), .Y(n1790) );
  INVX1 U5069 ( .A(n1787), .Y(n1788) );
  INVX1 U5070 ( .A(n2039), .Y(n2040) );
  INVX1 U5071 ( .A(n2149), .Y(n2150) );
  INVX1 U5072 ( .A(n2141), .Y(n2142) );
  INVX1 U5073 ( .A(n2135), .Y(n2136) );
  INVX1 U5074 ( .A(n2151), .Y(n2152) );
  INVX1 U5075 ( .A(n1678), .Y(n1679) );
  INVX1 U5076 ( .A(n1867), .Y(n1868) );
  INVX1 U5077 ( .A(n1676), .Y(n1677) );
  INVX1 U5078 ( .A(n1674), .Y(n1675) );
  INVX1 U5079 ( .A(n2082), .Y(n2083) );
  INVX1 U5080 ( .A(n2078), .Y(n2079) );
  INVX1 U5081 ( .A(n2064), .Y(n2065) );
  INVX1 U5082 ( .A(n2060), .Y(n2061) );
  INVX1 U5083 ( .A(n1600), .Y(n1601) );
  INVX1 U5084 ( .A(n1639), .Y(n1640) );
  INVX1 U5085 ( .A(n1572), .Y(n1573) );
  INVX1 U5086 ( .A(n1570), .Y(n1571) );
  INVX1 U5087 ( .A(n1621), .Y(n1622) );
  INVX1 U5088 ( .A(n1960), .Y(n1961) );
  INVX1 U5089 ( .A(n2015), .Y(n2016) );
  INVX1 U5090 ( .A(n1808), .Y(n1809) );
  INVX1 U5091 ( .A(n4971), .Y(n4970) );
  INVX1 U5092 ( .A(n4982), .Y(n4981) );
  OR2X1 U5093 ( .A(n1389), .B(n1398), .Y(n4805) );
  OR2X1 U5094 ( .A(n1427), .B(n1434), .Y(n4807) );
  INVX1 U5095 ( .A(n5037), .Y(n5035) );
  INVX1 U5096 ( .A(n5014), .Y(n5013) );
  INVX1 U5097 ( .A(n4992), .Y(n4991) );
  INVX1 U5098 ( .A(n5016), .Y(n5015) );
  INVX1 U5099 ( .A(n4984), .Y(n4983) );
  INVX1 U5100 ( .A(n4986), .Y(n4985) );
  INVX1 U5101 ( .A(n4996), .Y(n4995) );
  INVX1 U5102 ( .A(n4814), .Y(n4938) );
  INVX1 U5103 ( .A(n5022), .Y(n5021) );
  INVX1 U5104 ( .A(n5024), .Y(n5023) );
  INVX1 U5105 ( .A(n4998), .Y(n4997) );
  INVX1 U5106 ( .A(n5012), .Y(n5011) );
  INVX1 U5107 ( .A(n4988), .Y(n4987) );
  INVX1 U5108 ( .A(n1544), .Y(n1545) );
  INVX1 U5109 ( .A(n1542), .Y(n1543) );
  INVX1 U5110 ( .A(n1489), .Y(n1490) );
  INVX1 U5111 ( .A(n1525), .Y(n1526) );
  INVX1 U5112 ( .A(n1519), .Y(n1520) );
  INVX1 U5113 ( .A(n1517), .Y(n1518) );
  INVX1 U5114 ( .A(n1507), .Y(n1508) );
  INVX1 U5115 ( .A(n1501), .Y(n1502) );
  INVX1 U5116 ( .A(n1495), .Y(n1496) );
  INVX1 U5117 ( .A(n1483), .Y(n1484) );
  INVX1 U5118 ( .A(n1513), .Y(n1514) );
  INVX1 U5119 ( .A(b[16]), .Y(n5012) );
  INVX1 U5120 ( .A(n24), .Y(n4967) );
  AND2X1 U5121 ( .A(n3701), .B(n3723), .Y(n2198) );
  INVX1 U5122 ( .A(n1011), .Y(n1012) );
  INVX1 U5123 ( .A(n2131), .Y(n2132) );
  INVX1 U5124 ( .A(n2129), .Y(n2130) );
  INVX1 U5125 ( .A(n2094), .Y(n2095) );
  INVX1 U5126 ( .A(n2033), .Y(n2034) );
  INVX1 U5127 ( .A(n1970), .Y(n1971) );
  INVX1 U5128 ( .A(n2031), .Y(n2032) );
  INVX1 U5129 ( .A(n1907), .Y(n1908) );
  INVX1 U5130 ( .A(n2157), .Y(n2158) );
  INVX1 U5131 ( .A(n1594), .Y(n1595) );
  INVX1 U5132 ( .A(n1653), .Y(n1654) );
  INVX1 U5133 ( .A(n1716), .Y(n1717) );
  INVX1 U5134 ( .A(n1655), .Y(n1656) );
  INVX1 U5135 ( .A(n1590), .Y(n1591) );
  INVX1 U5136 ( .A(n1592), .Y(n1593) );
  INVX1 U5137 ( .A(n1844), .Y(n1845) );
  INVX1 U5138 ( .A(n2127), .Y(n2128) );
  INVX1 U5139 ( .A(n1842), .Y(n1843) );
  INVX1 U5140 ( .A(n2068), .Y(n2069) );
  INVX1 U5141 ( .A(n2066), .Y(n2067) );
  INVX1 U5142 ( .A(n1781), .Y(n1782) );
  INVX1 U5143 ( .A(n1779), .Y(n1780) );
  INVX1 U5144 ( .A(n1718), .Y(n1719) );
  INVX1 U5145 ( .A(n1879), .Y(n1880) );
  INVX1 U5146 ( .A(n1942), .Y(n1943) );
  INVX1 U5147 ( .A(n1938), .Y(n1939) );
  INVX1 U5148 ( .A(n1749), .Y(n1750) );
  INVX1 U5149 ( .A(n1690), .Y(n1691) );
  INVX1 U5150 ( .A(n1688), .Y(n1689) );
  INVX1 U5151 ( .A(n1686), .Y(n1687) );
  INVX1 U5152 ( .A(n1627), .Y(n1628) );
  INVX1 U5153 ( .A(n1625), .Y(n1626) );
  INVX1 U5154 ( .A(n1877), .Y(n1878) );
  INVX1 U5155 ( .A(n1875), .Y(n1876) );
  INVX1 U5156 ( .A(n1816), .Y(n1817) );
  INVX1 U5157 ( .A(n1812), .Y(n1813) );
  INVX1 U5158 ( .A(n1751), .Y(n1752) );
  INVX1 U5159 ( .A(n1753), .Y(n1754) );
  INVX1 U5160 ( .A(n1623), .Y(n1624) );
  INVX1 U5161 ( .A(n1564), .Y(n1565) );
  INVX1 U5162 ( .A(n1562), .Y(n1563) );
  INVX1 U5163 ( .A(n1560), .Y(n1561) );
  INVX1 U5164 ( .A(n1814), .Y(n1815) );
  INVX1 U5165 ( .A(n1521), .Y(n1522) );
  INVX1 U5166 ( .A(n1540), .Y(n2922) );
  XNOR2X1 U5167 ( .A(n2516), .B(n821), .Y(n232) );
  INVX1 U5168 ( .A(n5050), .Y(n5049) );
  INVX1 U5169 ( .A(n5047), .Y(n5046) );
  INVX1 U5170 ( .A(n5047), .Y(n5045) );
  INVX1 U5171 ( .A(n5050), .Y(n5048) );
  XNOR2X1 U5172 ( .A(n2238), .B(b[31]), .Y(n4809) );
  INVX1 U5173 ( .A(n16), .Y(n4971) );
  INVX1 U5174 ( .A(n3712), .Y(n2200) );
  INVX1 U5175 ( .A(n40), .Y(n4954) );
  INVX1 U5176 ( .A(n3710), .Y(n2194) );
  INVX1 U5177 ( .A(n3706), .Y(n2182) );
  AND2X1 U5178 ( .A(n3695), .B(n3717), .Y(n2180) );
  AND2X1 U5179 ( .A(n3697), .B(n3719), .Y(n2186) );
  INVX1 U5180 ( .A(n48), .Y(n4950) );
  AND2X1 U5181 ( .A(n3699), .B(n3721), .Y(n2192) );
  INVX1 U5182 ( .A(n12), .Y(n4976) );
  INVX1 U5183 ( .A(a[0]), .Y(n3702) );
  OR2X1 U5184 ( .A(n3701), .B(n3723), .Y(n4810) );
  OR2X1 U5185 ( .A(n3724), .B(n3702), .Y(n4811) );
  OR2X1 U5186 ( .A(n3721), .B(n3699), .Y(n4812) );
  OR2X1 U5187 ( .A(n3717), .B(n3695), .Y(n4814) );
  INVX1 U5188 ( .A(b[2]), .Y(n4984) );
  INVX1 U5189 ( .A(n2044), .Y(n3458) );
  INVX1 U5190 ( .A(n1981), .Y(n3391) );
  INVX1 U5191 ( .A(n22), .Y(n4969) );
  INVX1 U5192 ( .A(n3723), .Y(n2199) );
  INVX1 U5193 ( .A(n94), .Y(n4937) );
  INVX1 U5194 ( .A(n3717), .Y(n2181) );
  INVX1 U5195 ( .A(n70), .Y(n4943) );
  INVX1 U5196 ( .A(n3719), .Y(n2187) );
  INVX1 U5197 ( .A(n46), .Y(n4952) );
  INVX1 U5198 ( .A(n3721), .Y(n2193) );
  INVX1 U5199 ( .A(n1537), .Y(n1538) );
  INVX1 U5200 ( .A(n1968), .Y(n1969) );
  INVX1 U5201 ( .A(n1909), .Y(n1910) );
  INVX1 U5202 ( .A(n1972), .Y(n1973) );
  INVX1 U5203 ( .A(n1905), .Y(n1906) );
  INVX1 U5204 ( .A(n1846), .Y(n1847) );
  INVX1 U5205 ( .A(n1940), .Y(n1941) );
  INVX1 U5206 ( .A(n1535), .Y(n1536) );
  INVX1 U5207 ( .A(n1515), .Y(n1516) );
  INVX1 U5208 ( .A(n1487), .Y(n1488) );
  INVX1 U5209 ( .A(n2001), .Y(n2002) );
  INVX1 U5210 ( .A(n2096), .Y(n2097) );
  INVX1 U5211 ( .A(n2098), .Y(n2099) );
  INVX1 U5212 ( .A(n2035), .Y(n2036) );
  INVX1 U5213 ( .A(n1783), .Y(n1784) );
  INVX1 U5214 ( .A(n1720), .Y(n1721) );
  INVX1 U5215 ( .A(n1657), .Y(n1658) );
  INVX1 U5216 ( .A(n2003), .Y(n2004) );
  INVX1 U5217 ( .A(n4962), .Y(n4961) );
  INVX1 U5218 ( .A(n4958), .Y(n4956) );
  INVX1 U5219 ( .A(n4927), .Y(n4926) );
  INVX1 U5220 ( .A(n4826), .Y(n4931) );
  INVX1 U5221 ( .A(n4826), .Y(n4932) );
  INVX1 U5222 ( .A(n3724), .Y(n2202) );
  INVX1 U5223 ( .A(n4825), .Y(n4941) );
  INVX1 U5224 ( .A(n4824), .Y(n4963) );
  INVX1 U5225 ( .A(n4822), .Y(n4947) );
  INVX1 U5226 ( .A(n4946), .Y(n4945) );
  INVX1 U5227 ( .A(n4940), .Y(n4939) );
  INVX1 U5228 ( .A(n4960), .Y(n4959) );
  INVX1 U5229 ( .A(n4934), .Y(n4933) );
  INVX1 U5230 ( .A(n4930), .Y(n4929) );
  INVX1 U5231 ( .A(n3708), .Y(n2188) );
  INVX1 U5232 ( .A(n1527), .Y(n1528) );
  INVX1 U5233 ( .A(n1523), .Y(n1524) );
  INVX1 U5234 ( .A(n1533), .Y(n1534) );
  INVX1 U5235 ( .A(n1531), .Y(n1532) );
  INVX1 U5236 ( .A(n1511), .Y(n1512) );
  INVX1 U5237 ( .A(n1505), .Y(n1506) );
  INVX1 U5238 ( .A(n1529), .Y(n1530) );
  INVX1 U5239 ( .A(n1499), .Y(n1500) );
  INVX1 U5240 ( .A(n1493), .Y(n1494) );
  INVX1 U5241 ( .A(n2005), .Y(n2006) );
  OR2X1 U5242 ( .A(n1464), .B(n1461), .Y(n4815) );
  OR2X1 U5243 ( .A(n1435), .B(n1442), .Y(n4816) );
  OR2X1 U5244 ( .A(n1455), .B(n1460), .Y(n4817) );
  INVX1 U5245 ( .A(n4994), .Y(n4993) );
  INVX1 U5246 ( .A(n5002), .Y(n5001) );
  INVX1 U5247 ( .A(n5004), .Y(n5003) );
  INVX1 U5248 ( .A(n5006), .Y(n5005) );
  INVX1 U5249 ( .A(n5020), .Y(n5019) );
  INVX1 U5250 ( .A(n5008), .Y(n5007) );
  INVX1 U5251 ( .A(n5018), .Y(n5017) );
  INVX1 U5252 ( .A(n5026), .Y(n5025) );
  INVX1 U5253 ( .A(n5030), .Y(n5029) );
  INVX1 U5254 ( .A(n5032), .Y(n5031) );
  INVX1 U5255 ( .A(n4822), .Y(n4948) );
  INVX1 U5256 ( .A(n5000), .Y(n4999) );
  INVX1 U5257 ( .A(n5034), .Y(n5033) );
  INVX1 U5258 ( .A(n5028), .Y(n5027) );
  OR2X1 U5259 ( .A(n2886), .B(n1477), .Y(n4818) );
  OR2X1 U5260 ( .A(n2884), .B(n1473), .Y(n4819) );
  OR2X1 U5261 ( .A(n1465), .B(n1468), .Y(n4820) );
  INVX1 U5262 ( .A(n4823), .Y(n4935) );
  INVX1 U5263 ( .A(b[31]), .Y(n5037) );
  INVX1 U5264 ( .A(b[0]), .Y(n4982) );
  OR2X1 U5265 ( .A(n823), .B(n822), .Y(n4821) );
  INVX1 U5266 ( .A(b[4]), .Y(n4988) );
  INVX1 U5267 ( .A(b[19]), .Y(n5016) );
  INVX1 U5268 ( .A(b[24]), .Y(n5022) );
  INVX1 U5269 ( .A(b[25]), .Y(n5024) );
  INVX1 U5270 ( .A(b[6]), .Y(n4992) );
  INVX1 U5271 ( .A(b[3]), .Y(n4986) );
  INVX1 U5272 ( .A(b[8]), .Y(n4996) );
  XOR2X1 U5273 ( .A(n754), .B(n758), .Y(product[1]) );
  INVX1 U5274 ( .A(n1481), .Y(n1482) );
  INVX1 U5275 ( .A(n1479), .Y(n1480) );
  INVX1 U5276 ( .A(b[15]), .Y(n5010) );
  INVX1 U5277 ( .A(n1497), .Y(n1498) );
  INVX1 U5278 ( .A(n1509), .Y(n1510) );
  INVX1 U5279 ( .A(n1485), .Y(n1486) );
  INVX1 U5280 ( .A(n1503), .Y(n1504) );
  INVX1 U5281 ( .A(n82), .Y(n4940) );
  INVX1 U5282 ( .A(n3718), .Y(n2184) );
  INVX1 U5283 ( .A(n2159), .Y(n2160) );
  INVX1 U5284 ( .A(n2165), .Y(n2166) );
  INVX1 U5285 ( .A(n2163), .Y(n2164) );
  INVX1 U5286 ( .A(n2161), .Y(n2162) );
  INVX1 U5287 ( .A(n2170), .Y(n3592) );
  INVX1 U5288 ( .A(n1491), .Y(n1492) );
  INVX1 U5289 ( .A(n5059), .Y(n5058) );
  INVX1 U5290 ( .A(n5044), .Y(n5043) );
  INVX1 U5291 ( .A(n5056), .Y(n5055) );
  INVX1 U5292 ( .A(n5062), .Y(n5061) );
  INVX1 U5293 ( .A(n5053), .Y(n5052) );
  INVX1 U5294 ( .A(n5044), .Y(n5042) );
  INVX1 U5295 ( .A(n5056), .Y(n5054) );
  INVX1 U5296 ( .A(n5065), .Y(n5064) );
  INVX1 U5297 ( .A(n5062), .Y(n5060) );
  INVX1 U5298 ( .A(n5053), .Y(n5051) );
  INVX1 U5299 ( .A(n5065), .Y(n5063) );
  INVX1 U5300 ( .A(n5068), .Y(n5067) );
  INVX1 U5301 ( .A(n5068), .Y(n5066) );
  INVX1 U5302 ( .A(n124), .Y(n4927) );
  INVX1 U5303 ( .A(n3703), .Y(n2173) );
  INVX1 U5304 ( .A(n3707), .Y(n2185) );
  INVX1 U5305 ( .A(n28), .Y(n4962) );
  INVX1 U5306 ( .A(n3711), .Y(n2197) );
  INVX1 U5307 ( .A(n3709), .Y(n2191) );
  INVX1 U5308 ( .A(n3705), .Y(n2179) );
  INVX1 U5309 ( .A(n3704), .Y(n2176) );
  AND2X1 U5310 ( .A(n3696), .B(n3718), .Y(n2183) );
  AND2X1 U5311 ( .A(n3694), .B(n3716), .Y(n2177) );
  INVX1 U5312 ( .A(n36), .Y(n4958) );
  AND2X1 U5313 ( .A(n3700), .B(n3722), .Y(n2195) );
  AND2X1 U5314 ( .A(n3693), .B(n3715), .Y(n2174) );
  OR2X1 U5315 ( .A(n3720), .B(n3698), .Y(n4822) );
  OR2X1 U5316 ( .A(n3716), .B(n3694), .Y(n4823) );
  OR2X1 U5317 ( .A(n3722), .B(n3700), .Y(n4824) );
  OR2X1 U5318 ( .A(n3718), .B(n3696), .Y(n4825) );
  OR2X1 U5319 ( .A(n3715), .B(n3693), .Y(n4826) );
  INVX1 U5320 ( .A(b[30]), .Y(n5034) );
  INVX1 U5321 ( .A(b[27]), .Y(n5028) );
  INVX1 U5322 ( .A(b[28]), .Y(n5030) );
  INVX1 U5323 ( .A(b[29]), .Y(n5032) );
  INVX1 U5324 ( .A(b[23]), .Y(n5020) );
  INVX1 U5325 ( .A(n1792), .Y(n3190) );
  INVX1 U5326 ( .A(n2107), .Y(n3525) );
  INVX1 U5327 ( .A(n1918), .Y(n3324) );
  INVX1 U5328 ( .A(n1855), .Y(n3257) );
  INVX1 U5329 ( .A(n1729), .Y(n3123) );
  INVX1 U5330 ( .A(n1666), .Y(n3056) );
  INVX1 U5331 ( .A(n1603), .Y(n2989) );
  INVX1 U5332 ( .A(n58), .Y(n4946) );
  INVX1 U5333 ( .A(n3720), .Y(n2190) );
  INVX1 U5334 ( .A(n34), .Y(n4960) );
  INVX1 U5335 ( .A(n3722), .Y(n2196) );
  INVX1 U5336 ( .A(n118), .Y(n4930) );
  INVX1 U5337 ( .A(n3715), .Y(n2175) );
  INVX1 U5338 ( .A(n106), .Y(n4934) );
  INVX1 U5339 ( .A(n3716), .Y(n2178) );
  INVX1 U5340 ( .A(n4829), .Y(n4928) );
  XNOR2X1 U5341 ( .A(n3557), .B(n5038), .Y(n4827) );
  INVX1 U5342 ( .A(n4925), .Y(n4924) );
  INVX1 U5343 ( .A(n4990), .Y(n4989) );
  INVX1 U5344 ( .A(a[11]), .Y(n5050) );
  INVX1 U5345 ( .A(b[10]), .Y(n5000) );
  INVX1 U5346 ( .A(b[7]), .Y(n4994) );
  INVX1 U5347 ( .A(b[12]), .Y(n5004) );
  INVX1 U5348 ( .A(b[13]), .Y(n5006) );
  INVX1 U5349 ( .A(b[26]), .Y(n5026) );
  INVX1 U5350 ( .A(b[14]), .Y(n5008) );
  INVX1 U5351 ( .A(a[8]), .Y(n5047) );
  INVX1 U5352 ( .A(n5059), .Y(n5057) );
  OR2X1 U5353 ( .A(n2889), .B(n5039), .Y(n4828) );
  INVX1 U5354 ( .A(n508), .Y(n506) );
  INVX1 U5355 ( .A(n4609), .Y(n783) );
  INVX1 U5356 ( .A(a[2]), .Y(n5041) );
  INVX1 U5357 ( .A(n345), .Y(n343) );
  INVX1 U5358 ( .A(n3958), .Y(n326) );
  INVX1 U5359 ( .A(n5040), .Y(n5038) );
  INVX1 U5360 ( .A(a[2]), .Y(n5040) );
  AND2X1 U5361 ( .A(n3692), .B(n3703), .Y(n2171) );
  INVX1 U5362 ( .A(a[20]), .Y(n5059) );
  OR2X1 U5363 ( .A(n3692), .B(a[31]), .Y(n4829) );
  INVX1 U5364 ( .A(b[5]), .Y(n4990) );
  INVX1 U5365 ( .A(n4688), .Y(n420) );
  INVX1 U5366 ( .A(n127), .Y(n4925) );
  INVX1 U5367 ( .A(a[31]), .Y(n2172) );
  INVX1 U5368 ( .A(n419), .Y(n417) );
  INVX1 U5369 ( .A(n4621), .Y(n552) );
  INVX1 U5370 ( .A(a[5]), .Y(n5044) );
  INVX1 U5371 ( .A(a[14]), .Y(n5053) );
  INVX1 U5372 ( .A(a[29]), .Y(n5068) );
  INVX1 U5373 ( .A(a[26]), .Y(n5065) );
  INVX1 U5374 ( .A(a[17]), .Y(n5056) );
  INVX1 U5375 ( .A(a[23]), .Y(n5062) );
  INVX1 U5376 ( .A(n230), .Y(n421) );
  INVX1 U5377 ( .A(n569), .Y(n567) );
  INVX1 U5378 ( .A(n4670), .Y(n553) );
  INVX1 U5379 ( .A(n353), .Y(n351) );
  INVX1 U5380 ( .A(n4666), .Y(n399) );
  INVX1 U5381 ( .A(n305), .Y(n303) );
  INVX1 U5382 ( .A(n4730), .Y(n593) );
  INVX1 U5383 ( .A(n635), .Y(n634) );
  INVX1 U5384 ( .A(n4733), .Y(n605) );
  INVX1 U5385 ( .A(n4758), .Y(n472) );
  INVX1 U5386 ( .A(n371), .Y(n373) );
  INVX1 U5387 ( .A(n227), .Y(n4921) );
  INVX1 U5388 ( .A(n441), .Y(n439) );
  INVX1 U5389 ( .A(n4663), .Y(n456) );
  INVX1 U5390 ( .A(n4658), .Y(n350) );
  INVX1 U5391 ( .A(n4665), .Y(n492) );
  INVX1 U5392 ( .A(n4608), .Y(n316) );
  INVX1 U5393 ( .A(n4664), .Y(n327) );
  INVX1 U5394 ( .A(n4877), .Y(n480) );
  INVX1 U5395 ( .A(n4888), .Y(n379) );
  INVX1 U5396 ( .A(n4870), .Y(n788) );
  INVX1 U5397 ( .A(n4855), .Y(n639) );
  INVX1 U5398 ( .A(n395), .Y(n393) );
  INVX1 U5399 ( .A(n4889), .Y(n360) );
  INVX1 U5400 ( .A(n4893), .Y(n338) );
  INVX1 U5401 ( .A(n367), .Y(n365) );
  INVX1 U5402 ( .A(n4864), .Y(n791) );
  INVX1 U5403 ( .A(n4866), .Y(n790) );
  INVX1 U5404 ( .A(n4892), .Y(n764) );
  INVX1 U5405 ( .A(n4896), .Y(n762) );
  INVX1 U5406 ( .A(n4898), .Y(n761) );
  INVX1 U5407 ( .A(n4900), .Y(n760) );
  INVX1 U5408 ( .A(n4886), .Y(n403) );
  INVX1 U5409 ( .A(n4875), .Y(n496) );
  INVX1 U5410 ( .A(n4862), .Y(n597) );
  INVX1 U5411 ( .A(n4879), .Y(n460) );
  INVX1 U5412 ( .A(n4868), .Y(n789) );
  INVX1 U5413 ( .A(n4884), .Y(n770) );
  INVX1 U5414 ( .A(n4858), .Y(n624) );
  INVX1 U5415 ( .A(n4856), .Y(n631) );
  INVX1 U5416 ( .A(n4860), .Y(n612) );
  INVX1 U5417 ( .A(n4881), .Y(n434) );
  INVX1 U5418 ( .A(n4849), .Y(n652) );
  INVX1 U5419 ( .A(n4882), .Y(n771) );
  INVX1 U5420 ( .A(n4890), .Y(n765) );
  INVX1 U5421 ( .A(n4894), .Y(n763) );
  INVX1 U5422 ( .A(n4874), .Y(n778) );
  INVX1 U5423 ( .A(n4878), .Y(n465) );
  INVX1 U5424 ( .A(n4873), .Y(n501) );
  INVX1 U5425 ( .A(n4876), .Y(n485) );
  INVX1 U5426 ( .A(n4885), .Y(n412) );
  INVX1 U5427 ( .A(n4861), .Y(n602) );
  INVX1 U5428 ( .A(n4859), .Y(n617) );
  INVX1 U5429 ( .A(n4880), .Y(n447) );
  INVX1 U5430 ( .A(n4887), .Y(n388) );
  INVX1 U5431 ( .A(n4872), .Y(n786) );
  INVX1 U5432 ( .A(n3915), .Y(n800) );
  INVX1 U5433 ( .A(n4871), .Y(n562) );
  INVX1 U5434 ( .A(n4851), .Y(n649) );
  INVX1 U5435 ( .A(n4857), .Y(n797) );
  INVX1 U5436 ( .A(n4854), .Y(n799) );
  INVX1 U5437 ( .A(n4901), .Y(n298) );
  AOI22X1 U5438 ( .A(n4980), .B(b[1]), .C(n4), .D(n4981), .Y(n2169) );
  AOI22X1 U5439 ( .A(n4983), .B(n4980), .C(n4), .D(b[1]), .Y(n2167) );
  AOI22X1 U5440 ( .A(n4985), .B(n4980), .C(n4983), .D(n4), .Y(n2165) );
  AOI22X1 U5441 ( .A(n4987), .B(n4979), .C(n4985), .D(n4), .Y(n2163) );
  AOI22X1 U5442 ( .A(n4989), .B(n4980), .C(n4987), .D(n4), .Y(n2161) );
  AOI22X1 U5443 ( .A(n4991), .B(n4979), .C(n4989), .D(n4), .Y(n2159) );
  AOI22X1 U5444 ( .A(n4993), .B(n4979), .C(n4991), .D(n4), .Y(n2157) );
  AOI22X1 U5445 ( .A(n4995), .B(n4980), .C(n4993), .D(n4), .Y(n2155) );
  AOI22X1 U5446 ( .A(n4997), .B(n4980), .C(n4995), .D(n4), .Y(n2153) );
  AOI22X1 U5447 ( .A(n4999), .B(n4980), .C(n4997), .D(n4), .Y(n2151) );
  AOI22X1 U5448 ( .A(n5001), .B(n4980), .C(n4999), .D(n4), .Y(n2149) );
  AOI22X1 U5449 ( .A(n5003), .B(n4980), .C(n5001), .D(n4), .Y(n2147) );
  AOI22X1 U5450 ( .A(n5005), .B(n4980), .C(n5003), .D(n4), .Y(n2145) );
  AOI22X1 U5451 ( .A(n5007), .B(n4980), .C(n5005), .D(n4), .Y(n2143) );
  AOI22X1 U5452 ( .A(n5009), .B(n4980), .C(n5007), .D(n4), .Y(n2141) );
  AOI22X1 U5453 ( .A(n5011), .B(n4980), .C(n5009), .D(n4), .Y(n2139) );
  AOI22X1 U5454 ( .A(n5011), .B(n4), .C(b[17]), .D(n4979), .Y(n2137) );
  AOI22X1 U5455 ( .A(b[17]), .B(n4), .C(n5013), .D(n4980), .Y(n2135) );
  AOI22X1 U5456 ( .A(n5013), .B(n4), .C(n5015), .D(n4980), .Y(n2133) );
  AOI22X1 U5457 ( .A(n5015), .B(n4), .C(b[20]), .D(n4979), .Y(n2131) );
  AOI22X1 U5458 ( .A(b[20]), .B(n4), .C(n5017), .D(n4979), .Y(n2129) );
  AOI22X1 U5459 ( .A(n5017), .B(n4), .C(b[22]), .D(n4979), .Y(n2127) );
  AOI22X1 U5460 ( .A(b[22]), .B(n4), .C(n5019), .D(n4979), .Y(n2125) );
  AOI22X1 U5461 ( .A(n5019), .B(n4), .C(n5021), .D(n4979), .Y(n2123) );
  AOI22X1 U5462 ( .A(n5021), .B(n4), .C(n5023), .D(n4979), .Y(n2121) );
  AOI22X1 U5463 ( .A(n5023), .B(n4), .C(n5025), .D(n4979), .Y(n2119) );
  AOI22X1 U5464 ( .A(n5025), .B(n4), .C(n5027), .D(n4979), .Y(n2117) );
  AOI22X1 U5465 ( .A(n5027), .B(n4), .C(n5029), .D(n4979), .Y(n2115) );
  AOI22X1 U5466 ( .A(n5029), .B(n4), .C(n5031), .D(n4979), .Y(n2113) );
  AOI22X1 U5467 ( .A(n5031), .B(n4), .C(n5033), .D(n4979), .Y(n2111) );
  AOI22X1 U5468 ( .A(n5033), .B(n4), .C(n4980), .D(n5035), .Y(n2109) );
  AOI22X1 U5469 ( .A(n4972), .B(b[1]), .C(n16), .D(n4981), .Y(n2106) );
  AOI22X1 U5470 ( .A(n4972), .B(n4983), .C(n16), .D(b[1]), .Y(n2104) );
  AOI22X1 U5471 ( .A(n4972), .B(n4985), .C(n16), .D(n4983), .Y(n2102) );
  AOI22X1 U5472 ( .A(n4972), .B(n4987), .C(n16), .D(n4985), .Y(n2100) );
  AOI22X1 U5473 ( .A(n4972), .B(n4989), .C(n16), .D(n4987), .Y(n2098) );
  AOI22X1 U5474 ( .A(n4972), .B(n4991), .C(n16), .D(n4989), .Y(n2096) );
  AOI22X1 U5475 ( .A(n4972), .B(n4993), .C(n16), .D(n4991), .Y(n2094) );
  AOI22X1 U5476 ( .A(n4972), .B(n4995), .C(n16), .D(n4993), .Y(n2092) );
  AOI22X1 U5477 ( .A(n4972), .B(n4997), .C(n16), .D(n4995), .Y(n2090) );
  AOI22X1 U5478 ( .A(n4972), .B(n4999), .C(n16), .D(n4997), .Y(n2088) );
  AOI22X1 U5479 ( .A(n4972), .B(n5001), .C(n16), .D(n4999), .Y(n2086) );
  AOI22X1 U5480 ( .A(n4972), .B(n5003), .C(n16), .D(n5001), .Y(n2084) );
  AOI22X1 U5481 ( .A(n4972), .B(n5005), .C(n4970), .D(n5003), .Y(n2082) );
  AOI22X1 U5482 ( .A(n4973), .B(n5007), .C(n4970), .D(n5005), .Y(n2080) );
  AOI22X1 U5483 ( .A(n4973), .B(n5009), .C(n4970), .D(n5007), .Y(n2078) );
  AOI22X1 U5484 ( .A(n4973), .B(n5011), .C(n4970), .D(n5009), .Y(n2076) );
  AOI22X1 U5485 ( .A(n4973), .B(b[17]), .C(n4970), .D(n5011), .Y(n2074) );
  AOI22X1 U5486 ( .A(n4973), .B(n5013), .C(n4970), .D(b[17]), .Y(n2072) );
  AOI22X1 U5487 ( .A(n4973), .B(n5015), .C(n4970), .D(n5013), .Y(n2070) );
  AOI22X1 U5488 ( .A(n4973), .B(b[20]), .C(n4970), .D(n5015), .Y(n2068) );
  AOI22X1 U5489 ( .A(n4973), .B(n5017), .C(n4970), .D(b[20]), .Y(n2066) );
  AOI22X1 U5490 ( .A(n4973), .B(b[22]), .C(n4970), .D(n5017), .Y(n2064) );
  AOI22X1 U5491 ( .A(n4973), .B(n5019), .C(n4970), .D(b[22]), .Y(n2062) );
  AOI22X1 U5492 ( .A(n4973), .B(n5021), .C(n4970), .D(n5019), .Y(n2060) );
  AOI22X1 U5493 ( .A(n4973), .B(n5023), .C(n4970), .D(n5021), .Y(n2058) );
  AOI22X1 U5494 ( .A(n4973), .B(n5025), .C(n4970), .D(n5023), .Y(n2056) );
  AOI22X1 U5495 ( .A(n4973), .B(n5027), .C(n4970), .D(n5025), .Y(n2054) );
  AOI22X1 U5496 ( .A(n4972), .B(n5029), .C(n4970), .D(n5027), .Y(n2052) );
  AOI22X1 U5497 ( .A(n4973), .B(n5031), .C(n4970), .D(n5029), .Y(n2050) );
  AOI22X1 U5498 ( .A(n4972), .B(n5033), .C(n4970), .D(n5031), .Y(n2048) );
  AOI22X1 U5499 ( .A(n4973), .B(n5035), .C(n4970), .D(n5033), .Y(n2046) );
  AOI22X1 U5500 ( .A(n4964), .B(b[1]), .C(n28), .D(n4981), .Y(n2043) );
  AOI22X1 U5501 ( .A(n4963), .B(n4983), .C(n28), .D(b[1]), .Y(n2041) );
  AOI22X1 U5502 ( .A(n4963), .B(n4985), .C(n28), .D(n4983), .Y(n2039) );
  AOI22X1 U5503 ( .A(n4964), .B(n4987), .C(n28), .D(n4985), .Y(n2037) );
  AOI22X1 U5504 ( .A(n4963), .B(n4989), .C(n28), .D(n4987), .Y(n2035) );
  AOI22X1 U5505 ( .A(n4964), .B(n4991), .C(n28), .D(n4989), .Y(n2033) );
  AOI22X1 U5506 ( .A(n4963), .B(n4993), .C(n28), .D(n4991), .Y(n2031) );
  AOI22X1 U5507 ( .A(n4964), .B(n4995), .C(n28), .D(n4993), .Y(n2029) );
  AOI22X1 U5508 ( .A(n4964), .B(n4997), .C(n28), .D(n4995), .Y(n2027) );
  AOI22X1 U5509 ( .A(n4964), .B(n4999), .C(n28), .D(n4997), .Y(n2025) );
  AOI22X1 U5510 ( .A(n4964), .B(n5001), .C(n28), .D(n4999), .Y(n2023) );
  AOI22X1 U5511 ( .A(n4964), .B(n5003), .C(n28), .D(n5001), .Y(n2021) );
  AOI22X1 U5512 ( .A(n4964), .B(n5005), .C(n4961), .D(n5003), .Y(n2019) );
  AOI22X1 U5513 ( .A(n4964), .B(n5007), .C(n4961), .D(n5005), .Y(n2017) );
  AOI22X1 U5514 ( .A(n4964), .B(n5009), .C(n4961), .D(n5007), .Y(n2015) );
  AOI22X1 U5515 ( .A(n4964), .B(n5011), .C(n4961), .D(n5009), .Y(n2013) );
  AOI22X1 U5516 ( .A(n4961), .B(n5011), .C(n4964), .D(b[17]), .Y(n2011) );
  AOI22X1 U5517 ( .A(n4961), .B(b[17]), .C(n4964), .D(n5013), .Y(n2009) );
  AOI22X1 U5518 ( .A(n4961), .B(n5013), .C(n4964), .D(n5015), .Y(n2007) );
  AOI22X1 U5519 ( .A(n4961), .B(n5015), .C(n4963), .D(b[20]), .Y(n2005) );
  AOI22X1 U5520 ( .A(n4961), .B(b[20]), .C(n4963), .D(n5017), .Y(n2003) );
  AOI22X1 U5521 ( .A(n4961), .B(n5017), .C(n4963), .D(b[22]), .Y(n2001) );
  AOI22X1 U5522 ( .A(n4961), .B(b[22]), .C(n4963), .D(n5019), .Y(n1999) );
  AOI22X1 U5523 ( .A(n4961), .B(n5019), .C(n4963), .D(n5021), .Y(n1997) );
  AOI22X1 U5524 ( .A(n4961), .B(n5021), .C(n4963), .D(n5023), .Y(n1995) );
  AOI22X1 U5525 ( .A(n4961), .B(n5023), .C(n4963), .D(n5025), .Y(n1993) );
  AOI22X1 U5526 ( .A(n4961), .B(n5025), .C(n4963), .D(n5027), .Y(n1991) );
  AOI22X1 U5527 ( .A(n4961), .B(n5027), .C(n4963), .D(n5029), .Y(n1989) );
  AOI22X1 U5528 ( .A(n4961), .B(n5029), .C(n4963), .D(n5031), .Y(n1987) );
  AOI22X1 U5529 ( .A(n4961), .B(n5031), .C(n4963), .D(n5033), .Y(n1985) );
  AOI22X1 U5530 ( .A(n4961), .B(n5033), .C(n4963), .D(n5035), .Y(n1983) );
  AOI22X1 U5531 ( .A(n4955), .B(b[1]), .C(n4953), .D(n4981), .Y(n1980) );
  AOI22X1 U5532 ( .A(n4955), .B(n4983), .C(n4953), .D(b[1]), .Y(n1978) );
  AOI22X1 U5533 ( .A(n4955), .B(n4985), .C(n4953), .D(n4983), .Y(n1976) );
  AOI22X1 U5534 ( .A(n4955), .B(n4987), .C(n4953), .D(n4985), .Y(n1974) );
  AOI22X1 U5535 ( .A(n4955), .B(n4989), .C(n40), .D(n4987), .Y(n1972) );
  AOI22X1 U5536 ( .A(n4955), .B(n4991), .C(n40), .D(n4989), .Y(n1970) );
  AOI22X1 U5537 ( .A(n4955), .B(n4993), .C(n40), .D(n4991), .Y(n1968) );
  AOI22X1 U5538 ( .A(n4955), .B(n4995), .C(n40), .D(n4993), .Y(n1966) );
  AOI22X1 U5539 ( .A(n4955), .B(n4997), .C(n40), .D(n4995), .Y(n1964) );
  AOI22X1 U5540 ( .A(n4955), .B(n4999), .C(n40), .D(n4997), .Y(n1962) );
  AOI22X1 U5541 ( .A(n4955), .B(n5001), .C(n40), .D(n4999), .Y(n1960) );
  AOI22X1 U5542 ( .A(n4955), .B(n5003), .C(n40), .D(n5001), .Y(n1958) );
  AOI22X1 U5543 ( .A(n4955), .B(n5005), .C(n40), .D(n5003), .Y(n1956) );
  AOI22X1 U5544 ( .A(n4955), .B(n5007), .C(n40), .D(n5005), .Y(n1954) );
  AOI22X1 U5545 ( .A(n4955), .B(n5009), .C(n40), .D(n5007), .Y(n1952) );
  AOI22X1 U5546 ( .A(n4955), .B(n5011), .C(n40), .D(n5009), .Y(n1950) );
  AOI22X1 U5547 ( .A(n4953), .B(n5011), .C(n4955), .D(b[17]), .Y(n1948) );
  AOI22X1 U5548 ( .A(n4953), .B(b[17]), .C(n4955), .D(n5013), .Y(n1946) );
  AOI22X1 U5549 ( .A(n4953), .B(n5013), .C(n4955), .D(n5015), .Y(n1944) );
  AOI22X1 U5550 ( .A(n4953), .B(n5015), .C(n4955), .D(b[20]), .Y(n1942) );
  AOI22X1 U5551 ( .A(n4953), .B(b[20]), .C(n4955), .D(n5017), .Y(n1940) );
  AOI22X1 U5552 ( .A(n4953), .B(n5017), .C(n4955), .D(b[22]), .Y(n1938) );
  AOI22X1 U5553 ( .A(n4953), .B(b[22]), .C(n4955), .D(n5019), .Y(n1936) );
  AOI22X1 U5554 ( .A(n4953), .B(n5019), .C(n4955), .D(n5021), .Y(n1934) );
  AOI22X1 U5555 ( .A(n40), .B(n5021), .C(n4955), .D(n5023), .Y(n1932) );
  AOI22X1 U5556 ( .A(n40), .B(n5023), .C(n4955), .D(n5025), .Y(n1930) );
  AOI22X1 U5557 ( .A(n40), .B(n5025), .C(n4955), .D(n5027), .Y(n1928) );
  AOI22X1 U5558 ( .A(n40), .B(n5027), .C(n4955), .D(n5029), .Y(n1926) );
  AOI22X1 U5559 ( .A(n40), .B(n5029), .C(n4955), .D(n5031), .Y(n1924) );
  AOI22X1 U5560 ( .A(n40), .B(n5031), .C(n4955), .D(n5033), .Y(n1922) );
  AOI22X1 U5561 ( .A(n4953), .B(n5033), .C(n4955), .D(n5035), .Y(n1920) );
  AOI22X1 U5562 ( .A(n4948), .B(b[1]), .C(n52), .D(n4981), .Y(n1917) );
  AOI22X1 U5563 ( .A(n4948), .B(n4983), .C(n52), .D(b[1]), .Y(n1915) );
  AOI22X1 U5564 ( .A(n4948), .B(n4985), .C(n52), .D(n4983), .Y(n1913) );
  AOI22X1 U5565 ( .A(n4948), .B(n4987), .C(n52), .D(n4985), .Y(n1911) );
  AOI22X1 U5566 ( .A(n4948), .B(n4989), .C(n52), .D(n4987), .Y(n1909) );
  AOI22X1 U5567 ( .A(n4948), .B(n4991), .C(n52), .D(n4989), .Y(n1907) );
  AOI22X1 U5568 ( .A(n4947), .B(n4993), .C(n52), .D(n4991), .Y(n1905) );
  AOI22X1 U5569 ( .A(n4947), .B(n4995), .C(n52), .D(n4993), .Y(n1903) );
  AOI22X1 U5570 ( .A(n4947), .B(n4997), .C(n52), .D(n4995), .Y(n1901) );
  AOI22X1 U5571 ( .A(n4947), .B(n4999), .C(n52), .D(n4997), .Y(n1899) );
  AOI22X1 U5572 ( .A(n4947), .B(n5001), .C(n52), .D(n4999), .Y(n1897) );
  AOI22X1 U5573 ( .A(n4947), .B(n5003), .C(n52), .D(n5001), .Y(n1895) );
  AOI22X1 U5574 ( .A(n4947), .B(n5005), .C(n52), .D(n5003), .Y(n1893) );
  AOI22X1 U5575 ( .A(n4947), .B(n5007), .C(n52), .D(n5005), .Y(n1891) );
  AOI22X1 U5576 ( .A(n4947), .B(n5009), .C(n52), .D(n5007), .Y(n1889) );
  AOI22X1 U5577 ( .A(n4947), .B(n5011), .C(n52), .D(n5009), .Y(n1887) );
  AOI22X1 U5578 ( .A(n52), .B(n5011), .C(n4947), .D(b[17]), .Y(n1885) );
  AOI22X1 U5579 ( .A(n52), .B(b[17]), .C(n4947), .D(n5013), .Y(n1883) );
  AOI22X1 U5580 ( .A(n52), .B(n5013), .C(n4947), .D(n5015), .Y(n1881) );
  AOI22X1 U5581 ( .A(n52), .B(n5015), .C(n4947), .D(b[20]), .Y(n1879) );
  AOI22X1 U5582 ( .A(n52), .B(b[20]), .C(n4947), .D(n5017), .Y(n1877) );
  AOI22X1 U5583 ( .A(n52), .B(n5017), .C(n4947), .D(b[22]), .Y(n1875) );
  AOI22X1 U5584 ( .A(n52), .B(b[22]), .C(n4947), .D(n5019), .Y(n1873) );
  AOI22X1 U5585 ( .A(n52), .B(n5019), .C(n4947), .D(n5021), .Y(n1871) );
  AOI22X1 U5586 ( .A(n52), .B(n5021), .C(n4947), .D(n5023), .Y(n1869) );
  AOI22X1 U5587 ( .A(n52), .B(n5023), .C(n4947), .D(n5025), .Y(n1867) );
  AOI22X1 U5588 ( .A(n52), .B(n5025), .C(n4947), .D(n5027), .Y(n1865) );
  AOI22X1 U5589 ( .A(n52), .B(n5027), .C(n4947), .D(n5029), .Y(n1863) );
  AOI22X1 U5590 ( .A(n52), .B(n5029), .C(n4947), .D(n5031), .Y(n1861) );
  AOI22X1 U5591 ( .A(n52), .B(n5031), .C(n4947), .D(n5033), .Y(n1859) );
  AOI22X1 U5592 ( .A(n52), .B(n5033), .C(n4947), .D(n5035), .Y(n1857) );
  AOI22X1 U5593 ( .A(n4944), .B(b[1]), .C(n64), .D(n4981), .Y(n1854) );
  AOI22X1 U5594 ( .A(n4944), .B(n4983), .C(n64), .D(b[1]), .Y(n1852) );
  AOI22X1 U5595 ( .A(n4944), .B(n4985), .C(n64), .D(n4983), .Y(n1850) );
  AOI22X1 U5596 ( .A(n4944), .B(n4987), .C(n64), .D(n4985), .Y(n1848) );
  AOI22X1 U5597 ( .A(n4944), .B(n4989), .C(n64), .D(n4987), .Y(n1846) );
  AOI22X1 U5598 ( .A(n4944), .B(n4991), .C(n64), .D(n4989), .Y(n1844) );
  AOI22X1 U5599 ( .A(n4944), .B(n4993), .C(n64), .D(n4991), .Y(n1842) );
  AOI22X1 U5600 ( .A(n4944), .B(n4995), .C(n64), .D(n4993), .Y(n1840) );
  AOI22X1 U5601 ( .A(n4944), .B(n4997), .C(n64), .D(n4995), .Y(n1838) );
  AOI22X1 U5602 ( .A(n4944), .B(n4999), .C(n64), .D(n4997), .Y(n1836) );
  AOI22X1 U5603 ( .A(n4944), .B(n5001), .C(n64), .D(n4999), .Y(n1834) );
  AOI22X1 U5604 ( .A(n4944), .B(n5003), .C(n64), .D(n5001), .Y(n1832) );
  AOI22X1 U5605 ( .A(n4944), .B(n5005), .C(n64), .D(n5003), .Y(n1830) );
  AOI22X1 U5606 ( .A(n4944), .B(n5007), .C(n64), .D(n5005), .Y(n1828) );
  AOI22X1 U5607 ( .A(n4944), .B(n5009), .C(n64), .D(n5007), .Y(n1826) );
  AOI22X1 U5608 ( .A(n4944), .B(n5011), .C(n64), .D(n5009), .Y(n1824) );
  AOI22X1 U5609 ( .A(n64), .B(n5011), .C(n4944), .D(b[17]), .Y(n1822) );
  AOI22X1 U5610 ( .A(n64), .B(b[17]), .C(n4944), .D(n5013), .Y(n1820) );
  AOI22X1 U5611 ( .A(n64), .B(n5013), .C(n4944), .D(n5015), .Y(n1818) );
  AOI22X1 U5612 ( .A(n64), .B(n5015), .C(n4944), .D(b[20]), .Y(n1816) );
  AOI22X1 U5613 ( .A(n64), .B(b[20]), .C(n4944), .D(n5017), .Y(n1814) );
  AOI22X1 U5614 ( .A(n64), .B(n5017), .C(n4944), .D(b[22]), .Y(n1812) );
  AOI22X1 U5615 ( .A(n64), .B(b[22]), .C(n4944), .D(n5019), .Y(n1810) );
  AOI22X1 U5616 ( .A(n64), .B(n5019), .C(n4944), .D(n5021), .Y(n1808) );
  AOI22X1 U5617 ( .A(n64), .B(n5021), .C(n4944), .D(n5023), .Y(n1806) );
  AOI22X1 U5618 ( .A(n64), .B(n5023), .C(n4944), .D(n5025), .Y(n1804) );
  AOI22X1 U5619 ( .A(n64), .B(n5025), .C(n4944), .D(n5027), .Y(n1802) );
  AOI22X1 U5620 ( .A(n64), .B(n5027), .C(n4944), .D(n5029), .Y(n1800) );
  AOI22X1 U5621 ( .A(n64), .B(n5029), .C(n4944), .D(n5031), .Y(n1798) );
  AOI22X1 U5622 ( .A(n64), .B(n5031), .C(n4944), .D(n5033), .Y(n1796) );
  AOI22X1 U5623 ( .A(n64), .B(n5033), .C(n4944), .D(n5035), .Y(n1794) );
  AOI22X1 U5624 ( .A(n4941), .B(b[1]), .C(n76), .D(n4981), .Y(n1791) );
  AOI22X1 U5625 ( .A(n4941), .B(n4983), .C(n76), .D(b[1]), .Y(n1789) );
  AOI22X1 U5626 ( .A(n4941), .B(n4985), .C(n76), .D(n4983), .Y(n1787) );
  AOI22X1 U5627 ( .A(n4941), .B(n4987), .C(n76), .D(n4985), .Y(n1785) );
  AOI22X1 U5628 ( .A(n4941), .B(n4989), .C(n76), .D(n4987), .Y(n1783) );
  AOI22X1 U5629 ( .A(n4941), .B(n4991), .C(n76), .D(n4989), .Y(n1781) );
  AOI22X1 U5630 ( .A(n4941), .B(n4993), .C(n76), .D(n4991), .Y(n1779) );
  AOI22X1 U5631 ( .A(n4941), .B(n4995), .C(n76), .D(n4993), .Y(n1777) );
  AOI22X1 U5632 ( .A(n4941), .B(n4997), .C(n76), .D(n4995), .Y(n1775) );
  AOI22X1 U5633 ( .A(n4941), .B(n4999), .C(n76), .D(n4997), .Y(n1773) );
  AOI22X1 U5634 ( .A(n4941), .B(n5001), .C(n76), .D(n4999), .Y(n1771) );
  AOI22X1 U5635 ( .A(n4941), .B(n5003), .C(n76), .D(n5001), .Y(n1769) );
  AOI22X1 U5636 ( .A(n4941), .B(n5005), .C(n76), .D(n5003), .Y(n1767) );
  AOI22X1 U5637 ( .A(n4941), .B(n5007), .C(n76), .D(n5005), .Y(n1765) );
  AOI22X1 U5638 ( .A(n4941), .B(n5009), .C(n76), .D(n5007), .Y(n1763) );
  AOI22X1 U5639 ( .A(n4941), .B(n5011), .C(n76), .D(n5009), .Y(n1761) );
  AOI22X1 U5640 ( .A(n76), .B(n5011), .C(n4941), .D(b[17]), .Y(n1759) );
  AOI22X1 U5641 ( .A(n76), .B(b[17]), .C(n4941), .D(n5013), .Y(n1757) );
  AOI22X1 U5642 ( .A(n76), .B(n5013), .C(n4941), .D(n5015), .Y(n1755) );
  AOI22X1 U5643 ( .A(n76), .B(n5015), .C(n4941), .D(b[20]), .Y(n1753) );
  AOI22X1 U5644 ( .A(n76), .B(b[20]), .C(n4941), .D(n5017), .Y(n1751) );
  AOI22X1 U5645 ( .A(n76), .B(n5017), .C(n4941), .D(b[22]), .Y(n1749) );
  AOI22X1 U5646 ( .A(n76), .B(b[22]), .C(n4941), .D(n5019), .Y(n1747) );
  AOI22X1 U5647 ( .A(n76), .B(n5019), .C(n4941), .D(n5021), .Y(n1745) );
  AOI22X1 U5648 ( .A(n76), .B(n5021), .C(n4941), .D(n5023), .Y(n1743) );
  AOI22X1 U5649 ( .A(n76), .B(n5023), .C(n4941), .D(n5025), .Y(n1741) );
  AOI22X1 U5650 ( .A(n76), .B(n5025), .C(n4941), .D(n5027), .Y(n1739) );
  AOI22X1 U5651 ( .A(n76), .B(n5027), .C(n4941), .D(n5029), .Y(n1737) );
  AOI22X1 U5652 ( .A(n76), .B(n5029), .C(n4941), .D(n5031), .Y(n1735) );
  AOI22X1 U5653 ( .A(n76), .B(n5031), .C(n4941), .D(n5033), .Y(n1733) );
  AOI22X1 U5654 ( .A(n76), .B(n5033), .C(n4941), .D(n5035), .Y(n1731) );
  AOI22X1 U5655 ( .A(n4938), .B(b[1]), .C(n88), .D(n4981), .Y(n1728) );
  AOI22X1 U5656 ( .A(n4938), .B(n4983), .C(n88), .D(b[1]), .Y(n1726) );
  AOI22X1 U5657 ( .A(n4938), .B(n4985), .C(n88), .D(n4983), .Y(n1724) );
  AOI22X1 U5658 ( .A(n4938), .B(n4987), .C(n88), .D(n4985), .Y(n1722) );
  AOI22X1 U5659 ( .A(n4938), .B(n4989), .C(n88), .D(n4987), .Y(n1720) );
  AOI22X1 U5660 ( .A(n4938), .B(n4991), .C(n88), .D(n4989), .Y(n1718) );
  AOI22X1 U5661 ( .A(n4938), .B(n4993), .C(n88), .D(n4991), .Y(n1716) );
  AOI22X1 U5662 ( .A(n4938), .B(n4995), .C(n88), .D(n4993), .Y(n1714) );
  AOI22X1 U5663 ( .A(n4938), .B(n4997), .C(n88), .D(n4995), .Y(n1712) );
  AOI22X1 U5664 ( .A(n4938), .B(n4999), .C(n88), .D(n4997), .Y(n1710) );
  AOI22X1 U5665 ( .A(n4938), .B(n5001), .C(n88), .D(n4999), .Y(n1708) );
  AOI22X1 U5666 ( .A(n4938), .B(n5003), .C(n88), .D(n5001), .Y(n1706) );
  AOI22X1 U5667 ( .A(n4938), .B(n5005), .C(n88), .D(n5003), .Y(n1704) );
  AOI22X1 U5668 ( .A(n4938), .B(n5007), .C(n88), .D(n5005), .Y(n1702) );
  AOI22X1 U5669 ( .A(n4938), .B(n5009), .C(n88), .D(n5007), .Y(n1700) );
  AOI22X1 U5670 ( .A(n4938), .B(n5011), .C(n88), .D(n5009), .Y(n1698) );
  AOI22X1 U5671 ( .A(n88), .B(n5011), .C(n4938), .D(b[17]), .Y(n1696) );
  AOI22X1 U5672 ( .A(n88), .B(b[17]), .C(n4938), .D(n5013), .Y(n1694) );
  AOI22X1 U5673 ( .A(n88), .B(n5013), .C(n4938), .D(n5015), .Y(n1692) );
  AOI22X1 U5674 ( .A(n88), .B(n5015), .C(n4938), .D(b[20]), .Y(n1690) );
  AOI22X1 U5675 ( .A(n88), .B(b[20]), .C(n4938), .D(n5017), .Y(n1688) );
  AOI22X1 U5676 ( .A(n88), .B(n5017), .C(n4938), .D(b[22]), .Y(n1686) );
  AOI22X1 U5677 ( .A(n88), .B(b[22]), .C(n4938), .D(n5019), .Y(n1684) );
  AOI22X1 U5678 ( .A(n88), .B(n5019), .C(n4938), .D(n5021), .Y(n1682) );
  AOI22X1 U5679 ( .A(n88), .B(n5021), .C(n4938), .D(n5023), .Y(n1680) );
  AOI22X1 U5680 ( .A(n88), .B(n5023), .C(n4938), .D(n5025), .Y(n1678) );
  AOI22X1 U5681 ( .A(n88), .B(n5025), .C(n4938), .D(n5027), .Y(n1676) );
  AOI22X1 U5682 ( .A(n88), .B(n5027), .C(n4938), .D(n5029), .Y(n1674) );
  AOI22X1 U5683 ( .A(n88), .B(n5029), .C(n4938), .D(n5031), .Y(n1672) );
  AOI22X1 U5684 ( .A(n88), .B(n5031), .C(n4938), .D(n5033), .Y(n1670) );
  AOI22X1 U5685 ( .A(n88), .B(n5033), .C(n4938), .D(n5035), .Y(n1668) );
  AOI22X1 U5686 ( .A(n4935), .B(b[1]), .C(n100), .D(n4981), .Y(n1665) );
  AOI22X1 U5687 ( .A(n4935), .B(n4983), .C(n100), .D(b[1]), .Y(n1663) );
  AOI22X1 U5688 ( .A(n4935), .B(n4985), .C(n100), .D(n4983), .Y(n1661) );
  AOI22X1 U5689 ( .A(n4935), .B(n4987), .C(n100), .D(n4985), .Y(n1659) );
  AOI22X1 U5690 ( .A(n4935), .B(n4989), .C(n100), .D(n4987), .Y(n1657) );
  AOI22X1 U5691 ( .A(n4935), .B(n4991), .C(n100), .D(n4989), .Y(n1655) );
  AOI22X1 U5692 ( .A(n4935), .B(n4993), .C(n100), .D(n4991), .Y(n1653) );
  AOI22X1 U5693 ( .A(n4935), .B(n4995), .C(n100), .D(n4993), .Y(n1651) );
  AOI22X1 U5694 ( .A(n4935), .B(n4997), .C(n100), .D(n4995), .Y(n1649) );
  AOI22X1 U5695 ( .A(n4935), .B(n4999), .C(n100), .D(n4997), .Y(n1647) );
  AOI22X1 U5696 ( .A(n4935), .B(n5001), .C(n100), .D(n4999), .Y(n1645) );
  AOI22X1 U5697 ( .A(n4935), .B(n5003), .C(n100), .D(n5001), .Y(n1643) );
  AOI22X1 U5698 ( .A(n4935), .B(n5005), .C(n100), .D(n5003), .Y(n1641) );
  AOI22X1 U5699 ( .A(n4935), .B(n5007), .C(n100), .D(n5005), .Y(n1639) );
  AOI22X1 U5700 ( .A(n4935), .B(n5009), .C(n100), .D(n5007), .Y(n1637) );
  AOI22X1 U5701 ( .A(n4935), .B(n5011), .C(n100), .D(n5009), .Y(n1635) );
  AOI22X1 U5702 ( .A(n4935), .B(b[17]), .C(n100), .D(n5011), .Y(n1633) );
  AOI22X1 U5703 ( .A(n4935), .B(n5013), .C(n100), .D(b[17]), .Y(n1631) );
  AOI22X1 U5704 ( .A(n4935), .B(n5015), .C(n100), .D(n5013), .Y(n1629) );
  AOI22X1 U5705 ( .A(n4935), .B(b[20]), .C(n100), .D(n5015), .Y(n1627) );
  AOI22X1 U5706 ( .A(n4935), .B(n5017), .C(n100), .D(b[20]), .Y(n1625) );
  AOI22X1 U5707 ( .A(n4935), .B(b[22]), .C(n100), .D(n5017), .Y(n1623) );
  AOI22X1 U5708 ( .A(n4935), .B(n5019), .C(n100), .D(b[22]), .Y(n1621) );
  AOI22X1 U5709 ( .A(n4935), .B(n5021), .C(n100), .D(n5019), .Y(n1619) );
  AOI22X1 U5710 ( .A(n4935), .B(n5023), .C(n100), .D(n5021), .Y(n1617) );
  AOI22X1 U5711 ( .A(n4935), .B(n5025), .C(n100), .D(n5023), .Y(n1615) );
  AOI22X1 U5712 ( .A(n4935), .B(n5027), .C(n100), .D(n5025), .Y(n1613) );
  AOI22X1 U5713 ( .A(n4935), .B(n5029), .C(n100), .D(n5027), .Y(n1611) );
  AOI22X1 U5714 ( .A(n4935), .B(n5031), .C(n100), .D(n5029), .Y(n1609) );
  AOI22X1 U5715 ( .A(n4935), .B(n5033), .C(n100), .D(n5031), .Y(n1607) );
  AOI22X1 U5716 ( .A(n4935), .B(n5035), .C(n100), .D(n5033), .Y(n1605) );
  AOI22X1 U5717 ( .A(n4931), .B(b[1]), .C(n112), .D(n4981), .Y(n1602) );
  AOI22X1 U5718 ( .A(n4931), .B(n4983), .C(n112), .D(b[1]), .Y(n1600) );
  AOI22X1 U5719 ( .A(n4931), .B(n4985), .C(n112), .D(n4983), .Y(n1598) );
  AOI22X1 U5720 ( .A(n4931), .B(n4987), .C(n112), .D(n4985), .Y(n1596) );
  AOI22X1 U5721 ( .A(n4931), .B(n4989), .C(n112), .D(n4987), .Y(n1594) );
  AOI22X1 U5722 ( .A(n4931), .B(n4991), .C(n112), .D(n4989), .Y(n1592) );
  AOI22X1 U5723 ( .A(n4931), .B(n4993), .C(n112), .D(n4991), .Y(n1590) );
  AOI22X1 U5724 ( .A(n4931), .B(n4995), .C(n112), .D(n4993), .Y(n1588) );
  AOI22X1 U5725 ( .A(n4931), .B(n4997), .C(n112), .D(n4995), .Y(n1586) );
  AOI22X1 U5726 ( .A(n4931), .B(n4999), .C(n112), .D(n4997), .Y(n1584) );
  AOI22X1 U5727 ( .A(n4931), .B(n5001), .C(n112), .D(n4999), .Y(n1582) );
  AOI22X1 U5728 ( .A(n4931), .B(n5003), .C(n112), .D(n5001), .Y(n1580) );
  AOI22X1 U5729 ( .A(n4931), .B(n5005), .C(n112), .D(n5003), .Y(n1578) );
  AOI22X1 U5730 ( .A(n4932), .B(n5007), .C(n112), .D(n5005), .Y(n1576) );
  AOI22X1 U5731 ( .A(n4932), .B(n5009), .C(n112), .D(n5007), .Y(n1574) );
  AOI22X1 U5732 ( .A(n4932), .B(n5011), .C(n112), .D(n5009), .Y(n1572) );
  AOI22X1 U5733 ( .A(n4932), .B(b[17]), .C(n112), .D(n5011), .Y(n1570) );
  AOI22X1 U5734 ( .A(n4932), .B(n5013), .C(n112), .D(b[17]), .Y(n1568) );
  AOI22X1 U5735 ( .A(n4932), .B(n5015), .C(n112), .D(n5013), .Y(n1566) );
  AOI22X1 U5736 ( .A(n4932), .B(b[20]), .C(n112), .D(n5015), .Y(n1564) );
  AOI22X1 U5737 ( .A(n4932), .B(n5017), .C(n112), .D(b[20]), .Y(n1562) );
  AOI22X1 U5738 ( .A(n4932), .B(b[22]), .C(n112), .D(n5017), .Y(n1560) );
  AOI22X1 U5739 ( .A(n4932), .B(n5019), .C(n112), .D(b[22]), .Y(n1558) );
  AOI22X1 U5740 ( .A(n4932), .B(n5021), .C(n112), .D(n5019), .Y(n1556) );
  AOI22X1 U5741 ( .A(n4932), .B(n5023), .C(n112), .D(n5021), .Y(n1554) );
  AOI22X1 U5742 ( .A(n4932), .B(n5025), .C(n112), .D(n5023), .Y(n1552) );
  AOI22X1 U5743 ( .A(n4931), .B(n5027), .C(n112), .D(n5025), .Y(n1550) );
  AOI22X1 U5744 ( .A(n4932), .B(n5029), .C(n112), .D(n5027), .Y(n1548) );
  AOI22X1 U5745 ( .A(n4932), .B(n5031), .C(n112), .D(n5029), .Y(n1546) );
  AOI22X1 U5746 ( .A(n4932), .B(n5033), .C(n112), .D(n5031), .Y(n1544) );
  AOI22X1 U5747 ( .A(n4931), .B(n5035), .C(n112), .D(n5033), .Y(n1542) );
  AOI22X1 U5748 ( .A(n4928), .B(b[1]), .C(n4926), .D(n4981), .Y(n1539) );
  AOI22X1 U5749 ( .A(n4928), .B(b[2]), .C(n4926), .D(b[1]), .Y(n1537) );
  AOI22X1 U5750 ( .A(n4928), .B(n4985), .C(n4926), .D(n4983), .Y(n1535) );
  AOI22X1 U5751 ( .A(n4928), .B(n4987), .C(n4926), .D(n4985), .Y(n1533) );
  AOI22X1 U5752 ( .A(n4928), .B(n4989), .C(n4926), .D(n4987), .Y(n1531) );
  AOI22X1 U5753 ( .A(n4928), .B(n4991), .C(n4926), .D(n4989), .Y(n1529) );
  AOI22X1 U5754 ( .A(n4928), .B(n4993), .C(n4926), .D(n4991), .Y(n1527) );
  AOI22X1 U5755 ( .A(n4928), .B(n4995), .C(n4926), .D(n4993), .Y(n1525) );
  AOI22X1 U5756 ( .A(n4928), .B(n4997), .C(n4926), .D(n4995), .Y(n1523) );
  AOI22X1 U5757 ( .A(n4928), .B(n4999), .C(n4926), .D(n4997), .Y(n1521) );
  AOI22X1 U5758 ( .A(n4928), .B(n5001), .C(n4926), .D(n4999), .Y(n1519) );
  AOI22X1 U5759 ( .A(n4928), .B(n5003), .C(n4926), .D(n5001), .Y(n1517) );
  AOI22X1 U5760 ( .A(n4928), .B(n5005), .C(n124), .D(n5003), .Y(n1515) );
  AOI22X1 U5761 ( .A(n4928), .B(n5007), .C(n124), .D(n5005), .Y(n1513) );
  AOI22X1 U5762 ( .A(n4928), .B(n5009), .C(n124), .D(n5007), .Y(n1511) );
  AOI22X1 U5763 ( .A(n4928), .B(n5011), .C(n124), .D(n5009), .Y(n1509) );
  AOI22X1 U5764 ( .A(n4928), .B(b[17]), .C(n124), .D(n5011), .Y(n1507) );
  AOI22X1 U5765 ( .A(n4928), .B(n5013), .C(n124), .D(b[17]), .Y(n1505) );
  AOI22X1 U5766 ( .A(n4928), .B(n5015), .C(n124), .D(n5013), .Y(n1503) );
  AOI22X1 U5767 ( .A(n4928), .B(b[20]), .C(n124), .D(n5015), .Y(n1501) );
  AOI22X1 U5768 ( .A(n4928), .B(n5017), .C(n124), .D(b[20]), .Y(n1499) );
  AOI22X1 U5769 ( .A(n4928), .B(b[22]), .C(n124), .D(n5017), .Y(n1497) );
  AOI22X1 U5770 ( .A(n4928), .B(n5019), .C(n124), .D(b[22]), .Y(n1495) );
  AOI22X1 U5771 ( .A(n4928), .B(n5021), .C(n124), .D(n5019), .Y(n1493) );
  AOI22X1 U5772 ( .A(n4928), .B(n5023), .C(n124), .D(n5021), .Y(n1491) );
  AOI22X1 U5773 ( .A(n4928), .B(n5025), .C(n124), .D(n5023), .Y(n1489) );
  AOI22X1 U5774 ( .A(n4928), .B(n5027), .C(n124), .D(n5025), .Y(n1487) );
  AOI22X1 U5775 ( .A(n4928), .B(n5029), .C(n124), .D(n5027), .Y(n1485) );
  AOI22X1 U5776 ( .A(n4928), .B(n5031), .C(n124), .D(n5029), .Y(n1483) );
  AOI22X1 U5777 ( .A(n4928), .B(n5033), .C(n124), .D(n5031), .Y(n1481) );
  AOI22X1 U5778 ( .A(n4928), .B(n5035), .C(n124), .D(n5033), .Y(n1479) );
endmodule


module alu_DW02_mult_2_stage_0 ( A, B, TC, CLK, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC, CLK;
  wire   n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2;

  alu_DW_mult_tc_1 mult_96 ( .a({1'b0, A}), .b({1'b0, B}), .product({
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, PRODUCT[63:20], n26, 
        n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, 
        n41, n42, n43, n44, n45}), .ALU1ALU_MUL32_CLK(CLK) );
  DFFPOSX1 clk_r_REG89_S1 ( .D(n26), .CLK(CLK), .Q(PRODUCT[19]) );
  DFFPOSX1 clk_r_REG91_S1 ( .D(n27), .CLK(CLK), .Q(PRODUCT[18]) );
  DFFPOSX1 clk_r_REG92_S1 ( .D(n28), .CLK(CLK), .Q(PRODUCT[17]) );
  DFFPOSX1 clk_r_REG93_S1 ( .D(n29), .CLK(CLK), .Q(PRODUCT[16]) );
  DFFPOSX1 clk_r_REG94_S1 ( .D(n30), .CLK(CLK), .Q(PRODUCT[15]) );
  DFFPOSX1 clk_r_REG95_S1 ( .D(n31), .CLK(CLK), .Q(PRODUCT[14]) );
  DFFPOSX1 clk_r_REG96_S1 ( .D(n32), .CLK(CLK), .Q(PRODUCT[13]) );
  DFFPOSX1 clk_r_REG97_S1 ( .D(n33), .CLK(CLK), .Q(PRODUCT[12]) );
  DFFPOSX1 clk_r_REG98_S1 ( .D(n34), .CLK(CLK), .Q(PRODUCT[11]) );
  DFFPOSX1 clk_r_REG99_S1 ( .D(n35), .CLK(CLK), .Q(PRODUCT[10]) );
  DFFPOSX1 clk_r_REG100_S1 ( .D(n36), .CLK(CLK), .Q(PRODUCT[9]) );
  DFFPOSX1 clk_r_REG101_S1 ( .D(n37), .CLK(CLK), .Q(PRODUCT[8]) );
  DFFPOSX1 clk_r_REG102_S1 ( .D(n38), .CLK(CLK), .Q(PRODUCT[7]) );
  DFFPOSX1 clk_r_REG103_S1 ( .D(n39), .CLK(CLK), .Q(PRODUCT[6]) );
  DFFPOSX1 clk_r_REG104_S1 ( .D(n40), .CLK(CLK), .Q(PRODUCT[5]) );
  DFFPOSX1 clk_r_REG105_S1 ( .D(n41), .CLK(CLK), .Q(PRODUCT[4]) );
  DFFPOSX1 clk_r_REG106_S1 ( .D(n42), .CLK(CLK), .Q(PRODUCT[3]) );
  DFFPOSX1 clk_r_REG107_S1 ( .D(n43), .CLK(CLK), .Q(PRODUCT[2]) );
  DFFPOSX1 clk_r_REG108_S1 ( .D(n44), .CLK(CLK), .Q(PRODUCT[1]) );
  DFFPOSX1 clk_r_REG109_S1 ( .D(n45), .CLK(CLK), .Q(PRODUCT[0]) );
endmodule


module alu_DW_rightsh_0 ( A, DATA_TC, SH, B );
  input [63:0] A;
  input [4:0] SH;
  output [63:0] B;
  input DATA_TC;
  wire   n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076;

  INVX2 U659 ( .A(SH[0]), .Y(n735) );
  INVX1 U660 ( .A(n860), .Y(n801) );
  INVX1 U661 ( .A(n1042), .Y(n805) );
  INVX1 U662 ( .A(n1005), .Y(n810) );
  INVX1 U663 ( .A(n1003), .Y(n806) );
  INVX1 U664 ( .A(n1073), .Y(n797) );
  INVX1 U665 ( .A(n982), .Y(n798) );
  INVX1 U666 ( .A(n788), .Y(B[63]) );
  INVX1 U667 ( .A(n1055), .Y(n815) );
  INVX1 U668 ( .A(A[59]), .Y(n783) );
  INVX1 U669 ( .A(n1062), .Y(n803) );
  INVX1 U670 ( .A(A[62]), .Y(n786) );
  INVX1 U671 ( .A(n1029), .Y(n816) );
  INVX1 U672 ( .A(n887), .Y(n792) );
  INVX1 U673 ( .A(n931), .Y(n791) );
  INVX1 U674 ( .A(n844), .Y(n802) );
  INVX1 U675 ( .A(n1056), .Y(n811) );
  INVX1 U676 ( .A(n1027), .Y(n814) );
  INVX1 U677 ( .A(A[54]), .Y(n778) );
  INVX1 U678 ( .A(n747), .Y(n746) );
  INVX1 U679 ( .A(n747), .Y(n744) );
  INVX1 U680 ( .A(n747), .Y(n743) );
  INVX1 U681 ( .A(n747), .Y(n745) );
  INVX1 U682 ( .A(n735), .Y(n734) );
  INVX1 U683 ( .A(n735), .Y(n731) );
  INVX1 U684 ( .A(n735), .Y(n732) );
  INVX1 U685 ( .A(n735), .Y(n733) );
  INVX1 U686 ( .A(A[53]), .Y(n777) );
  INVX1 U687 ( .A(A[63]), .Y(n788) );
  INVX1 U688 ( .A(n1072), .Y(n809) );
  INVX1 U689 ( .A(n884), .Y(n796) );
  INVX1 U690 ( .A(n1065), .Y(n799) );
  INVX1 U691 ( .A(n1048), .Y(n812) );
  INVX1 U692 ( .A(n1071), .Y(n813) );
  INVX1 U693 ( .A(n1059), .Y(n807) );
  INVX1 U694 ( .A(n1050), .Y(n804) );
  INVX1 U695 ( .A(n1051), .Y(n800) );
  INVX1 U696 ( .A(n928), .Y(n795) );
  INVX1 U697 ( .A(n1049), .Y(n808) );
  INVX1 U698 ( .A(A[38]), .Y(n762) );
  INVX1 U699 ( .A(A[40]), .Y(n764) );
  INVX1 U700 ( .A(A[46]), .Y(n770) );
  INVX1 U701 ( .A(A[42]), .Y(n766) );
  INVX1 U702 ( .A(n1069), .Y(n819) );
  INVX1 U703 ( .A(A[44]), .Y(n768) );
  INVX1 U704 ( .A(A[60]), .Y(n784) );
  INVX1 U705 ( .A(n842), .Y(n794) );
  INVX1 U706 ( .A(n1074), .Y(n789) );
  INVX1 U707 ( .A(n858), .Y(n793) );
  INVX1 U708 ( .A(A[48]), .Y(n772) );
  INVX1 U709 ( .A(n753), .Y(n750) );
  INVX1 U710 ( .A(n753), .Y(n749) );
  INVX1 U711 ( .A(n753), .Y(n748) );
  INVX1 U712 ( .A(n753), .Y(n751) );
  INVX1 U713 ( .A(n753), .Y(n752) );
  INVX1 U714 ( .A(n742), .Y(n736) );
  INVX1 U715 ( .A(n741), .Y(n739) );
  INVX1 U716 ( .A(n742), .Y(n738) );
  INVX1 U717 ( .A(n742), .Y(n737) );
  INVX1 U718 ( .A(n741), .Y(n740) );
  INVX1 U719 ( .A(SH[2]), .Y(n747) );
  INVX1 U720 ( .A(n1044), .Y(n824) );
  INVX1 U721 ( .A(n1053), .Y(n823) );
  INVX1 U722 ( .A(n1045), .Y(n822) );
  INVX1 U723 ( .A(n1046), .Y(n820) );
  INVX1 U724 ( .A(n1054), .Y(n821) );
  INVX1 U725 ( .A(n1047), .Y(n818) );
  INVX1 U726 ( .A(n1070), .Y(n817) );
  INVX1 U727 ( .A(A[36]), .Y(n760) );
  INVX1 U728 ( .A(A[58]), .Y(n782) );
  INVX1 U729 ( .A(A[47]), .Y(n771) );
  INVX1 U730 ( .A(A[45]), .Y(n769) );
  INVX1 U731 ( .A(A[57]), .Y(n781) );
  INVX1 U732 ( .A(n985), .Y(n790) );
  INVX1 U733 ( .A(A[41]), .Y(n765) );
  INVX1 U734 ( .A(A[50]), .Y(n774) );
  INVX1 U735 ( .A(A[39]), .Y(n763) );
  INVX1 U736 ( .A(A[55]), .Y(n779) );
  INVX1 U737 ( .A(A[43]), .Y(n767) );
  INVX1 U738 ( .A(A[56]), .Y(n780) );
  INVX1 U739 ( .A(A[52]), .Y(n776) );
  INVX1 U740 ( .A(SH[3]), .Y(n753) );
  INVX1 U741 ( .A(SH[1]), .Y(n742) );
  INVX1 U742 ( .A(SH[1]), .Y(n741) );
  INVX1 U743 ( .A(n759), .Y(n754) );
  INVX1 U744 ( .A(n759), .Y(n758) );
  INVX1 U745 ( .A(n759), .Y(n756) );
  INVX1 U746 ( .A(n759), .Y(n755) );
  INVX1 U747 ( .A(n759), .Y(n757) );
  INVX1 U748 ( .A(A[61]), .Y(n785) );
  INVX1 U749 ( .A(A[49]), .Y(n773) );
  INVX1 U750 ( .A(SH[4]), .Y(n759) );
  INVX1 U751 ( .A(A[37]), .Y(n761) );
  INVX1 U752 ( .A(A[51]), .Y(n775) );
  MUX2X1 U753 ( .B(n825), .A(n826), .S(n755), .Y(B[9]) );
  MUX2X1 U754 ( .B(n798), .A(n806), .S(n749), .Y(n825) );
  MUX2X1 U755 ( .B(n827), .A(n828), .S(n755), .Y(B[8]) );
  MUX2X1 U756 ( .B(n797), .A(n829), .S(n750), .Y(n827) );
  MUX2X1 U757 ( .B(n830), .A(n831), .S(n756), .Y(B[7]) );
  MUX2X1 U758 ( .B(n832), .A(n833), .S(n750), .Y(n830) );
  MUX2X1 U759 ( .B(n796), .A(n800), .S(n743), .Y(n832) );
  MUX2X1 U760 ( .B(n834), .A(n835), .S(n758), .Y(B[6]) );
  MUX2X1 U761 ( .B(n836), .A(n837), .S(n752), .Y(n834) );
  MUX2X1 U762 ( .B(n795), .A(n799), .S(n743), .Y(n836) );
  MUX2X1 U763 ( .B(n838), .A(n788), .S(n758), .Y(B[62]) );
  MUX2X1 U764 ( .B(n839), .A(n788), .S(n758), .Y(B[61]) );
  MUX2X1 U765 ( .B(n840), .A(n788), .S(n758), .Y(B[60]) );
  MUX2X1 U766 ( .B(n794), .A(n841), .S(n758), .Y(B[5]) );
  MUX2X1 U767 ( .B(n843), .A(n844), .S(n752), .Y(n842) );
  MUX2X1 U768 ( .B(n845), .A(n846), .S(n744), .Y(n843) );
  MUX2X1 U769 ( .B(n847), .A(n788), .S(n758), .Y(B[59]) );
  MUX2X1 U770 ( .B(n848), .A(n788), .S(n758), .Y(B[58]) );
  MUX2X1 U771 ( .B(n849), .A(n788), .S(n758), .Y(B[57]) );
  MUX2X1 U772 ( .B(n850), .A(n788), .S(n758), .Y(B[56]) );
  MUX2X1 U773 ( .B(n851), .A(n788), .S(n758), .Y(B[55]) );
  MUX2X1 U774 ( .B(n852), .A(n788), .S(n758), .Y(B[54]) );
  MUX2X1 U775 ( .B(n853), .A(n788), .S(n758), .Y(B[53]) );
  MUX2X1 U776 ( .B(n854), .A(n788), .S(n757), .Y(B[52]) );
  MUX2X1 U777 ( .B(n855), .A(n788), .S(n757), .Y(B[51]) );
  MUX2X1 U778 ( .B(n856), .A(n788), .S(n757), .Y(B[50]) );
  MUX2X1 U779 ( .B(n793), .A(n857), .S(n757), .Y(B[4]) );
  MUX2X1 U780 ( .B(n859), .A(n860), .S(n752), .Y(n858) );
  MUX2X1 U781 ( .B(n861), .A(n862), .S(n746), .Y(n859) );
  MUX2X1 U782 ( .B(n863), .A(n788), .S(n757), .Y(B[49]) );
  MUX2X1 U783 ( .B(n864), .A(n788), .S(n757), .Y(B[48]) );
  MUX2X1 U784 ( .B(n865), .A(n788), .S(n757), .Y(B[47]) );
  MUX2X1 U785 ( .B(n866), .A(n838), .S(n757), .Y(B[46]) );
  MUX2X1 U786 ( .B(n867), .A(A[63]), .S(n752), .Y(n838) );
  MUX2X1 U787 ( .B(n868), .A(n839), .S(n757), .Y(B[45]) );
  MUX2X1 U788 ( .B(n869), .A(A[63]), .S(n752), .Y(n839) );
  MUX2X1 U789 ( .B(n870), .A(n840), .S(n757), .Y(B[44]) );
  MUX2X1 U790 ( .B(n871), .A(A[63]), .S(n752), .Y(n840) );
  MUX2X1 U791 ( .B(n872), .A(n847), .S(n757), .Y(B[43]) );
  MUX2X1 U792 ( .B(n873), .A(A[63]), .S(n752), .Y(n847) );
  MUX2X1 U793 ( .B(n874), .A(n848), .S(n757), .Y(B[42]) );
  MUX2X1 U794 ( .B(n875), .A(B[63]), .S(n752), .Y(n848) );
  MUX2X1 U795 ( .B(n876), .A(n849), .S(n756), .Y(B[41]) );
  MUX2X1 U796 ( .B(n877), .A(B[63]), .S(n752), .Y(n849) );
  MUX2X1 U797 ( .B(n878), .A(n850), .S(n756), .Y(B[40]) );
  MUX2X1 U798 ( .B(n879), .A(B[63]), .S(n752), .Y(n850) );
  MUX2X1 U799 ( .B(n880), .A(n881), .S(n756), .Y(B[3]) );
  MUX2X1 U800 ( .B(n882), .A(n883), .S(n752), .Y(n880) );
  MUX2X1 U801 ( .B(n792), .A(n796), .S(n746), .Y(n882) );
  MUX2X1 U802 ( .B(n885), .A(n886), .S(n736), .Y(n884) );
  MUX2X1 U803 ( .B(n888), .A(n889), .S(n738), .Y(n887) );
  MUX2X1 U804 ( .B(n890), .A(n851), .S(n756), .Y(B[39]) );
  MUX2X1 U805 ( .B(n891), .A(B[63]), .S(n752), .Y(n851) );
  MUX2X1 U806 ( .B(n892), .A(n852), .S(n756), .Y(B[38]) );
  MUX2X1 U807 ( .B(n893), .A(n867), .S(n751), .Y(n852) );
  MUX2X1 U808 ( .B(n894), .A(n788), .S(n746), .Y(n867) );
  MUX2X1 U809 ( .B(n895), .A(n853), .S(n756), .Y(B[37]) );
  MUX2X1 U810 ( .B(n896), .A(n869), .S(n751), .Y(n853) );
  MUX2X1 U811 ( .B(n897), .A(n788), .S(n746), .Y(n869) );
  MUX2X1 U812 ( .B(n898), .A(n854), .S(n756), .Y(B[36]) );
  MUX2X1 U813 ( .B(n899), .A(n871), .S(n751), .Y(n854) );
  MUX2X1 U814 ( .B(n900), .A(n788), .S(n746), .Y(n871) );
  MUX2X1 U815 ( .B(n901), .A(n855), .S(n756), .Y(B[35]) );
  MUX2X1 U816 ( .B(n902), .A(n873), .S(n751), .Y(n855) );
  MUX2X1 U817 ( .B(n903), .A(n788), .S(n746), .Y(n873) );
  MUX2X1 U818 ( .B(n904), .A(n856), .S(n756), .Y(B[34]) );
  MUX2X1 U819 ( .B(n905), .A(n875), .S(n751), .Y(n856) );
  MUX2X1 U820 ( .B(n906), .A(n894), .S(n746), .Y(n875) );
  MUX2X1 U821 ( .B(n907), .A(B[63]), .S(n736), .Y(n894) );
  MUX2X1 U822 ( .B(n908), .A(n863), .S(n756), .Y(B[33]) );
  MUX2X1 U823 ( .B(n909), .A(n877), .S(n751), .Y(n863) );
  MUX2X1 U824 ( .B(n910), .A(n897), .S(n746), .Y(n877) );
  MUX2X1 U825 ( .B(n911), .A(B[63]), .S(n740), .Y(n897) );
  MUX2X1 U826 ( .B(n912), .A(n864), .S(n756), .Y(B[32]) );
  MUX2X1 U827 ( .B(n913), .A(n879), .S(n751), .Y(n864) );
  MUX2X1 U828 ( .B(n914), .A(n900), .S(n746), .Y(n879) );
  MUX2X1 U829 ( .B(n915), .A(n907), .S(n740), .Y(n900) );
  MUX2X1 U830 ( .B(n786), .A(n788), .S(n732), .Y(n907) );
  MUX2X1 U831 ( .B(n916), .A(n865), .S(n756), .Y(B[31]) );
  MUX2X1 U832 ( .B(n917), .A(n891), .S(n751), .Y(n865) );
  MUX2X1 U833 ( .B(n918), .A(n903), .S(n746), .Y(n891) );
  MUX2X1 U834 ( .B(n919), .A(n911), .S(n740), .Y(n903) );
  MUX2X1 U835 ( .B(n785), .A(n786), .S(n732), .Y(n911) );
  MUX2X1 U836 ( .B(n920), .A(n866), .S(n755), .Y(B[30]) );
  MUX2X1 U837 ( .B(n921), .A(n893), .S(n751), .Y(n866) );
  MUX2X1 U838 ( .B(n922), .A(n906), .S(n746), .Y(n893) );
  MUX2X1 U839 ( .B(n923), .A(n915), .S(n740), .Y(n906) );
  MUX2X1 U840 ( .B(n784), .A(n785), .S(n732), .Y(n915) );
  MUX2X1 U841 ( .B(n924), .A(n925), .S(n755), .Y(B[2]) );
  MUX2X1 U842 ( .B(n926), .A(n927), .S(n751), .Y(n924) );
  MUX2X1 U843 ( .B(n791), .A(n795), .S(n746), .Y(n926) );
  MUX2X1 U844 ( .B(n929), .A(n930), .S(n740), .Y(n928) );
  MUX2X1 U845 ( .B(n932), .A(n933), .S(n740), .Y(n931) );
  MUX2X1 U846 ( .B(n934), .A(n868), .S(n755), .Y(B[29]) );
  MUX2X1 U847 ( .B(n935), .A(n896), .S(n751), .Y(n868) );
  MUX2X1 U848 ( .B(n936), .A(n910), .S(n745), .Y(n896) );
  MUX2X1 U849 ( .B(n937), .A(n919), .S(n740), .Y(n910) );
  MUX2X1 U850 ( .B(n783), .A(n784), .S(n734), .Y(n919) );
  MUX2X1 U851 ( .B(n938), .A(n870), .S(n755), .Y(B[28]) );
  MUX2X1 U852 ( .B(n939), .A(n899), .S(n751), .Y(n870) );
  MUX2X1 U853 ( .B(n940), .A(n914), .S(n745), .Y(n899) );
  MUX2X1 U854 ( .B(n941), .A(n923), .S(n740), .Y(n914) );
  MUX2X1 U855 ( .B(n782), .A(n783), .S(n734), .Y(n923) );
  MUX2X1 U856 ( .B(n942), .A(n872), .S(n755), .Y(B[27]) );
  MUX2X1 U857 ( .B(n943), .A(n902), .S(n750), .Y(n872) );
  MUX2X1 U858 ( .B(n944), .A(n918), .S(n745), .Y(n902) );
  MUX2X1 U859 ( .B(n945), .A(n937), .S(n740), .Y(n918) );
  MUX2X1 U860 ( .B(n781), .A(n782), .S(n734), .Y(n937) );
  MUX2X1 U861 ( .B(n946), .A(n874), .S(n755), .Y(B[26]) );
  MUX2X1 U862 ( .B(n947), .A(n905), .S(n750), .Y(n874) );
  MUX2X1 U863 ( .B(n948), .A(n922), .S(n745), .Y(n905) );
  MUX2X1 U864 ( .B(n949), .A(n941), .S(n740), .Y(n922) );
  MUX2X1 U865 ( .B(n780), .A(n781), .S(n734), .Y(n941) );
  MUX2X1 U866 ( .B(n826), .A(n876), .S(n755), .Y(B[25]) );
  MUX2X1 U867 ( .B(n950), .A(n909), .S(n750), .Y(n876) );
  MUX2X1 U868 ( .B(n951), .A(n936), .S(n745), .Y(n909) );
  MUX2X1 U869 ( .B(n952), .A(n945), .S(n740), .Y(n936) );
  MUX2X1 U870 ( .B(n779), .A(n780), .S(n734), .Y(n945) );
  MUX2X1 U871 ( .B(n953), .A(n954), .S(n750), .Y(n826) );
  MUX2X1 U872 ( .B(n828), .A(n878), .S(n755), .Y(B[24]) );
  MUX2X1 U873 ( .B(n955), .A(n913), .S(n750), .Y(n878) );
  MUX2X1 U874 ( .B(n956), .A(n940), .S(n745), .Y(n913) );
  MUX2X1 U875 ( .B(n957), .A(n949), .S(n740), .Y(n940) );
  MUX2X1 U876 ( .B(n778), .A(n779), .S(n734), .Y(n949) );
  MUX2X1 U877 ( .B(n958), .A(n959), .S(n750), .Y(n828) );
  MUX2X1 U878 ( .B(n831), .A(n890), .S(n755), .Y(B[23]) );
  MUX2X1 U879 ( .B(n960), .A(n917), .S(n750), .Y(n890) );
  MUX2X1 U880 ( .B(n961), .A(n944), .S(n745), .Y(n917) );
  MUX2X1 U881 ( .B(n962), .A(n952), .S(n739), .Y(n944) );
  MUX2X1 U882 ( .B(n777), .A(n778), .S(n734), .Y(n952) );
  MUX2X1 U883 ( .B(n963), .A(n964), .S(n750), .Y(n831) );
  MUX2X1 U884 ( .B(n835), .A(n892), .S(n755), .Y(B[22]) );
  MUX2X1 U885 ( .B(n965), .A(n921), .S(n750), .Y(n892) );
  MUX2X1 U886 ( .B(n966), .A(n948), .S(n745), .Y(n921) );
  MUX2X1 U887 ( .B(n967), .A(n957), .S(n739), .Y(n948) );
  MUX2X1 U888 ( .B(n776), .A(n777), .S(n734), .Y(n957) );
  MUX2X1 U889 ( .B(n968), .A(n969), .S(n750), .Y(n835) );
  MUX2X1 U890 ( .B(n841), .A(n895), .S(n755), .Y(B[21]) );
  MUX2X1 U891 ( .B(n970), .A(n935), .S(n750), .Y(n895) );
  MUX2X1 U892 ( .B(n971), .A(n951), .S(n745), .Y(n935) );
  MUX2X1 U893 ( .B(n972), .A(n962), .S(n739), .Y(n951) );
  MUX2X1 U894 ( .B(n775), .A(n776), .S(n734), .Y(n962) );
  MUX2X1 U895 ( .B(n973), .A(n974), .S(n750), .Y(n841) );
  MUX2X1 U896 ( .B(n857), .A(n898), .S(n755), .Y(B[20]) );
  MUX2X1 U897 ( .B(n975), .A(n939), .S(n749), .Y(n898) );
  MUX2X1 U898 ( .B(n976), .A(n956), .S(n745), .Y(n939) );
  MUX2X1 U899 ( .B(n977), .A(n967), .S(n739), .Y(n956) );
  MUX2X1 U900 ( .B(n774), .A(n775), .S(n734), .Y(n967) );
  MUX2X1 U901 ( .B(n978), .A(n979), .S(n749), .Y(n857) );
  MUX2X1 U902 ( .B(n980), .A(n981), .S(n754), .Y(B[1]) );
  MUX2X1 U903 ( .B(n790), .A(n798), .S(n749), .Y(n980) );
  MUX2X1 U904 ( .B(n846), .A(n983), .S(n745), .Y(n982) );
  MUX2X1 U905 ( .B(n886), .A(n984), .S(n739), .Y(n846) );
  MUX2X1 U906 ( .B(A[9]), .A(A[10]), .S(n734), .Y(n886) );
  MUX2X1 U907 ( .B(n986), .A(n845), .S(n745), .Y(n985) );
  MUX2X1 U908 ( .B(n889), .A(n885), .S(n739), .Y(n845) );
  MUX2X1 U909 ( .B(A[7]), .A(A[8]), .S(n734), .Y(n885) );
  MUX2X1 U910 ( .B(A[5]), .A(A[6]), .S(n733), .Y(n889) );
  MUX2X1 U911 ( .B(n987), .A(n888), .S(n739), .Y(n986) );
  MUX2X1 U912 ( .B(A[3]), .A(A[4]), .S(n733), .Y(n888) );
  MUX2X1 U913 ( .B(A[1]), .A(A[2]), .S(n733), .Y(n987) );
  MUX2X1 U914 ( .B(n881), .A(n901), .S(n754), .Y(B[19]) );
  MUX2X1 U915 ( .B(n988), .A(n943), .S(n749), .Y(n901) );
  MUX2X1 U916 ( .B(n989), .A(n961), .S(n744), .Y(n943) );
  MUX2X1 U917 ( .B(n990), .A(n972), .S(n739), .Y(n961) );
  MUX2X1 U918 ( .B(n773), .A(n774), .S(n733), .Y(n972) );
  MUX2X1 U919 ( .B(n991), .A(n992), .S(n749), .Y(n881) );
  MUX2X1 U920 ( .B(n925), .A(n904), .S(n754), .Y(B[18]) );
  MUX2X1 U921 ( .B(n993), .A(n947), .S(n749), .Y(n904) );
  MUX2X1 U922 ( .B(n994), .A(n966), .S(n744), .Y(n947) );
  MUX2X1 U923 ( .B(n995), .A(n977), .S(n739), .Y(n966) );
  MUX2X1 U924 ( .B(n772), .A(n773), .S(n733), .Y(n977) );
  MUX2X1 U925 ( .B(n996), .A(n997), .S(n749), .Y(n925) );
  MUX2X1 U926 ( .B(n981), .A(n908), .S(n754), .Y(B[17]) );
  MUX2X1 U927 ( .B(n954), .A(n950), .S(n749), .Y(n908) );
  MUX2X1 U928 ( .B(n998), .A(n971), .S(n744), .Y(n950) );
  MUX2X1 U929 ( .B(n999), .A(n990), .S(n739), .Y(n971) );
  MUX2X1 U930 ( .B(n771), .A(n772), .S(n733), .Y(n990) );
  MUX2X1 U931 ( .B(n1000), .A(n1001), .S(n744), .Y(n954) );
  MUX2X1 U932 ( .B(n806), .A(n953), .S(n749), .Y(n981) );
  MUX2X1 U933 ( .B(n814), .A(n1002), .S(n744), .Y(n953) );
  MUX2X1 U934 ( .B(n1004), .A(n1005), .S(n744), .Y(n1003) );
  MUX2X1 U935 ( .B(n1006), .A(n912), .S(n754), .Y(B[16]) );
  MUX2X1 U936 ( .B(n959), .A(n955), .S(n749), .Y(n912) );
  MUX2X1 U937 ( .B(n1007), .A(n976), .S(n744), .Y(n955) );
  MUX2X1 U938 ( .B(n1008), .A(n995), .S(n739), .Y(n976) );
  MUX2X1 U939 ( .B(n770), .A(n771), .S(n733), .Y(n995) );
  MUX2X1 U940 ( .B(n1009), .A(n1010), .S(n744), .Y(n959) );
  MUX2X1 U941 ( .B(n1011), .A(n916), .S(n754), .Y(B[15]) );
  MUX2X1 U942 ( .B(n964), .A(n960), .S(n749), .Y(n916) );
  MUX2X1 U943 ( .B(n1012), .A(n989), .S(n744), .Y(n960) );
  MUX2X1 U944 ( .B(n1013), .A(n999), .S(n739), .Y(n989) );
  MUX2X1 U945 ( .B(n769), .A(n770), .S(n733), .Y(n999) );
  MUX2X1 U946 ( .B(n1014), .A(n1015), .S(n744), .Y(n964) );
  MUX2X1 U947 ( .B(n833), .A(n963), .S(n749), .Y(n1011) );
  MUX2X1 U948 ( .B(n812), .A(n1016), .S(n744), .Y(n963) );
  MUX2X1 U949 ( .B(n804), .A(n808), .S(n744), .Y(n833) );
  MUX2X1 U950 ( .B(n1017), .A(n920), .S(n754), .Y(B[14]) );
  MUX2X1 U951 ( .B(n969), .A(n965), .S(n748), .Y(n920) );
  MUX2X1 U952 ( .B(n1018), .A(n994), .S(n744), .Y(n965) );
  MUX2X1 U953 ( .B(n1019), .A(n1008), .S(n738), .Y(n994) );
  MUX2X1 U954 ( .B(n768), .A(n769), .S(n733), .Y(n1008) );
  MUX2X1 U955 ( .B(n1020), .A(n1021), .S(n746), .Y(n969) );
  MUX2X1 U956 ( .B(n837), .A(n968), .S(n748), .Y(n1017) );
  MUX2X1 U957 ( .B(n811), .A(n1022), .S(n743), .Y(n968) );
  MUX2X1 U958 ( .B(n803), .A(n807), .S(n745), .Y(n837) );
  MUX2X1 U959 ( .B(n1023), .A(n934), .S(n754), .Y(B[13]) );
  MUX2X1 U960 ( .B(n974), .A(n970), .S(n748), .Y(n934) );
  MUX2X1 U961 ( .B(n1001), .A(n998), .S(SH[2]), .Y(n970) );
  MUX2X1 U962 ( .B(n1024), .A(n1013), .S(n738), .Y(n998) );
  MUX2X1 U963 ( .B(n767), .A(n768), .S(n733), .Y(n1013) );
  MUX2X1 U964 ( .B(n1025), .A(n1026), .S(n738), .Y(n1001) );
  MUX2X1 U965 ( .B(n1002), .A(n1000), .S(SH[2]), .Y(n974) );
  MUX2X1 U966 ( .B(n822), .A(n824), .S(n738), .Y(n1000) );
  MUX2X1 U967 ( .B(n818), .A(n820), .S(n738), .Y(n1002) );
  MUX2X1 U968 ( .B(n802), .A(n973), .S(n748), .Y(n1023) );
  MUX2X1 U969 ( .B(n810), .A(n814), .S(SH[2]), .Y(n973) );
  MUX2X1 U970 ( .B(n1028), .A(n1029), .S(n738), .Y(n1027) );
  MUX2X1 U971 ( .B(n1030), .A(n1031), .S(n738), .Y(n1005) );
  MUX2X1 U972 ( .B(n983), .A(n1004), .S(SH[2]), .Y(n844) );
  MUX2X1 U973 ( .B(n1032), .A(n1033), .S(n738), .Y(n1004) );
  MUX2X1 U974 ( .B(n1034), .A(n1035), .S(n738), .Y(n983) );
  MUX2X1 U975 ( .B(n1036), .A(n938), .S(n754), .Y(B[12]) );
  MUX2X1 U976 ( .B(n979), .A(n975), .S(n748), .Y(n938) );
  MUX2X1 U977 ( .B(n1010), .A(n1007), .S(SH[2]), .Y(n975) );
  MUX2X1 U978 ( .B(n1037), .A(n1019), .S(n738), .Y(n1007) );
  MUX2X1 U979 ( .B(n766), .A(n767), .S(n733), .Y(n1019) );
  MUX2X1 U980 ( .B(n1038), .A(n1039), .S(n738), .Y(n1010) );
  MUX2X1 U981 ( .B(n1040), .A(n1009), .S(SH[2]), .Y(n979) );
  MUX2X1 U982 ( .B(n821), .A(n823), .S(n738), .Y(n1009) );
  MUX2X1 U983 ( .B(n801), .A(n978), .S(n748), .Y(n1036) );
  MUX2X1 U984 ( .B(n809), .A(n813), .S(SH[2]), .Y(n978) );
  MUX2X1 U985 ( .B(n1041), .A(n1042), .S(SH[2]), .Y(n860) );
  MUX2X1 U986 ( .B(n1043), .A(n942), .S(n754), .Y(B[11]) );
  MUX2X1 U987 ( .B(n992), .A(n988), .S(n748), .Y(n942) );
  MUX2X1 U988 ( .B(n1015), .A(n1012), .S(n743), .Y(n988) );
  MUX2X1 U989 ( .B(n1026), .A(n1024), .S(n737), .Y(n1012) );
  MUX2X1 U990 ( .B(n765), .A(n766), .S(n733), .Y(n1024) );
  MUX2X1 U991 ( .B(n763), .A(n764), .S(n732), .Y(n1026) );
  MUX2X1 U992 ( .B(n824), .A(n1025), .S(n737), .Y(n1015) );
  MUX2X1 U993 ( .B(n761), .A(n762), .S(n732), .Y(n1025) );
  MUX2X1 U994 ( .B(A[35]), .A(A[36]), .S(n732), .Y(n1044) );
  MUX2X1 U995 ( .B(n1016), .A(n1014), .S(n743), .Y(n992) );
  MUX2X1 U996 ( .B(n820), .A(n822), .S(n737), .Y(n1014) );
  MUX2X1 U997 ( .B(A[33]), .A(A[34]), .S(n732), .Y(n1045) );
  MUX2X1 U998 ( .B(A[31]), .A(A[32]), .S(n732), .Y(n1046) );
  MUX2X1 U999 ( .B(n816), .A(n818), .S(n737), .Y(n1016) );
  MUX2X1 U1000 ( .B(A[29]), .A(A[30]), .S(n732), .Y(n1047) );
  MUX2X1 U1001 ( .B(A[27]), .A(A[28]), .S(n732), .Y(n1029) );
  MUX2X1 U1002 ( .B(n883), .A(n991), .S(n748), .Y(n1043) );
  MUX2X1 U1003 ( .B(n808), .A(n812), .S(n743), .Y(n991) );
  MUX2X1 U1004 ( .B(n1031), .A(n1028), .S(n737), .Y(n1048) );
  MUX2X1 U1005 ( .B(A[25]), .A(A[26]), .S(n732), .Y(n1028) );
  MUX2X1 U1006 ( .B(A[23]), .A(A[24]), .S(n732), .Y(n1031) );
  MUX2X1 U1007 ( .B(n1033), .A(n1030), .S(n737), .Y(n1049) );
  MUX2X1 U1008 ( .B(A[21]), .A(A[22]), .S(n732), .Y(n1030) );
  MUX2X1 U1009 ( .B(A[19]), .A(A[20]), .S(n732), .Y(n1033) );
  MUX2X1 U1010 ( .B(n800), .A(n804), .S(n743), .Y(n883) );
  MUX2X1 U1011 ( .B(n1035), .A(n1032), .S(n737), .Y(n1050) );
  MUX2X1 U1012 ( .B(A[17]), .A(A[18]), .S(n732), .Y(n1032) );
  MUX2X1 U1013 ( .B(A[15]), .A(A[16]), .S(n731), .Y(n1035) );
  MUX2X1 U1014 ( .B(n984), .A(n1034), .S(n737), .Y(n1051) );
  MUX2X1 U1015 ( .B(A[13]), .A(A[14]), .S(n731), .Y(n1034) );
  MUX2X1 U1016 ( .B(A[11]), .A(A[12]), .S(n731), .Y(n984) );
  MUX2X1 U1017 ( .B(n1052), .A(n946), .S(n754), .Y(B[10]) );
  MUX2X1 U1018 ( .B(n997), .A(n993), .S(n748), .Y(n946) );
  MUX2X1 U1019 ( .B(n1021), .A(n1018), .S(n743), .Y(n993) );
  MUX2X1 U1020 ( .B(n1039), .A(n1037), .S(n737), .Y(n1018) );
  MUX2X1 U1021 ( .B(n764), .A(n765), .S(n731), .Y(n1037) );
  MUX2X1 U1022 ( .B(n762), .A(n763), .S(n731), .Y(n1039) );
  MUX2X1 U1023 ( .B(n823), .A(n1038), .S(n737), .Y(n1021) );
  MUX2X1 U1024 ( .B(n760), .A(n761), .S(n731), .Y(n1038) );
  MUX2X1 U1025 ( .B(A[34]), .A(A[35]), .S(n731), .Y(n1053) );
  MUX2X1 U1026 ( .B(n1022), .A(n1020), .S(n743), .Y(n997) );
  MUX2X1 U1027 ( .B(n819), .A(n821), .S(n737), .Y(n1020) );
  MUX2X1 U1028 ( .B(A[32]), .A(A[33]), .S(n731), .Y(n1054) );
  MUX2X1 U1029 ( .B(n815), .A(n817), .S(n737), .Y(n1022) );
  MUX2X1 U1030 ( .B(n927), .A(n996), .S(n748), .Y(n1052) );
  MUX2X1 U1031 ( .B(n807), .A(n811), .S(n743), .Y(n996) );
  MUX2X1 U1032 ( .B(n1057), .A(n1058), .S(n736), .Y(n1056) );
  MUX2X1 U1033 ( .B(n1060), .A(n1061), .S(n736), .Y(n1059) );
  MUX2X1 U1034 ( .B(n799), .A(n803), .S(n743), .Y(n927) );
  MUX2X1 U1035 ( .B(n1063), .A(n1064), .S(n736), .Y(n1062) );
  MUX2X1 U1036 ( .B(n1066), .A(n1067), .S(n736), .Y(n1065) );
  MUX2X1 U1037 ( .B(n1068), .A(n1006), .S(n754), .Y(B[0]) );
  MUX2X1 U1038 ( .B(n829), .A(n958), .S(n748), .Y(n1006) );
  MUX2X1 U1039 ( .B(n813), .A(n1040), .S(n743), .Y(n958) );
  MUX2X1 U1040 ( .B(n817), .A(n819), .S(n736), .Y(n1040) );
  MUX2X1 U1041 ( .B(A[30]), .A(A[31]), .S(n731), .Y(n1069) );
  MUX2X1 U1042 ( .B(A[28]), .A(A[29]), .S(n731), .Y(n1070) );
  MUX2X1 U1043 ( .B(n1058), .A(n1055), .S(n736), .Y(n1071) );
  MUX2X1 U1044 ( .B(A[26]), .A(A[27]), .S(n731), .Y(n1055) );
  MUX2X1 U1045 ( .B(A[24]), .A(A[25]), .S(n731), .Y(n1058) );
  MUX2X1 U1046 ( .B(n805), .A(n809), .S(n743), .Y(n829) );
  MUX2X1 U1047 ( .B(n1061), .A(n1057), .S(n736), .Y(n1072) );
  MUX2X1 U1048 ( .B(A[22]), .A(A[23]), .S(n731), .Y(n1057) );
  MUX2X1 U1049 ( .B(A[20]), .A(A[21]), .S(n733), .Y(n1061) );
  MUX2X1 U1050 ( .B(n1064), .A(n1060), .S(n736), .Y(n1042) );
  MUX2X1 U1051 ( .B(A[18]), .A(A[19]), .S(n734), .Y(n1060) );
  MUX2X1 U1052 ( .B(A[16]), .A(A[17]), .S(n733), .Y(n1064) );
  MUX2X1 U1053 ( .B(n789), .A(n797), .S(n748), .Y(n1068) );
  MUX2X1 U1054 ( .B(n862), .A(n1041), .S(n743), .Y(n1073) );
  MUX2X1 U1055 ( .B(n1067), .A(n1063), .S(n736), .Y(n1041) );
  MUX2X1 U1056 ( .B(A[14]), .A(A[15]), .S(n734), .Y(n1063) );
  MUX2X1 U1057 ( .B(A[12]), .A(A[13]), .S(n731), .Y(n1067) );
  MUX2X1 U1058 ( .B(n930), .A(n1066), .S(n736), .Y(n862) );
  MUX2X1 U1059 ( .B(A[10]), .A(A[11]), .S(n733), .Y(n1066) );
  MUX2X1 U1060 ( .B(A[8]), .A(A[9]), .S(n734), .Y(n930) );
  MUX2X1 U1061 ( .B(n1075), .A(n861), .S(n743), .Y(n1074) );
  MUX2X1 U1062 ( .B(n933), .A(n929), .S(n736), .Y(n861) );
  MUX2X1 U1063 ( .B(A[6]), .A(A[7]), .S(n733), .Y(n929) );
  MUX2X1 U1064 ( .B(A[4]), .A(A[5]), .S(n732), .Y(n933) );
  MUX2X1 U1065 ( .B(n1076), .A(n932), .S(n736), .Y(n1075) );
  MUX2X1 U1066 ( .B(A[2]), .A(A[3]), .S(SH[0]), .Y(n932) );
  MUX2X1 U1067 ( .B(A[0]), .A(A[1]), .S(SH[0]), .Y(n1076) );
endmodule


module alu_DW_rightsh_1 ( A, DATA_TC, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC;
  wire   n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539;
  assign B[31] = A[31];

  INVX1 U329 ( .A(n431), .Y(n393) );
  INVX1 U330 ( .A(n485), .Y(n408) );
  INVX1 U331 ( .A(n500), .Y(n404) );
  INVX1 U332 ( .A(n505), .Y(n396) );
  INVX1 U333 ( .A(n429), .Y(n389) );
  INVX1 U334 ( .A(n417), .Y(n400) );
  INVX1 U335 ( .A(n488), .Y(B[16]) );
  INVX1 U336 ( .A(n535), .Y(B[0]) );
  INVX1 U337 ( .A(n434), .Y(n388) );
  INVX1 U338 ( .A(n454), .Y(n385) );
  INVX1 U339 ( .A(n421), .Y(n390) );
  INVX1 U340 ( .A(n437), .Y(n387) );
  INVX1 U341 ( .A(n498), .Y(n412) );
  INVX1 U342 ( .A(n465), .Y(n406) );
  INVX1 U343 ( .A(n527), .Y(n401) );
  INVX1 U344 ( .A(n512), .Y(n395) );
  INVX1 U345 ( .A(n518), .Y(n394) );
  INVX1 U346 ( .A(n418), .Y(n391) );
  INVX1 U347 ( .A(n470), .Y(n403) );
  INVX1 U348 ( .A(n480), .Y(n402) );
  INVX1 U349 ( .A(n370), .Y(n369) );
  INVX1 U350 ( .A(n375), .Y(n374) );
  INVX1 U351 ( .A(n520), .Y(n413) );
  INVX1 U352 ( .A(n510), .Y(n411) );
  INVX1 U353 ( .A(n517), .Y(n410) );
  INVX1 U354 ( .A(n463), .Y(n407) );
  INVX1 U355 ( .A(n530), .Y(n397) );
  INVX1 U356 ( .A(n521), .Y(n409) );
  INVX1 U357 ( .A(n524), .Y(n405) );
  INVX1 U358 ( .A(n442), .Y(n386) );
  INVX1 U359 ( .A(n415), .Y(n392) );
  INVX1 U360 ( .A(n490), .Y(n398) );
  INVX1 U361 ( .A(n474), .Y(n384) );
  INVX1 U362 ( .A(n378), .Y(n376) );
  INVX1 U363 ( .A(n378), .Y(n377) );
  INVX1 U364 ( .A(n373), .Y(n372) );
  INVX1 U365 ( .A(n373), .Y(n371) );
  INVX1 U366 ( .A(A[31]), .Y(n382) );
  INVX1 U367 ( .A(SH[0]), .Y(n370) );
  INVX1 U368 ( .A(SH[2]), .Y(n375) );
  INVX1 U369 ( .A(SH[3]), .Y(n378) );
  INVX1 U370 ( .A(SH[1]), .Y(n373) );
  INVX1 U371 ( .A(n381), .Y(n380) );
  INVX1 U372 ( .A(n381), .Y(n379) );
  INVX1 U373 ( .A(SH[4]), .Y(n381) );
  MUX2X1 U374 ( .B(n392), .A(n414), .S(n380), .Y(B[9]) );
  MUX2X1 U375 ( .B(n416), .A(n417), .S(n376), .Y(n415) );
  MUX2X1 U376 ( .B(n391), .A(n407), .S(SH[4]), .Y(B[8]) );
  MUX2X1 U377 ( .B(n419), .A(n420), .S(SH[3]), .Y(n418) );
  MUX2X1 U378 ( .B(n390), .A(n406), .S(SH[4]), .Y(B[7]) );
  MUX2X1 U379 ( .B(n422), .A(n423), .S(SH[3]), .Y(n421) );
  MUX2X1 U380 ( .B(n424), .A(n425), .S(SH[2]), .Y(n422) );
  MUX2X1 U381 ( .B(n426), .A(n427), .S(SH[4]), .Y(B[6]) );
  MUX2X1 U382 ( .B(n389), .A(n428), .S(n376), .Y(n426) );
  MUX2X1 U383 ( .B(n430), .A(n431), .S(n374), .Y(n429) );
  MUX2X1 U384 ( .B(n432), .A(n433), .S(SH[4]), .Y(B[5]) );
  MUX2X1 U385 ( .B(n388), .A(n396), .S(n376), .Y(n432) );
  MUX2X1 U386 ( .B(n435), .A(n436), .S(SH[2]), .Y(n434) );
  MUX2X1 U387 ( .B(n387), .A(n403), .S(SH[4]), .Y(B[4]) );
  MUX2X1 U388 ( .B(n438), .A(n439), .S(SH[3]), .Y(n437) );
  MUX2X1 U389 ( .B(n440), .A(n441), .S(SH[2]), .Y(n438) );
  MUX2X1 U390 ( .B(n386), .A(n402), .S(SH[4]), .Y(B[3]) );
  MUX2X1 U391 ( .B(n443), .A(n444), .S(SH[3]), .Y(n442) );
  MUX2X1 U392 ( .B(n445), .A(n424), .S(SH[2]), .Y(n443) );
  MUX2X1 U393 ( .B(n446), .A(n447), .S(SH[1]), .Y(n424) );
  MUX2X1 U394 ( .B(n448), .A(n449), .S(SH[1]), .Y(n445) );
  MUX2X1 U395 ( .B(n450), .A(n382), .S(n380), .Y(B[30]) );
  MUX2X1 U396 ( .B(n451), .A(n452), .S(n380), .Y(B[2]) );
  MUX2X1 U397 ( .B(n385), .A(n453), .S(n377), .Y(n451) );
  MUX2X1 U398 ( .B(n455), .A(n430), .S(n374), .Y(n454) );
  MUX2X1 U399 ( .B(n456), .A(n457), .S(n371), .Y(n430) );
  MUX2X1 U400 ( .B(n458), .A(n459), .S(SH[1]), .Y(n455) );
  MUX2X1 U401 ( .B(n460), .A(n382), .S(n380), .Y(B[29]) );
  MUX2X1 U402 ( .B(n411), .A(n382), .S(n380), .Y(B[28]) );
  MUX2X1 U403 ( .B(n410), .A(n382), .S(n380), .Y(B[27]) );
  MUX2X1 U404 ( .B(n461), .A(n382), .S(n380), .Y(B[26]) );
  MUX2X1 U405 ( .B(n414), .A(n382), .S(n380), .Y(B[25]) );
  MUX2X1 U406 ( .B(n462), .A(A[31]), .S(n377), .Y(n414) );
  MUX2X1 U407 ( .B(n407), .A(n382), .S(n380), .Y(B[24]) );
  MUX2X1 U408 ( .B(n464), .A(n382), .S(n377), .Y(n463) );
  MUX2X1 U409 ( .B(n406), .A(n382), .S(n380), .Y(B[23]) );
  MUX2X1 U410 ( .B(n466), .A(n382), .S(n377), .Y(n465) );
  MUX2X1 U411 ( .B(n427), .A(n382), .S(n380), .Y(B[22]) );
  MUX2X1 U412 ( .B(n467), .A(n468), .S(n377), .Y(n427) );
  MUX2X1 U413 ( .B(n433), .A(n382), .S(n380), .Y(B[21]) );
  MUX2X1 U414 ( .B(n404), .A(n469), .S(n377), .Y(n433) );
  MUX2X1 U415 ( .B(n403), .A(n382), .S(n380), .Y(B[20]) );
  MUX2X1 U416 ( .B(n471), .A(n472), .S(n377), .Y(n470) );
  MUX2X1 U417 ( .B(n384), .A(n473), .S(n379), .Y(B[1]) );
  MUX2X1 U418 ( .B(n475), .A(n416), .S(n377), .Y(n474) );
  MUX2X1 U419 ( .B(n436), .A(n476), .S(SH[2]), .Y(n416) );
  MUX2X1 U420 ( .B(n447), .A(n477), .S(SH[1]), .Y(n436) );
  MUX2X1 U421 ( .B(A[9]), .A(A[10]), .S(SH[0]), .Y(n447) );
  MUX2X1 U422 ( .B(n478), .A(n435), .S(SH[2]), .Y(n475) );
  MUX2X1 U423 ( .B(n449), .A(n446), .S(n372), .Y(n435) );
  MUX2X1 U424 ( .B(A[7]), .A(A[8]), .S(n369), .Y(n446) );
  MUX2X1 U425 ( .B(A[5]), .A(A[6]), .S(SH[0]), .Y(n449) );
  MUX2X1 U426 ( .B(n479), .A(n448), .S(SH[1]), .Y(n478) );
  MUX2X1 U427 ( .B(A[3]), .A(A[4]), .S(SH[0]), .Y(n448) );
  MUX2X1 U428 ( .B(A[1]), .A(A[2]), .S(SH[0]), .Y(n479) );
  MUX2X1 U429 ( .B(n402), .A(n382), .S(n379), .Y(B[19]) );
  MUX2X1 U430 ( .B(n481), .A(n482), .S(n377), .Y(n480) );
  MUX2X1 U431 ( .B(n452), .A(n382), .S(n379), .Y(B[18]) );
  MUX2X1 U432 ( .B(n483), .A(n484), .S(n377), .Y(n452) );
  MUX2X1 U433 ( .B(n473), .A(n382), .S(n379), .Y(B[17]) );
  MUX2X1 U434 ( .B(n400), .A(n462), .S(n377), .Y(n473) );
  MUX2X1 U435 ( .B(n408), .A(n412), .S(SH[2]), .Y(n462) );
  MUX2X1 U436 ( .B(n486), .A(n487), .S(SH[2]), .Y(n417) );
  MUX2X1 U437 ( .B(n489), .A(A[31]), .S(n379), .Y(n488) );
  MUX2X1 U438 ( .B(n398), .A(n382), .S(n379), .Y(B[15]) );
  MUX2X1 U439 ( .B(n423), .A(n466), .S(n377), .Y(n490) );
  MUX2X1 U440 ( .B(n491), .A(n492), .S(SH[2]), .Y(n466) );
  MUX2X1 U441 ( .B(n493), .A(n494), .S(SH[2]), .Y(n423) );
  MUX2X1 U442 ( .B(n495), .A(n450), .S(n379), .Y(B[14]) );
  MUX2X1 U443 ( .B(n468), .A(A[31]), .S(n376), .Y(n450) );
  MUX2X1 U444 ( .B(n496), .A(n382), .S(SH[2]), .Y(n468) );
  MUX2X1 U445 ( .B(n428), .A(n467), .S(n376), .Y(n495) );
  MUX2X1 U446 ( .B(n405), .A(n409), .S(SH[2]), .Y(n467) );
  MUX2X1 U447 ( .B(n397), .A(n401), .S(SH[2]), .Y(n428) );
  MUX2X1 U448 ( .B(n497), .A(n460), .S(n379), .Y(B[13]) );
  MUX2X1 U449 ( .B(n469), .A(A[31]), .S(n376), .Y(n460) );
  MUX2X1 U450 ( .B(n412), .A(n382), .S(SH[2]), .Y(n469) );
  MUX2X1 U451 ( .B(n499), .A(n382), .S(n372), .Y(n498) );
  MUX2X1 U452 ( .B(n396), .A(n404), .S(n376), .Y(n497) );
  MUX2X1 U453 ( .B(n487), .A(n485), .S(SH[2]), .Y(n500) );
  MUX2X1 U454 ( .B(n501), .A(n502), .S(n372), .Y(n485) );
  MUX2X1 U455 ( .B(n503), .A(n504), .S(n372), .Y(n487) );
  MUX2X1 U456 ( .B(n476), .A(n486), .S(SH[2]), .Y(n505) );
  MUX2X1 U457 ( .B(n506), .A(n507), .S(n372), .Y(n486) );
  MUX2X1 U458 ( .B(n508), .A(n509), .S(n372), .Y(n476) );
  MUX2X1 U459 ( .B(n395), .A(n411), .S(n379), .Y(B[12]) );
  MUX2X1 U460 ( .B(n472), .A(n382), .S(n376), .Y(n510) );
  MUX2X1 U461 ( .B(n511), .A(A[31]), .S(SH[2]), .Y(n472) );
  MUX2X1 U462 ( .B(n439), .A(n471), .S(n376), .Y(n512) );
  MUX2X1 U463 ( .B(n513), .A(n514), .S(n374), .Y(n471) );
  MUX2X1 U464 ( .B(n515), .A(n516), .S(n374), .Y(n439) );
  MUX2X1 U465 ( .B(n394), .A(n410), .S(n379), .Y(B[11]) );
  MUX2X1 U466 ( .B(n482), .A(n382), .S(n376), .Y(n517) );
  MUX2X1 U467 ( .B(n492), .A(A[31]), .S(n374), .Y(n482) );
  MUX2X1 U468 ( .B(n502), .A(n499), .S(n372), .Y(n492) );
  MUX2X1 U469 ( .B(A[29]), .A(A[30]), .S(SH[0]), .Y(n499) );
  MUX2X1 U470 ( .B(A[27]), .A(A[28]), .S(n369), .Y(n502) );
  MUX2X1 U471 ( .B(n444), .A(n481), .S(n376), .Y(n518) );
  MUX2X1 U472 ( .B(n494), .A(n491), .S(n374), .Y(n481) );
  MUX2X1 U473 ( .B(n504), .A(n501), .S(n372), .Y(n491) );
  MUX2X1 U474 ( .B(A[25]), .A(A[26]), .S(SH[0]), .Y(n501) );
  MUX2X1 U475 ( .B(A[23]), .A(A[24]), .S(SH[0]), .Y(n504) );
  MUX2X1 U476 ( .B(n507), .A(n503), .S(n372), .Y(n494) );
  MUX2X1 U477 ( .B(A[21]), .A(A[22]), .S(SH[0]), .Y(n503) );
  MUX2X1 U478 ( .B(A[19]), .A(A[20]), .S(SH[0]), .Y(n507) );
  MUX2X1 U479 ( .B(n425), .A(n493), .S(n374), .Y(n444) );
  MUX2X1 U480 ( .B(n509), .A(n506), .S(n372), .Y(n493) );
  MUX2X1 U481 ( .B(A[17]), .A(A[18]), .S(SH[0]), .Y(n506) );
  MUX2X1 U482 ( .B(A[15]), .A(A[16]), .S(SH[0]), .Y(n509) );
  MUX2X1 U483 ( .B(n477), .A(n508), .S(n372), .Y(n425) );
  MUX2X1 U484 ( .B(A[13]), .A(A[14]), .S(SH[0]), .Y(n508) );
  MUX2X1 U485 ( .B(A[11]), .A(A[12]), .S(SH[0]), .Y(n477) );
  MUX2X1 U486 ( .B(n519), .A(n461), .S(n379), .Y(B[10]) );
  MUX2X1 U487 ( .B(n484), .A(A[31]), .S(n376), .Y(n461) );
  MUX2X1 U488 ( .B(n409), .A(n496), .S(n374), .Y(n484) );
  MUX2X1 U489 ( .B(n413), .A(A[31]), .S(n372), .Y(n496) );
  MUX2X1 U490 ( .B(n522), .A(n523), .S(n372), .Y(n521) );
  MUX2X1 U491 ( .B(n453), .A(n483), .S(n376), .Y(n519) );
  MUX2X1 U492 ( .B(n401), .A(n405), .S(n374), .Y(n483) );
  MUX2X1 U493 ( .B(n525), .A(n526), .S(n371), .Y(n524) );
  MUX2X1 U494 ( .B(n528), .A(n529), .S(n371), .Y(n527) );
  MUX2X1 U495 ( .B(n393), .A(n397), .S(n374), .Y(n453) );
  MUX2X1 U496 ( .B(n531), .A(n532), .S(n371), .Y(n530) );
  MUX2X1 U497 ( .B(n533), .A(n534), .S(n371), .Y(n431) );
  MUX2X1 U498 ( .B(n536), .A(n489), .S(n379), .Y(n535) );
  MUX2X1 U499 ( .B(n420), .A(n464), .S(n376), .Y(n489) );
  MUX2X1 U500 ( .B(n514), .A(n511), .S(n374), .Y(n464) );
  MUX2X1 U501 ( .B(n523), .A(n520), .S(n371), .Y(n511) );
  MUX2X1 U502 ( .B(A[30]), .A(A[31]), .S(SH[0]), .Y(n520) );
  MUX2X1 U503 ( .B(A[28]), .A(A[29]), .S(SH[0]), .Y(n523) );
  MUX2X1 U504 ( .B(n526), .A(n522), .S(n371), .Y(n514) );
  MUX2X1 U505 ( .B(A[26]), .A(A[27]), .S(SH[0]), .Y(n522) );
  MUX2X1 U506 ( .B(A[24]), .A(A[25]), .S(SH[0]), .Y(n526) );
  MUX2X1 U507 ( .B(n516), .A(n513), .S(n374), .Y(n420) );
  MUX2X1 U508 ( .B(n529), .A(n525), .S(n371), .Y(n513) );
  MUX2X1 U509 ( .B(A[22]), .A(A[23]), .S(n369), .Y(n525) );
  MUX2X1 U510 ( .B(A[20]), .A(A[21]), .S(n369), .Y(n529) );
  MUX2X1 U511 ( .B(n532), .A(n528), .S(n371), .Y(n516) );
  MUX2X1 U512 ( .B(A[18]), .A(A[19]), .S(n369), .Y(n528) );
  MUX2X1 U513 ( .B(A[16]), .A(A[17]), .S(n369), .Y(n532) );
  MUX2X1 U514 ( .B(n537), .A(n419), .S(n376), .Y(n536) );
  MUX2X1 U515 ( .B(n441), .A(n515), .S(n374), .Y(n419) );
  MUX2X1 U516 ( .B(n534), .A(n531), .S(n371), .Y(n515) );
  MUX2X1 U517 ( .B(A[14]), .A(A[15]), .S(n369), .Y(n531) );
  MUX2X1 U518 ( .B(A[12]), .A(A[13]), .S(n369), .Y(n534) );
  MUX2X1 U519 ( .B(n457), .A(n533), .S(n371), .Y(n441) );
  MUX2X1 U520 ( .B(A[10]), .A(A[11]), .S(n369), .Y(n533) );
  MUX2X1 U521 ( .B(A[8]), .A(A[9]), .S(n369), .Y(n457) );
  MUX2X1 U522 ( .B(n538), .A(n440), .S(n374), .Y(n537) );
  MUX2X1 U523 ( .B(n459), .A(n456), .S(n371), .Y(n440) );
  MUX2X1 U524 ( .B(A[6]), .A(A[7]), .S(n369), .Y(n456) );
  MUX2X1 U525 ( .B(A[4]), .A(A[5]), .S(n369), .Y(n459) );
  MUX2X1 U526 ( .B(n539), .A(n458), .S(n371), .Y(n538) );
  MUX2X1 U527 ( .B(A[2]), .A(A[3]), .S(n369), .Y(n458) );
  MUX2X1 U528 ( .B(A[0]), .A(A[1]), .S(n369), .Y(n539) );
endmodule


module alu_DW_rightsh_2 ( A, DATA_TC, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC;
  wire   n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537;
  assign B[31] = A[31];

  INVX1 U329 ( .A(n427), .Y(n387) );
  INVX1 U330 ( .A(n498), .Y(n402) );
  INVX1 U331 ( .A(n429), .Y(n391) );
  INVX1 U332 ( .A(n415), .Y(n398) );
  INVX1 U333 ( .A(n486), .Y(B[16]) );
  INVX1 U334 ( .A(n533), .Y(B[0]) );
  INVX1 U335 ( .A(n432), .Y(n386) );
  INVX1 U336 ( .A(n452), .Y(n383) );
  INVX1 U337 ( .A(n419), .Y(n388) );
  INVX1 U338 ( .A(n435), .Y(n385) );
  INVX1 U339 ( .A(n508), .Y(n409) );
  INVX1 U340 ( .A(n515), .Y(n408) );
  INVX1 U341 ( .A(n461), .Y(n405) );
  INVX1 U342 ( .A(n463), .Y(n404) );
  INVX1 U343 ( .A(n522), .Y(n403) );
  INVX1 U344 ( .A(n488), .Y(n396) );
  INVX1 U345 ( .A(n510), .Y(n393) );
  INVX1 U346 ( .A(n516), .Y(n392) );
  INVX1 U347 ( .A(n416), .Y(n389) );
  INVX1 U348 ( .A(n373), .Y(n372) );
  INVX1 U349 ( .A(A[31]), .Y(n380) );
  INVX1 U350 ( .A(n518), .Y(n411) );
  INVX1 U351 ( .A(n483), .Y(n406) );
  INVX1 U352 ( .A(n503), .Y(n394) );
  INVX1 U353 ( .A(n468), .Y(n401) );
  INVX1 U354 ( .A(n478), .Y(n400) );
  INVX1 U355 ( .A(n440), .Y(n384) );
  INVX1 U356 ( .A(n413), .Y(n390) );
  INVX1 U357 ( .A(n472), .Y(n382) );
  INVX1 U358 ( .A(n376), .Y(n374) );
  INVX1 U359 ( .A(n376), .Y(n375) );
  INVX1 U360 ( .A(n371), .Y(n370) );
  INVX1 U361 ( .A(n371), .Y(n369) );
  INVX1 U362 ( .A(SH[2]), .Y(n373) );
  INVX1 U363 ( .A(n496), .Y(n410) );
  INVX1 U364 ( .A(n519), .Y(n407) );
  INVX1 U365 ( .A(n528), .Y(n395) );
  INVX1 U366 ( .A(n525), .Y(n399) );
  INVX1 U367 ( .A(SH[3]), .Y(n376) );
  INVX1 U368 ( .A(SH[1]), .Y(n371) );
  INVX1 U369 ( .A(n379), .Y(n378) );
  INVX1 U370 ( .A(n379), .Y(n377) );
  INVX1 U371 ( .A(SH[4]), .Y(n379) );
  MUX2X1 U372 ( .B(n390), .A(n412), .S(SH[4]), .Y(B[9]) );
  MUX2X1 U373 ( .B(n414), .A(n415), .S(SH[3]), .Y(n413) );
  MUX2X1 U374 ( .B(n389), .A(n405), .S(SH[4]), .Y(B[8]) );
  MUX2X1 U375 ( .B(n417), .A(n418), .S(SH[3]), .Y(n416) );
  MUX2X1 U376 ( .B(n388), .A(n404), .S(SH[4]), .Y(B[7]) );
  MUX2X1 U377 ( .B(n420), .A(n421), .S(SH[3]), .Y(n419) );
  MUX2X1 U378 ( .B(n422), .A(n423), .S(SH[2]), .Y(n420) );
  MUX2X1 U379 ( .B(n424), .A(n425), .S(SH[4]), .Y(B[6]) );
  MUX2X1 U380 ( .B(n387), .A(n426), .S(n374), .Y(n424) );
  MUX2X1 U381 ( .B(n428), .A(n429), .S(SH[2]), .Y(n427) );
  MUX2X1 U382 ( .B(n430), .A(n431), .S(SH[4]), .Y(B[5]) );
  MUX2X1 U383 ( .B(n386), .A(n394), .S(SH[3]), .Y(n430) );
  MUX2X1 U384 ( .B(n433), .A(n434), .S(SH[2]), .Y(n432) );
  MUX2X1 U385 ( .B(n385), .A(n401), .S(SH[4]), .Y(B[4]) );
  MUX2X1 U386 ( .B(n436), .A(n437), .S(SH[3]), .Y(n435) );
  MUX2X1 U387 ( .B(n438), .A(n439), .S(SH[2]), .Y(n436) );
  MUX2X1 U388 ( .B(n384), .A(n400), .S(SH[4]), .Y(B[3]) );
  MUX2X1 U389 ( .B(n441), .A(n442), .S(SH[3]), .Y(n440) );
  MUX2X1 U390 ( .B(n443), .A(n422), .S(SH[2]), .Y(n441) );
  MUX2X1 U391 ( .B(n444), .A(n445), .S(SH[1]), .Y(n422) );
  MUX2X1 U392 ( .B(n446), .A(n447), .S(SH[1]), .Y(n443) );
  MUX2X1 U393 ( .B(n448), .A(n380), .S(n378), .Y(B[30]) );
  MUX2X1 U394 ( .B(n449), .A(n450), .S(n378), .Y(B[2]) );
  MUX2X1 U395 ( .B(n383), .A(n451), .S(n375), .Y(n449) );
  MUX2X1 U396 ( .B(n453), .A(n428), .S(n372), .Y(n452) );
  MUX2X1 U397 ( .B(n454), .A(n455), .S(n370), .Y(n428) );
  MUX2X1 U398 ( .B(n456), .A(n457), .S(n369), .Y(n453) );
  MUX2X1 U399 ( .B(n458), .A(n380), .S(n378), .Y(B[29]) );
  MUX2X1 U400 ( .B(n409), .A(n380), .S(n378), .Y(B[28]) );
  MUX2X1 U401 ( .B(n408), .A(n380), .S(n378), .Y(B[27]) );
  MUX2X1 U402 ( .B(n459), .A(n380), .S(n378), .Y(B[26]) );
  MUX2X1 U403 ( .B(n412), .A(n380), .S(n378), .Y(B[25]) );
  MUX2X1 U404 ( .B(n460), .A(A[31]), .S(n375), .Y(n412) );
  MUX2X1 U405 ( .B(n405), .A(n380), .S(n378), .Y(B[24]) );
  MUX2X1 U406 ( .B(n462), .A(n380), .S(n375), .Y(n461) );
  MUX2X1 U407 ( .B(n404), .A(n380), .S(n378), .Y(B[23]) );
  MUX2X1 U408 ( .B(n464), .A(n380), .S(n375), .Y(n463) );
  MUX2X1 U409 ( .B(n425), .A(n380), .S(n378), .Y(B[22]) );
  MUX2X1 U410 ( .B(n465), .A(n466), .S(n375), .Y(n425) );
  MUX2X1 U411 ( .B(n431), .A(n380), .S(n378), .Y(B[21]) );
  MUX2X1 U412 ( .B(n402), .A(n467), .S(n375), .Y(n431) );
  MUX2X1 U413 ( .B(n401), .A(n380), .S(n378), .Y(B[20]) );
  MUX2X1 U414 ( .B(n469), .A(n470), .S(n375), .Y(n468) );
  MUX2X1 U415 ( .B(n382), .A(n471), .S(n377), .Y(B[1]) );
  MUX2X1 U416 ( .B(n473), .A(n414), .S(n375), .Y(n472) );
  MUX2X1 U417 ( .B(n434), .A(n474), .S(SH[2]), .Y(n414) );
  MUX2X1 U418 ( .B(n445), .A(n475), .S(SH[1]), .Y(n434) );
  MUX2X1 U419 ( .B(A[9]), .A(A[10]), .S(SH[0]), .Y(n445) );
  MUX2X1 U420 ( .B(n476), .A(n433), .S(n372), .Y(n473) );
  MUX2X1 U421 ( .B(n447), .A(n444), .S(SH[1]), .Y(n433) );
  MUX2X1 U422 ( .B(A[7]), .A(A[8]), .S(SH[0]), .Y(n444) );
  MUX2X1 U423 ( .B(A[5]), .A(A[6]), .S(SH[0]), .Y(n447) );
  MUX2X1 U424 ( .B(n477), .A(n446), .S(SH[1]), .Y(n476) );
  MUX2X1 U425 ( .B(A[3]), .A(A[4]), .S(SH[0]), .Y(n446) );
  MUX2X1 U426 ( .B(A[1]), .A(A[2]), .S(SH[0]), .Y(n477) );
  MUX2X1 U427 ( .B(n400), .A(n380), .S(n377), .Y(B[19]) );
  MUX2X1 U428 ( .B(n479), .A(n480), .S(n375), .Y(n478) );
  MUX2X1 U429 ( .B(n450), .A(n380), .S(n377), .Y(B[18]) );
  MUX2X1 U430 ( .B(n481), .A(n482), .S(n375), .Y(n450) );
  MUX2X1 U431 ( .B(n471), .A(n380), .S(n377), .Y(B[17]) );
  MUX2X1 U432 ( .B(n398), .A(n460), .S(n375), .Y(n471) );
  MUX2X1 U433 ( .B(n406), .A(n410), .S(n372), .Y(n460) );
  MUX2X1 U434 ( .B(n484), .A(n485), .S(n372), .Y(n415) );
  MUX2X1 U435 ( .B(n487), .A(A[31]), .S(n377), .Y(n486) );
  MUX2X1 U436 ( .B(n396), .A(n380), .S(n377), .Y(B[15]) );
  MUX2X1 U437 ( .B(n421), .A(n464), .S(n375), .Y(n488) );
  MUX2X1 U438 ( .B(n489), .A(n490), .S(n372), .Y(n464) );
  MUX2X1 U439 ( .B(n491), .A(n492), .S(n372), .Y(n421) );
  MUX2X1 U440 ( .B(n493), .A(n448), .S(n377), .Y(B[14]) );
  MUX2X1 U441 ( .B(n466), .A(A[31]), .S(n374), .Y(n448) );
  MUX2X1 U442 ( .B(n494), .A(n380), .S(n372), .Y(n466) );
  MUX2X1 U443 ( .B(n426), .A(n465), .S(n374), .Y(n493) );
  MUX2X1 U444 ( .B(n403), .A(n407), .S(n372), .Y(n465) );
  MUX2X1 U445 ( .B(n395), .A(n399), .S(n372), .Y(n426) );
  MUX2X1 U446 ( .B(n495), .A(n458), .S(n377), .Y(B[13]) );
  MUX2X1 U447 ( .B(n467), .A(A[31]), .S(n374), .Y(n458) );
  MUX2X1 U448 ( .B(n410), .A(n380), .S(n372), .Y(n467) );
  MUX2X1 U449 ( .B(n497), .A(n380), .S(n370), .Y(n496) );
  MUX2X1 U450 ( .B(n394), .A(n402), .S(n374), .Y(n495) );
  MUX2X1 U451 ( .B(n485), .A(n483), .S(n372), .Y(n498) );
  MUX2X1 U452 ( .B(n499), .A(n500), .S(n370), .Y(n483) );
  MUX2X1 U453 ( .B(n501), .A(n502), .S(n370), .Y(n485) );
  MUX2X1 U454 ( .B(n474), .A(n484), .S(n372), .Y(n503) );
  MUX2X1 U455 ( .B(n504), .A(n505), .S(n370), .Y(n484) );
  MUX2X1 U456 ( .B(n506), .A(n507), .S(n370), .Y(n474) );
  MUX2X1 U457 ( .B(n393), .A(n409), .S(n377), .Y(B[12]) );
  MUX2X1 U458 ( .B(n470), .A(n380), .S(n374), .Y(n508) );
  MUX2X1 U459 ( .B(n509), .A(A[31]), .S(n372), .Y(n470) );
  MUX2X1 U460 ( .B(n437), .A(n469), .S(n374), .Y(n510) );
  MUX2X1 U461 ( .B(n511), .A(n512), .S(SH[2]), .Y(n469) );
  MUX2X1 U462 ( .B(n513), .A(n514), .S(SH[2]), .Y(n437) );
  MUX2X1 U463 ( .B(n392), .A(n408), .S(n377), .Y(B[11]) );
  MUX2X1 U464 ( .B(n480), .A(n380), .S(n374), .Y(n515) );
  MUX2X1 U465 ( .B(n490), .A(A[31]), .S(SH[2]), .Y(n480) );
  MUX2X1 U466 ( .B(n500), .A(n497), .S(n370), .Y(n490) );
  MUX2X1 U467 ( .B(A[29]), .A(A[30]), .S(SH[0]), .Y(n497) );
  MUX2X1 U468 ( .B(A[27]), .A(A[28]), .S(SH[0]), .Y(n500) );
  MUX2X1 U469 ( .B(n442), .A(n479), .S(n374), .Y(n516) );
  MUX2X1 U470 ( .B(n492), .A(n489), .S(SH[2]), .Y(n479) );
  MUX2X1 U471 ( .B(n502), .A(n499), .S(n370), .Y(n489) );
  MUX2X1 U472 ( .B(A[25]), .A(A[26]), .S(SH[0]), .Y(n499) );
  MUX2X1 U473 ( .B(A[23]), .A(A[24]), .S(SH[0]), .Y(n502) );
  MUX2X1 U474 ( .B(n505), .A(n501), .S(n370), .Y(n492) );
  MUX2X1 U475 ( .B(A[21]), .A(A[22]), .S(SH[0]), .Y(n501) );
  MUX2X1 U476 ( .B(A[19]), .A(A[20]), .S(SH[0]), .Y(n505) );
  MUX2X1 U477 ( .B(n423), .A(n491), .S(SH[2]), .Y(n442) );
  MUX2X1 U478 ( .B(n507), .A(n504), .S(n370), .Y(n491) );
  MUX2X1 U479 ( .B(A[17]), .A(A[18]), .S(SH[0]), .Y(n504) );
  MUX2X1 U480 ( .B(A[15]), .A(A[16]), .S(SH[0]), .Y(n507) );
  MUX2X1 U481 ( .B(n475), .A(n506), .S(n370), .Y(n423) );
  MUX2X1 U482 ( .B(A[13]), .A(A[14]), .S(SH[0]), .Y(n506) );
  MUX2X1 U483 ( .B(A[11]), .A(A[12]), .S(SH[0]), .Y(n475) );
  MUX2X1 U484 ( .B(n517), .A(n459), .S(n377), .Y(B[10]) );
  MUX2X1 U485 ( .B(n482), .A(A[31]), .S(n374), .Y(n459) );
  MUX2X1 U486 ( .B(n407), .A(n494), .S(SH[2]), .Y(n482) );
  MUX2X1 U487 ( .B(n411), .A(A[31]), .S(n370), .Y(n494) );
  MUX2X1 U488 ( .B(n520), .A(n521), .S(n370), .Y(n519) );
  MUX2X1 U489 ( .B(n451), .A(n481), .S(n374), .Y(n517) );
  MUX2X1 U490 ( .B(n399), .A(n403), .S(n372), .Y(n481) );
  MUX2X1 U491 ( .B(n523), .A(n524), .S(n369), .Y(n522) );
  MUX2X1 U492 ( .B(n526), .A(n527), .S(n369), .Y(n525) );
  MUX2X1 U493 ( .B(n391), .A(n395), .S(SH[2]), .Y(n451) );
  MUX2X1 U494 ( .B(n529), .A(n530), .S(n369), .Y(n528) );
  MUX2X1 U495 ( .B(n531), .A(n532), .S(n369), .Y(n429) );
  MUX2X1 U496 ( .B(n534), .A(n487), .S(n377), .Y(n533) );
  MUX2X1 U497 ( .B(n418), .A(n462), .S(n374), .Y(n487) );
  MUX2X1 U498 ( .B(n512), .A(n509), .S(SH[2]), .Y(n462) );
  MUX2X1 U499 ( .B(n521), .A(n518), .S(n369), .Y(n509) );
  MUX2X1 U500 ( .B(A[30]), .A(A[31]), .S(SH[0]), .Y(n518) );
  MUX2X1 U501 ( .B(A[28]), .A(A[29]), .S(SH[0]), .Y(n521) );
  MUX2X1 U502 ( .B(n524), .A(n520), .S(n369), .Y(n512) );
  MUX2X1 U503 ( .B(A[26]), .A(A[27]), .S(SH[0]), .Y(n520) );
  MUX2X1 U504 ( .B(A[24]), .A(A[25]), .S(SH[0]), .Y(n524) );
  MUX2X1 U505 ( .B(n514), .A(n511), .S(SH[2]), .Y(n418) );
  MUX2X1 U506 ( .B(n527), .A(n523), .S(n369), .Y(n511) );
  MUX2X1 U507 ( .B(A[22]), .A(A[23]), .S(SH[0]), .Y(n523) );
  MUX2X1 U508 ( .B(A[20]), .A(A[21]), .S(SH[0]), .Y(n527) );
  MUX2X1 U509 ( .B(n530), .A(n526), .S(n369), .Y(n514) );
  MUX2X1 U510 ( .B(A[18]), .A(A[19]), .S(SH[0]), .Y(n526) );
  MUX2X1 U511 ( .B(A[16]), .A(A[17]), .S(SH[0]), .Y(n530) );
  MUX2X1 U512 ( .B(n535), .A(n417), .S(n374), .Y(n534) );
  MUX2X1 U513 ( .B(n439), .A(n513), .S(SH[2]), .Y(n417) );
  MUX2X1 U514 ( .B(n532), .A(n529), .S(n369), .Y(n513) );
  MUX2X1 U515 ( .B(A[14]), .A(A[15]), .S(SH[0]), .Y(n529) );
  MUX2X1 U516 ( .B(A[12]), .A(A[13]), .S(SH[0]), .Y(n532) );
  MUX2X1 U517 ( .B(n455), .A(n531), .S(n369), .Y(n439) );
  MUX2X1 U518 ( .B(A[10]), .A(A[11]), .S(SH[0]), .Y(n531) );
  MUX2X1 U519 ( .B(A[8]), .A(A[9]), .S(SH[0]), .Y(n455) );
  MUX2X1 U520 ( .B(n536), .A(n438), .S(SH[2]), .Y(n535) );
  MUX2X1 U521 ( .B(n457), .A(n454), .S(n369), .Y(n438) );
  MUX2X1 U522 ( .B(A[6]), .A(A[7]), .S(SH[0]), .Y(n454) );
  MUX2X1 U523 ( .B(A[4]), .A(A[5]), .S(SH[0]), .Y(n457) );
  MUX2X1 U524 ( .B(n537), .A(n456), .S(n369), .Y(n536) );
  MUX2X1 U525 ( .B(A[2]), .A(A[3]), .S(SH[0]), .Y(n456) );
  MUX2X1 U526 ( .B(A[0]), .A(A[1]), .S(SH[0]), .Y(n537) );
endmodule


module alu_DW_rightsh_15 ( A, DATA_TC, SH, B );
  input [63:0] A;
  input [5:0] SH;
  output [63:0] B;
  input DATA_TC;
  wire   n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209;

  INVX1 U790 ( .A(B[63]), .Y(n894) );
  INVX1 U791 ( .A(n893), .Y(n892) );
  INVX1 U792 ( .A(n893), .Y(B[63]) );
  INVX1 U793 ( .A(n867), .Y(n863) );
  INVX1 U794 ( .A(n867), .Y(n866) );
  INVX1 U795 ( .A(n867), .Y(n864) );
  INVX1 U796 ( .A(A[63]), .Y(n893) );
  INVX1 U797 ( .A(n881), .Y(n877) );
  INVX1 U798 ( .A(n881), .Y(n879) );
  INVX1 U799 ( .A(n881), .Y(n878) );
  INVX1 U800 ( .A(n881), .Y(n880) );
  INVX1 U801 ( .A(n876), .Y(n874) );
  INVX1 U802 ( .A(n876), .Y(n872) );
  INVX1 U803 ( .A(n876), .Y(n873) );
  INVX1 U804 ( .A(n876), .Y(n875) );
  INVX1 U805 ( .A(n871), .Y(n868) );
  INVX1 U806 ( .A(n871), .Y(n869) );
  INVX1 U807 ( .A(n871), .Y(n870) );
  INVX1 U808 ( .A(n867), .Y(n865) );
  INVX1 U809 ( .A(n885), .Y(n883) );
  INVX1 U810 ( .A(n885), .Y(n882) );
  INVX1 U811 ( .A(n885), .Y(n884) );
  INVX1 U812 ( .A(SH[0]), .Y(n867) );
  INVX1 U813 ( .A(SH[3]), .Y(n881) );
  INVX1 U814 ( .A(SH[2]), .Y(n876) );
  INVX1 U815 ( .A(SH[1]), .Y(n871) );
  INVX1 U816 ( .A(SH[4]), .Y(n885) );
  INVX1 U817 ( .A(n890), .Y(n886) );
  INVX1 U818 ( .A(n890), .Y(n888) );
  INVX1 U819 ( .A(n890), .Y(n887) );
  INVX1 U820 ( .A(n890), .Y(n889) );
  INVX1 U821 ( .A(SH[5]), .Y(n890) );
  MUX2X1 U822 ( .B(n895), .A(n896), .S(n889), .Y(B[9]) );
  MUX2X1 U823 ( .B(n897), .A(n898), .S(n883), .Y(n895) );
  MUX2X1 U824 ( .B(n899), .A(n900), .S(n877), .Y(n897) );
  MUX2X1 U825 ( .B(n901), .A(n902), .S(n886), .Y(B[8]) );
  MUX2X1 U826 ( .B(n903), .A(n904), .S(n883), .Y(n901) );
  MUX2X1 U827 ( .B(n905), .A(n906), .S(n879), .Y(n903) );
  MUX2X1 U828 ( .B(n907), .A(n908), .S(n887), .Y(B[7]) );
  MUX2X1 U829 ( .B(n909), .A(n910), .S(n883), .Y(n907) );
  MUX2X1 U830 ( .B(n911), .A(n912), .S(n880), .Y(n909) );
  MUX2X1 U831 ( .B(n913), .A(n914), .S(n873), .Y(n911) );
  MUX2X1 U832 ( .B(n915), .A(n916), .S(n889), .Y(B[6]) );
  MUX2X1 U833 ( .B(n917), .A(n918), .S(n884), .Y(n915) );
  MUX2X1 U834 ( .B(n919), .A(n920), .S(n880), .Y(n917) );
  MUX2X1 U835 ( .B(n921), .A(n922), .S(n872), .Y(n919) );
  MUX2X1 U836 ( .B(n923), .A(n894), .S(n889), .Y(B[62]) );
  MUX2X1 U837 ( .B(n924), .A(n894), .S(n889), .Y(B[61]) );
  MUX2X1 U838 ( .B(n925), .A(n894), .S(n889), .Y(B[60]) );
  MUX2X1 U839 ( .B(n926), .A(n927), .S(n889), .Y(B[5]) );
  MUX2X1 U840 ( .B(n928), .A(n929), .S(n884), .Y(n926) );
  MUX2X1 U841 ( .B(n930), .A(n931), .S(n880), .Y(n928) );
  MUX2X1 U842 ( .B(n932), .A(n933), .S(n873), .Y(n930) );
  MUX2X1 U843 ( .B(n934), .A(n894), .S(n889), .Y(B[59]) );
  MUX2X1 U844 ( .B(n935), .A(n894), .S(n889), .Y(B[58]) );
  MUX2X1 U845 ( .B(n936), .A(n894), .S(n889), .Y(B[57]) );
  MUX2X1 U846 ( .B(n937), .A(n894), .S(n889), .Y(B[56]) );
  MUX2X1 U847 ( .B(n938), .A(n894), .S(n889), .Y(B[55]) );
  MUX2X1 U848 ( .B(n939), .A(n894), .S(n889), .Y(B[54]) );
  MUX2X1 U849 ( .B(n940), .A(n894), .S(n889), .Y(B[53]) );
  MUX2X1 U850 ( .B(n941), .A(n894), .S(n888), .Y(B[52]) );
  MUX2X1 U851 ( .B(n942), .A(n894), .S(n888), .Y(B[51]) );
  MUX2X1 U852 ( .B(n943), .A(n893), .S(n888), .Y(B[50]) );
  MUX2X1 U853 ( .B(n944), .A(n945), .S(n888), .Y(B[4]) );
  MUX2X1 U854 ( .B(n946), .A(n947), .S(n884), .Y(n944) );
  MUX2X1 U855 ( .B(n948), .A(n949), .S(n880), .Y(n946) );
  MUX2X1 U856 ( .B(n950), .A(n951), .S(n875), .Y(n948) );
  MUX2X1 U857 ( .B(n952), .A(n893), .S(n888), .Y(B[49]) );
  MUX2X1 U858 ( .B(n953), .A(n893), .S(n888), .Y(B[48]) );
  MUX2X1 U859 ( .B(n954), .A(n893), .S(n888), .Y(B[47]) );
  MUX2X1 U860 ( .B(n955), .A(n893), .S(n888), .Y(B[46]) );
  MUX2X1 U861 ( .B(n956), .A(n893), .S(n888), .Y(B[45]) );
  MUX2X1 U862 ( .B(n957), .A(n893), .S(n888), .Y(B[44]) );
  MUX2X1 U863 ( .B(n958), .A(n893), .S(n888), .Y(B[43]) );
  MUX2X1 U864 ( .B(n959), .A(n893), .S(n888), .Y(B[42]) );
  MUX2X1 U865 ( .B(n896), .A(n893), .S(n887), .Y(B[41]) );
  MUX2X1 U866 ( .B(n960), .A(n961), .S(n884), .Y(n896) );
  MUX2X1 U867 ( .B(n902), .A(n893), .S(n887), .Y(B[40]) );
  MUX2X1 U868 ( .B(n962), .A(n963), .S(n884), .Y(n902) );
  MUX2X1 U869 ( .B(n964), .A(n965), .S(n887), .Y(B[3]) );
  MUX2X1 U870 ( .B(n966), .A(n967), .S(n884), .Y(n964) );
  MUX2X1 U871 ( .B(n968), .A(n969), .S(n880), .Y(n966) );
  MUX2X1 U872 ( .B(n970), .A(n913), .S(n875), .Y(n968) );
  MUX2X1 U873 ( .B(n971), .A(n972), .S(n870), .Y(n913) );
  MUX2X1 U874 ( .B(n973), .A(n974), .S(n870), .Y(n970) );
  MUX2X1 U875 ( .B(n908), .A(n893), .S(n887), .Y(B[39]) );
  MUX2X1 U876 ( .B(n975), .A(n976), .S(n884), .Y(n908) );
  MUX2X1 U877 ( .B(n916), .A(n893), .S(n887), .Y(B[38]) );
  MUX2X1 U878 ( .B(n977), .A(n978), .S(n884), .Y(n916) );
  MUX2X1 U879 ( .B(n927), .A(n893), .S(n887), .Y(B[37]) );
  MUX2X1 U880 ( .B(n979), .A(n980), .S(n884), .Y(n927) );
  MUX2X1 U881 ( .B(n945), .A(n894), .S(n887), .Y(B[36]) );
  MUX2X1 U882 ( .B(n981), .A(n982), .S(n884), .Y(n945) );
  MUX2X1 U883 ( .B(n965), .A(n893), .S(n887), .Y(B[35]) );
  MUX2X1 U884 ( .B(n983), .A(n984), .S(n884), .Y(n965) );
  MUX2X1 U885 ( .B(n985), .A(n893), .S(n887), .Y(B[34]) );
  MUX2X1 U886 ( .B(n986), .A(n893), .S(n887), .Y(B[33]) );
  MUX2X1 U887 ( .B(n987), .A(n893), .S(n887), .Y(B[32]) );
  MUX2X1 U888 ( .B(n988), .A(n894), .S(n887), .Y(B[31]) );
  MUX2X1 U889 ( .B(n989), .A(n990), .S(n884), .Y(n988) );
  MUX2X1 U890 ( .B(n991), .A(n923), .S(n886), .Y(B[30]) );
  MUX2X1 U891 ( .B(n992), .A(B[63]), .S(n883), .Y(n923) );
  MUX2X1 U892 ( .B(n993), .A(n994), .S(n883), .Y(n991) );
  MUX2X1 U893 ( .B(n995), .A(n985), .S(n886), .Y(B[2]) );
  MUX2X1 U894 ( .B(n996), .A(n997), .S(n883), .Y(n985) );
  MUX2X1 U895 ( .B(n998), .A(n999), .S(n883), .Y(n995) );
  MUX2X1 U896 ( .B(n1000), .A(n1001), .S(n880), .Y(n998) );
  MUX2X1 U897 ( .B(n1002), .A(n921), .S(n875), .Y(n1000) );
  MUX2X1 U898 ( .B(n1003), .A(n1004), .S(n870), .Y(n921) );
  MUX2X1 U899 ( .B(n1005), .A(n1006), .S(n870), .Y(n1002) );
  MUX2X1 U900 ( .B(n1007), .A(n924), .S(n886), .Y(B[29]) );
  MUX2X1 U901 ( .B(n1008), .A(B[63]), .S(n883), .Y(n924) );
  MUX2X1 U902 ( .B(n1009), .A(n1010), .S(n883), .Y(n1007) );
  MUX2X1 U903 ( .B(n1011), .A(n925), .S(n886), .Y(B[28]) );
  MUX2X1 U904 ( .B(n1012), .A(B[63]), .S(n883), .Y(n925) );
  MUX2X1 U905 ( .B(n1013), .A(n1014), .S(n883), .Y(n1011) );
  MUX2X1 U906 ( .B(n1015), .A(n934), .S(n886), .Y(B[27]) );
  MUX2X1 U907 ( .B(n1016), .A(B[63]), .S(n883), .Y(n934) );
  MUX2X1 U908 ( .B(n1017), .A(n1018), .S(n883), .Y(n1015) );
  MUX2X1 U909 ( .B(n1019), .A(n935), .S(n886), .Y(B[26]) );
  MUX2X1 U910 ( .B(n1020), .A(B[63]), .S(n883), .Y(n935) );
  MUX2X1 U911 ( .B(n1021), .A(n1022), .S(n883), .Y(n1019) );
  MUX2X1 U912 ( .B(n1023), .A(n936), .S(n886), .Y(B[25]) );
  MUX2X1 U913 ( .B(n961), .A(B[63]), .S(n882), .Y(n936) );
  MUX2X1 U914 ( .B(n1024), .A(n894), .S(n880), .Y(n961) );
  MUX2X1 U915 ( .B(n898), .A(n960), .S(n882), .Y(n1023) );
  MUX2X1 U916 ( .B(n1025), .A(n1026), .S(n880), .Y(n960) );
  MUX2X1 U917 ( .B(n1027), .A(n1028), .S(n880), .Y(n898) );
  MUX2X1 U918 ( .B(n1029), .A(n937), .S(n886), .Y(B[24]) );
  MUX2X1 U919 ( .B(n963), .A(B[63]), .S(n882), .Y(n937) );
  MUX2X1 U920 ( .B(n1030), .A(n894), .S(n880), .Y(n963) );
  MUX2X1 U921 ( .B(n904), .A(n962), .S(n882), .Y(n1029) );
  MUX2X1 U922 ( .B(n1031), .A(n1032), .S(n880), .Y(n962) );
  MUX2X1 U923 ( .B(n1033), .A(n1034), .S(n880), .Y(n904) );
  MUX2X1 U924 ( .B(n1035), .A(n938), .S(n886), .Y(B[23]) );
  MUX2X1 U925 ( .B(n976), .A(n892), .S(n882), .Y(n938) );
  MUX2X1 U926 ( .B(n1036), .A(n894), .S(n880), .Y(n976) );
  MUX2X1 U927 ( .B(n910), .A(n975), .S(n882), .Y(n1035) );
  MUX2X1 U928 ( .B(n1037), .A(n1038), .S(n879), .Y(n975) );
  MUX2X1 U929 ( .B(n1039), .A(n1040), .S(n879), .Y(n910) );
  MUX2X1 U930 ( .B(n1041), .A(n939), .S(n886), .Y(B[22]) );
  MUX2X1 U931 ( .B(n978), .A(n892), .S(n882), .Y(n939) );
  MUX2X1 U932 ( .B(n1042), .A(n1043), .S(n879), .Y(n978) );
  MUX2X1 U933 ( .B(n918), .A(n977), .S(n882), .Y(n1041) );
  MUX2X1 U934 ( .B(n1044), .A(n1045), .S(n879), .Y(n977) );
  MUX2X1 U935 ( .B(n1046), .A(n1047), .S(n879), .Y(n918) );
  MUX2X1 U936 ( .B(n1048), .A(n940), .S(n886), .Y(B[21]) );
  MUX2X1 U937 ( .B(n980), .A(n892), .S(n882), .Y(n940) );
  MUX2X1 U938 ( .B(n1049), .A(n1050), .S(n879), .Y(n980) );
  MUX2X1 U939 ( .B(n929), .A(n979), .S(n882), .Y(n1048) );
  MUX2X1 U940 ( .B(n1051), .A(n1052), .S(n879), .Y(n979) );
  MUX2X1 U941 ( .B(n1053), .A(n1054), .S(n879), .Y(n929) );
  MUX2X1 U942 ( .B(n1055), .A(n941), .S(n886), .Y(B[20]) );
  MUX2X1 U943 ( .B(n982), .A(n892), .S(n882), .Y(n941) );
  MUX2X1 U944 ( .B(n1056), .A(n1057), .S(n879), .Y(n982) );
  MUX2X1 U945 ( .B(n947), .A(n981), .S(n882), .Y(n1055) );
  MUX2X1 U946 ( .B(n1058), .A(n1059), .S(n879), .Y(n981) );
  MUX2X1 U947 ( .B(n1060), .A(n1061), .S(n879), .Y(n947) );
  MUX2X1 U948 ( .B(n1062), .A(n986), .S(n886), .Y(B[1]) );
  MUX2X1 U949 ( .B(n1063), .A(n1064), .S(SH[4]), .Y(n986) );
  MUX2X1 U950 ( .B(n1065), .A(n1066), .S(SH[4]), .Y(n1062) );
  MUX2X1 U951 ( .B(n1067), .A(n899), .S(n879), .Y(n1065) );
  MUX2X1 U952 ( .B(n933), .A(n1068), .S(n875), .Y(n899) );
  MUX2X1 U953 ( .B(n972), .A(n1069), .S(n870), .Y(n933) );
  MUX2X1 U954 ( .B(A[9]), .A(A[10]), .S(n865), .Y(n972) );
  MUX2X1 U955 ( .B(n1070), .A(n932), .S(n875), .Y(n1067) );
  MUX2X1 U956 ( .B(n974), .A(n971), .S(n870), .Y(n932) );
  MUX2X1 U957 ( .B(A[7]), .A(A[8]), .S(n865), .Y(n971) );
  MUX2X1 U958 ( .B(A[5]), .A(A[6]), .S(n865), .Y(n974) );
  MUX2X1 U959 ( .B(n1071), .A(n973), .S(n870), .Y(n1070) );
  MUX2X1 U960 ( .B(A[3]), .A(A[4]), .S(n866), .Y(n973) );
  MUX2X1 U961 ( .B(A[1]), .A(A[2]), .S(n866), .Y(n1071) );
  MUX2X1 U962 ( .B(n1072), .A(n942), .S(n889), .Y(B[19]) );
  MUX2X1 U963 ( .B(n984), .A(n892), .S(SH[4]), .Y(n942) );
  MUX2X1 U964 ( .B(n1073), .A(n1074), .S(n877), .Y(n984) );
  MUX2X1 U965 ( .B(n967), .A(n983), .S(SH[4]), .Y(n1072) );
  MUX2X1 U966 ( .B(n1075), .A(n1076), .S(n880), .Y(n983) );
  MUX2X1 U967 ( .B(n1077), .A(n1078), .S(n879), .Y(n967) );
  MUX2X1 U968 ( .B(n1079), .A(n943), .S(n889), .Y(B[18]) );
  MUX2X1 U969 ( .B(n997), .A(n892), .S(SH[4]), .Y(n943) );
  MUX2X1 U970 ( .B(n1080), .A(n1081), .S(n879), .Y(n997) );
  MUX2X1 U971 ( .B(n999), .A(n996), .S(SH[4]), .Y(n1079) );
  MUX2X1 U972 ( .B(n1082), .A(n1083), .S(n877), .Y(n996) );
  MUX2X1 U973 ( .B(n1084), .A(n1085), .S(n877), .Y(n999) );
  MUX2X1 U974 ( .B(n1086), .A(n952), .S(n886), .Y(B[17]) );
  MUX2X1 U975 ( .B(n1064), .A(n892), .S(SH[4]), .Y(n952) );
  MUX2X1 U976 ( .B(n1026), .A(n1024), .S(n879), .Y(n1064) );
  MUX2X1 U977 ( .B(n1087), .A(n1088), .S(n875), .Y(n1024) );
  MUX2X1 U978 ( .B(n1089), .A(n1090), .S(n875), .Y(n1026) );
  MUX2X1 U979 ( .B(n1066), .A(n1063), .S(SH[4]), .Y(n1086) );
  MUX2X1 U980 ( .B(n1028), .A(n1025), .S(n880), .Y(n1063) );
  MUX2X1 U981 ( .B(n1091), .A(n1092), .S(n875), .Y(n1025) );
  MUX2X1 U982 ( .B(n1093), .A(n1094), .S(n875), .Y(n1028) );
  MUX2X1 U983 ( .B(n900), .A(n1027), .S(n880), .Y(n1066) );
  MUX2X1 U984 ( .B(n1095), .A(n1096), .S(n875), .Y(n1027) );
  MUX2X1 U985 ( .B(n1097), .A(n1098), .S(n875), .Y(n900) );
  MUX2X1 U986 ( .B(n1099), .A(n953), .S(n886), .Y(B[16]) );
  MUX2X1 U987 ( .B(n1100), .A(n892), .S(n884), .Y(n953) );
  MUX2X1 U988 ( .B(n1101), .A(n1102), .S(SH[4]), .Y(n1099) );
  MUX2X1 U989 ( .B(n1103), .A(n954), .S(n889), .Y(B[15]) );
  MUX2X1 U990 ( .B(n990), .A(n892), .S(SH[4]), .Y(n954) );
  MUX2X1 U991 ( .B(n1038), .A(n1036), .S(SH[3]), .Y(n990) );
  MUX2X1 U992 ( .B(n1104), .A(n1105), .S(n875), .Y(n1036) );
  MUX2X1 U993 ( .B(n1106), .A(n1107), .S(n874), .Y(n1038) );
  MUX2X1 U994 ( .B(n1108), .A(n989), .S(n882), .Y(n1103) );
  MUX2X1 U995 ( .B(n1040), .A(n1037), .S(n879), .Y(n989) );
  MUX2X1 U996 ( .B(n1109), .A(n1110), .S(n874), .Y(n1037) );
  MUX2X1 U997 ( .B(n1111), .A(n1112), .S(n874), .Y(n1040) );
  MUX2X1 U998 ( .B(n912), .A(n1039), .S(n880), .Y(n1108) );
  MUX2X1 U999 ( .B(n1113), .A(n1114), .S(n874), .Y(n1039) );
  MUX2X1 U1000 ( .B(n1115), .A(n1116), .S(n874), .Y(n912) );
  MUX2X1 U1001 ( .B(n1117), .A(n955), .S(n887), .Y(B[14]) );
  MUX2X1 U1002 ( .B(n994), .A(n992), .S(n882), .Y(n955) );
  MUX2X1 U1003 ( .B(n1043), .A(n893), .S(n878), .Y(n992) );
  MUX2X1 U1004 ( .B(n1118), .A(n892), .S(n874), .Y(n1043) );
  MUX2X1 U1005 ( .B(n1045), .A(n1042), .S(n878), .Y(n994) );
  MUX2X1 U1006 ( .B(n1119), .A(n1120), .S(n874), .Y(n1042) );
  MUX2X1 U1007 ( .B(n1121), .A(n1122), .S(n874), .Y(n1045) );
  MUX2X1 U1008 ( .B(n1123), .A(n993), .S(n884), .Y(n1117) );
  MUX2X1 U1009 ( .B(n1047), .A(n1044), .S(n878), .Y(n993) );
  MUX2X1 U1010 ( .B(n1124), .A(n1125), .S(n874), .Y(n1044) );
  MUX2X1 U1011 ( .B(n1126), .A(n1127), .S(n874), .Y(n1047) );
  MUX2X1 U1012 ( .B(n920), .A(n1046), .S(n878), .Y(n1123) );
  MUX2X1 U1013 ( .B(n1128), .A(n1129), .S(n874), .Y(n1046) );
  MUX2X1 U1014 ( .B(n1130), .A(n1131), .S(n874), .Y(n920) );
  MUX2X1 U1015 ( .B(n1132), .A(n956), .S(n889), .Y(B[13]) );
  MUX2X1 U1016 ( .B(n1010), .A(n1008), .S(n882), .Y(n956) );
  MUX2X1 U1017 ( .B(n1050), .A(n894), .S(n878), .Y(n1008) );
  MUX2X1 U1018 ( .B(n1088), .A(B[63]), .S(n873), .Y(n1050) );
  MUX2X1 U1019 ( .B(n1133), .A(n894), .S(n870), .Y(n1088) );
  MUX2X1 U1020 ( .B(n1052), .A(n1049), .S(n878), .Y(n1010) );
  MUX2X1 U1021 ( .B(n1090), .A(n1087), .S(n873), .Y(n1049) );
  MUX2X1 U1022 ( .B(n1134), .A(n1135), .S(n870), .Y(n1087) );
  MUX2X1 U1023 ( .B(n1136), .A(n1137), .S(n870), .Y(n1090) );
  MUX2X1 U1024 ( .B(n1092), .A(n1089), .S(n873), .Y(n1052) );
  MUX2X1 U1025 ( .B(n1138), .A(n1139), .S(n870), .Y(n1089) );
  MUX2X1 U1026 ( .B(n1140), .A(n1141), .S(n870), .Y(n1092) );
  MUX2X1 U1027 ( .B(n1142), .A(n1009), .S(n883), .Y(n1132) );
  MUX2X1 U1028 ( .B(n1054), .A(n1051), .S(n878), .Y(n1009) );
  MUX2X1 U1029 ( .B(n1094), .A(n1091), .S(n873), .Y(n1051) );
  MUX2X1 U1030 ( .B(n1143), .A(n1144), .S(n870), .Y(n1091) );
  MUX2X1 U1031 ( .B(n1145), .A(n1146), .S(n870), .Y(n1094) );
  MUX2X1 U1032 ( .B(n1096), .A(n1093), .S(n873), .Y(n1054) );
  MUX2X1 U1033 ( .B(n1147), .A(n1148), .S(n870), .Y(n1093) );
  MUX2X1 U1034 ( .B(n1149), .A(n1150), .S(SH[1]), .Y(n1096) );
  MUX2X1 U1035 ( .B(n931), .A(n1053), .S(n878), .Y(n1142) );
  MUX2X1 U1036 ( .B(n1098), .A(n1095), .S(n873), .Y(n1053) );
  MUX2X1 U1037 ( .B(n1151), .A(n1152), .S(n869), .Y(n1095) );
  MUX2X1 U1038 ( .B(n1153), .A(n1154), .S(SH[1]), .Y(n1098) );
  MUX2X1 U1039 ( .B(n1068), .A(n1097), .S(n873), .Y(n931) );
  MUX2X1 U1040 ( .B(n1155), .A(n1156), .S(SH[1]), .Y(n1097) );
  MUX2X1 U1041 ( .B(n1157), .A(n1158), .S(SH[1]), .Y(n1068) );
  MUX2X1 U1042 ( .B(n1159), .A(n957), .S(n889), .Y(B[12]) );
  MUX2X1 U1043 ( .B(n1014), .A(n1012), .S(n883), .Y(n957) );
  MUX2X1 U1044 ( .B(n1057), .A(n894), .S(n878), .Y(n1012) );
  MUX2X1 U1045 ( .B(n1160), .A(B[63]), .S(n873), .Y(n1057) );
  MUX2X1 U1046 ( .B(n1059), .A(n1056), .S(n878), .Y(n1014) );
  MUX2X1 U1047 ( .B(n1161), .A(n1162), .S(n873), .Y(n1056) );
  MUX2X1 U1048 ( .B(n1163), .A(n1164), .S(n873), .Y(n1059) );
  MUX2X1 U1049 ( .B(n1165), .A(n1013), .S(n883), .Y(n1159) );
  MUX2X1 U1050 ( .B(n1061), .A(n1058), .S(n878), .Y(n1013) );
  MUX2X1 U1051 ( .B(n1166), .A(n1167), .S(n873), .Y(n1058) );
  MUX2X1 U1052 ( .B(n1168), .A(n1169), .S(n873), .Y(n1061) );
  MUX2X1 U1053 ( .B(n949), .A(n1060), .S(n878), .Y(n1165) );
  MUX2X1 U1054 ( .B(n1170), .A(n1171), .S(n872), .Y(n1060) );
  MUX2X1 U1055 ( .B(n1172), .A(n1173), .S(n872), .Y(n949) );
  MUX2X1 U1056 ( .B(n1174), .A(n958), .S(n886), .Y(B[11]) );
  MUX2X1 U1057 ( .B(n1018), .A(n1016), .S(n883), .Y(n958) );
  MUX2X1 U1058 ( .B(n1074), .A(n894), .S(n877), .Y(n1016) );
  MUX2X1 U1059 ( .B(n1105), .A(B[63]), .S(n872), .Y(n1074) );
  MUX2X1 U1060 ( .B(n1135), .A(n1133), .S(SH[1]), .Y(n1105) );
  MUX2X1 U1061 ( .B(A[61]), .A(A[62]), .S(n866), .Y(n1133) );
  MUX2X1 U1062 ( .B(A[59]), .A(A[60]), .S(n866), .Y(n1135) );
  MUX2X1 U1063 ( .B(n1076), .A(n1073), .S(n877), .Y(n1018) );
  MUX2X1 U1064 ( .B(n1107), .A(n1104), .S(n872), .Y(n1073) );
  MUX2X1 U1065 ( .B(n1137), .A(n1134), .S(SH[1]), .Y(n1104) );
  MUX2X1 U1066 ( .B(A[57]), .A(A[58]), .S(n866), .Y(n1134) );
  MUX2X1 U1067 ( .B(A[55]), .A(A[56]), .S(n866), .Y(n1137) );
  MUX2X1 U1068 ( .B(n1139), .A(n1136), .S(SH[1]), .Y(n1107) );
  MUX2X1 U1069 ( .B(A[53]), .A(A[54]), .S(n866), .Y(n1136) );
  MUX2X1 U1070 ( .B(A[51]), .A(A[52]), .S(n866), .Y(n1139) );
  MUX2X1 U1071 ( .B(n1110), .A(n1106), .S(n872), .Y(n1076) );
  MUX2X1 U1072 ( .B(n1141), .A(n1138), .S(SH[1]), .Y(n1106) );
  MUX2X1 U1073 ( .B(A[49]), .A(A[50]), .S(n866), .Y(n1138) );
  MUX2X1 U1074 ( .B(A[47]), .A(A[48]), .S(n866), .Y(n1141) );
  MUX2X1 U1075 ( .B(n1144), .A(n1140), .S(n869), .Y(n1110) );
  MUX2X1 U1076 ( .B(A[45]), .A(A[46]), .S(n866), .Y(n1140) );
  MUX2X1 U1077 ( .B(A[43]), .A(A[44]), .S(n866), .Y(n1144) );
  MUX2X1 U1078 ( .B(n1175), .A(n1017), .S(n883), .Y(n1174) );
  MUX2X1 U1079 ( .B(n1078), .A(n1075), .S(n877), .Y(n1017) );
  MUX2X1 U1080 ( .B(n1112), .A(n1109), .S(n872), .Y(n1075) );
  MUX2X1 U1081 ( .B(n1146), .A(n1143), .S(n868), .Y(n1109) );
  MUX2X1 U1082 ( .B(A[41]), .A(A[42]), .S(n865), .Y(n1143) );
  MUX2X1 U1083 ( .B(A[39]), .A(A[40]), .S(n865), .Y(n1146) );
  MUX2X1 U1084 ( .B(n1148), .A(n1145), .S(n868), .Y(n1112) );
  MUX2X1 U1085 ( .B(A[37]), .A(A[38]), .S(n865), .Y(n1145) );
  MUX2X1 U1086 ( .B(A[35]), .A(A[36]), .S(n865), .Y(n1148) );
  MUX2X1 U1087 ( .B(n1114), .A(n1111), .S(n872), .Y(n1078) );
  MUX2X1 U1088 ( .B(n1150), .A(n1147), .S(n869), .Y(n1111) );
  MUX2X1 U1089 ( .B(A[33]), .A(A[34]), .S(n865), .Y(n1147) );
  MUX2X1 U1090 ( .B(A[31]), .A(A[32]), .S(n865), .Y(n1150) );
  MUX2X1 U1091 ( .B(n1152), .A(n1149), .S(n869), .Y(n1114) );
  MUX2X1 U1092 ( .B(A[29]), .A(A[30]), .S(n865), .Y(n1149) );
  MUX2X1 U1093 ( .B(A[27]), .A(A[28]), .S(n865), .Y(n1152) );
  MUX2X1 U1094 ( .B(n969), .A(n1077), .S(n877), .Y(n1175) );
  MUX2X1 U1095 ( .B(n1116), .A(n1113), .S(n872), .Y(n1077) );
  MUX2X1 U1096 ( .B(n1154), .A(n1151), .S(n869), .Y(n1113) );
  MUX2X1 U1097 ( .B(A[25]), .A(A[26]), .S(n865), .Y(n1151) );
  MUX2X1 U1098 ( .B(A[23]), .A(A[24]), .S(n865), .Y(n1154) );
  MUX2X1 U1099 ( .B(n1156), .A(n1153), .S(n869), .Y(n1116) );
  MUX2X1 U1100 ( .B(A[21]), .A(A[22]), .S(n865), .Y(n1153) );
  MUX2X1 U1101 ( .B(A[19]), .A(A[20]), .S(n865), .Y(n1156) );
  MUX2X1 U1102 ( .B(n914), .A(n1115), .S(n872), .Y(n969) );
  MUX2X1 U1103 ( .B(n1158), .A(n1155), .S(n869), .Y(n1115) );
  MUX2X1 U1104 ( .B(A[17]), .A(A[18]), .S(n864), .Y(n1155) );
  MUX2X1 U1105 ( .B(A[15]), .A(A[16]), .S(n864), .Y(n1158) );
  MUX2X1 U1106 ( .B(n1069), .A(n1157), .S(n869), .Y(n914) );
  MUX2X1 U1107 ( .B(A[13]), .A(A[14]), .S(n864), .Y(n1157) );
  MUX2X1 U1108 ( .B(A[11]), .A(A[12]), .S(n864), .Y(n1069) );
  MUX2X1 U1109 ( .B(n1176), .A(n959), .S(n886), .Y(B[10]) );
  MUX2X1 U1110 ( .B(n1022), .A(n1020), .S(n884), .Y(n959) );
  MUX2X1 U1111 ( .B(n1081), .A(n894), .S(n877), .Y(n1020) );
  MUX2X1 U1112 ( .B(n1120), .A(n1118), .S(n872), .Y(n1081) );
  MUX2X1 U1113 ( .B(n1177), .A(n893), .S(n869), .Y(n1118) );
  MUX2X1 U1114 ( .B(n1178), .A(n1179), .S(n869), .Y(n1120) );
  MUX2X1 U1115 ( .B(n1083), .A(n1080), .S(n877), .Y(n1022) );
  MUX2X1 U1116 ( .B(n1122), .A(n1119), .S(n872), .Y(n1080) );
  MUX2X1 U1117 ( .B(n1180), .A(n1181), .S(n869), .Y(n1119) );
  MUX2X1 U1118 ( .B(n1182), .A(n1183), .S(n869), .Y(n1122) );
  MUX2X1 U1119 ( .B(n1125), .A(n1121), .S(n872), .Y(n1083) );
  MUX2X1 U1120 ( .B(n1184), .A(n1185), .S(n869), .Y(n1121) );
  MUX2X1 U1121 ( .B(n1186), .A(n1187), .S(n869), .Y(n1125) );
  MUX2X1 U1122 ( .B(n1188), .A(n1021), .S(n884), .Y(n1176) );
  MUX2X1 U1123 ( .B(n1085), .A(n1082), .S(n877), .Y(n1021) );
  MUX2X1 U1124 ( .B(n1127), .A(n1124), .S(n873), .Y(n1082) );
  MUX2X1 U1125 ( .B(n1189), .A(n1190), .S(n868), .Y(n1124) );
  MUX2X1 U1126 ( .B(n1191), .A(n1192), .S(n868), .Y(n1127) );
  MUX2X1 U1127 ( .B(n1129), .A(n1126), .S(n872), .Y(n1085) );
  MUX2X1 U1128 ( .B(n1193), .A(n1194), .S(n868), .Y(n1126) );
  MUX2X1 U1129 ( .B(n1195), .A(n1196), .S(n868), .Y(n1129) );
  MUX2X1 U1130 ( .B(n1001), .A(n1084), .S(n877), .Y(n1188) );
  MUX2X1 U1131 ( .B(n1131), .A(n1128), .S(n873), .Y(n1084) );
  MUX2X1 U1132 ( .B(n1197), .A(n1198), .S(n868), .Y(n1128) );
  MUX2X1 U1133 ( .B(n1199), .A(n1200), .S(n868), .Y(n1131) );
  MUX2X1 U1134 ( .B(n922), .A(n1130), .S(n872), .Y(n1001) );
  MUX2X1 U1135 ( .B(n1201), .A(n1202), .S(n868), .Y(n1130) );
  MUX2X1 U1136 ( .B(n1203), .A(n1204), .S(n868), .Y(n922) );
  MUX2X1 U1137 ( .B(n1205), .A(n987), .S(n886), .Y(B[0]) );
  MUX2X1 U1138 ( .B(n1102), .A(n1100), .S(n883), .Y(n987) );
  MUX2X1 U1139 ( .B(n1032), .A(n1030), .S(n877), .Y(n1100) );
  MUX2X1 U1140 ( .B(n1162), .A(n1160), .S(n873), .Y(n1030) );
  MUX2X1 U1141 ( .B(n1179), .A(n1177), .S(n868), .Y(n1160) );
  MUX2X1 U1142 ( .B(A[62]), .A(n892), .S(n864), .Y(n1177) );
  MUX2X1 U1143 ( .B(A[60]), .A(A[61]), .S(n864), .Y(n1179) );
  MUX2X1 U1144 ( .B(n1181), .A(n1178), .S(n868), .Y(n1162) );
  MUX2X1 U1145 ( .B(A[58]), .A(A[59]), .S(n864), .Y(n1178) );
  MUX2X1 U1146 ( .B(A[56]), .A(A[57]), .S(n864), .Y(n1181) );
  MUX2X1 U1147 ( .B(n1164), .A(n1161), .S(n873), .Y(n1032) );
  MUX2X1 U1148 ( .B(n1183), .A(n1180), .S(n868), .Y(n1161) );
  MUX2X1 U1149 ( .B(A[54]), .A(A[55]), .S(n864), .Y(n1180) );
  MUX2X1 U1150 ( .B(A[52]), .A(A[53]), .S(n864), .Y(n1183) );
  MUX2X1 U1151 ( .B(n1185), .A(n1182), .S(n868), .Y(n1164) );
  MUX2X1 U1152 ( .B(A[50]), .A(A[51]), .S(n864), .Y(n1182) );
  MUX2X1 U1153 ( .B(A[48]), .A(A[49]), .S(n864), .Y(n1185) );
  MUX2X1 U1154 ( .B(n1034), .A(n1031), .S(n877), .Y(n1102) );
  MUX2X1 U1155 ( .B(n1167), .A(n1163), .S(n872), .Y(n1031) );
  MUX2X1 U1156 ( .B(n1187), .A(n1184), .S(n870), .Y(n1163) );
  MUX2X1 U1157 ( .B(A[46]), .A(A[47]), .S(n863), .Y(n1184) );
  MUX2X1 U1158 ( .B(A[44]), .A(A[45]), .S(n863), .Y(n1187) );
  MUX2X1 U1159 ( .B(n1190), .A(n1186), .S(n870), .Y(n1167) );
  MUX2X1 U1160 ( .B(A[42]), .A(A[43]), .S(n863), .Y(n1186) );
  MUX2X1 U1161 ( .B(A[40]), .A(A[41]), .S(n863), .Y(n1190) );
  MUX2X1 U1162 ( .B(n1169), .A(n1166), .S(n872), .Y(n1034) );
  MUX2X1 U1163 ( .B(n1192), .A(n1189), .S(n870), .Y(n1166) );
  MUX2X1 U1164 ( .B(A[38]), .A(A[39]), .S(n863), .Y(n1189) );
  MUX2X1 U1165 ( .B(A[36]), .A(A[37]), .S(n863), .Y(n1192) );
  MUX2X1 U1166 ( .B(n1194), .A(n1191), .S(n870), .Y(n1169) );
  MUX2X1 U1167 ( .B(A[34]), .A(A[35]), .S(n863), .Y(n1191) );
  MUX2X1 U1168 ( .B(A[32]), .A(A[33]), .S(n863), .Y(n1194) );
  MUX2X1 U1169 ( .B(n1206), .A(n1101), .S(n883), .Y(n1205) );
  MUX2X1 U1170 ( .B(n906), .A(n1033), .S(n877), .Y(n1101) );
  MUX2X1 U1171 ( .B(n1171), .A(n1168), .S(n873), .Y(n1033) );
  MUX2X1 U1172 ( .B(n1196), .A(n1193), .S(n870), .Y(n1168) );
  MUX2X1 U1173 ( .B(A[30]), .A(A[31]), .S(n863), .Y(n1193) );
  MUX2X1 U1174 ( .B(A[28]), .A(A[29]), .S(n863), .Y(n1196) );
  MUX2X1 U1175 ( .B(n1198), .A(n1195), .S(n868), .Y(n1171) );
  MUX2X1 U1176 ( .B(A[26]), .A(A[27]), .S(n863), .Y(n1195) );
  MUX2X1 U1177 ( .B(A[24]), .A(A[25]), .S(n863), .Y(n1198) );
  MUX2X1 U1178 ( .B(n1173), .A(n1170), .S(n872), .Y(n906) );
  MUX2X1 U1179 ( .B(n1200), .A(n1197), .S(n868), .Y(n1170) );
  MUX2X1 U1180 ( .B(A[22]), .A(A[23]), .S(n863), .Y(n1197) );
  MUX2X1 U1181 ( .B(A[20]), .A(A[21]), .S(n865), .Y(n1200) );
  MUX2X1 U1182 ( .B(n1202), .A(n1199), .S(n868), .Y(n1173) );
  MUX2X1 U1183 ( .B(A[18]), .A(A[19]), .S(n864), .Y(n1199) );
  MUX2X1 U1184 ( .B(A[16]), .A(A[17]), .S(n864), .Y(n1202) );
  MUX2X1 U1185 ( .B(n1207), .A(n905), .S(n877), .Y(n1206) );
  MUX2X1 U1186 ( .B(n951), .A(n1172), .S(n873), .Y(n905) );
  MUX2X1 U1187 ( .B(n1204), .A(n1201), .S(n870), .Y(n1172) );
  MUX2X1 U1188 ( .B(A[14]), .A(A[15]), .S(n863), .Y(n1201) );
  MUX2X1 U1189 ( .B(A[12]), .A(A[13]), .S(n864), .Y(n1204) );
  MUX2X1 U1190 ( .B(n1004), .A(n1203), .S(n869), .Y(n951) );
  MUX2X1 U1191 ( .B(A[10]), .A(A[11]), .S(n863), .Y(n1203) );
  MUX2X1 U1192 ( .B(A[8]), .A(A[9]), .S(n865), .Y(n1004) );
  MUX2X1 U1193 ( .B(n1208), .A(n950), .S(n872), .Y(n1207) );
  MUX2X1 U1194 ( .B(n1006), .A(n1003), .S(n870), .Y(n950) );
  MUX2X1 U1195 ( .B(A[6]), .A(A[7]), .S(n863), .Y(n1003) );
  MUX2X1 U1196 ( .B(A[4]), .A(A[5]), .S(n865), .Y(n1006) );
  MUX2X1 U1197 ( .B(n1209), .A(n1005), .S(n869), .Y(n1208) );
  MUX2X1 U1198 ( .B(A[2]), .A(A[3]), .S(n864), .Y(n1005) );
  MUX2X1 U1199 ( .B(A[0]), .A(A[1]), .S(n863), .Y(n1209) );
endmodule


module alu_DW_rightsh_16 ( A, DATA_TC, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC;
  wire   n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544;
  assign B[31] = A[31];

  INVX1 U329 ( .A(n525), .Y(n408) );
  INVX1 U330 ( .A(n436), .Y(n416) );
  INVX1 U331 ( .A(n490), .Y(n399) );
  INVX1 U332 ( .A(n422), .Y(n401) );
  INVX1 U333 ( .A(n468), .Y(n405) );
  INVX1 U334 ( .A(n470), .Y(n396) );
  INVX1 U335 ( .A(n434), .Y(n417) );
  INVX1 U336 ( .A(n485), .Y(n394) );
  INVX1 U337 ( .A(n515), .Y(n406) );
  INVX1 U338 ( .A(n522), .Y(n393) );
  INVX1 U339 ( .A(n505), .Y(n398) );
  INVX1 U340 ( .A(n510), .Y(n402) );
  INVX1 U341 ( .A(n475), .Y(n407) );
  INVX1 U342 ( .A(n439), .Y(n390) );
  INVX1 U343 ( .A(A[31]), .Y(n387) );
  INVX1 U344 ( .A(n493), .Y(B[16]) );
  INVX1 U345 ( .A(n540), .Y(B[0]) );
  INVX1 U346 ( .A(n459), .Y(n418) );
  INVX1 U347 ( .A(n379), .Y(n376) );
  INVX1 U348 ( .A(n379), .Y(n377) );
  INVX1 U349 ( .A(n382), .Y(n380) );
  INVX1 U350 ( .A(n382), .Y(n381) );
  INVX1 U351 ( .A(n375), .Y(n373) );
  INVX1 U352 ( .A(n375), .Y(n372) );
  INVX1 U353 ( .A(n371), .Y(n369) );
  INVX1 U354 ( .A(n386), .Y(n384) );
  INVX1 U355 ( .A(n386), .Y(n383) );
  INVX1 U356 ( .A(n503), .Y(n397) );
  INVX1 U357 ( .A(n535), .Y(n415) );
  INVX1 U358 ( .A(n532), .Y(n413) );
  INVX1 U359 ( .A(n526), .Y(n409) );
  INVX1 U360 ( .A(n529), .Y(n411) );
  INVX1 U361 ( .A(n479), .Y(n388) );
  INVX1 U362 ( .A(n379), .Y(n378) );
  INVX1 U363 ( .A(n375), .Y(n374) );
  INVX1 U364 ( .A(n371), .Y(n370) );
  INVX1 U365 ( .A(n386), .Y(n385) );
  INVX1 U366 ( .A(n420), .Y(n389) );
  INVX1 U367 ( .A(n423), .Y(n412) );
  INVX1 U368 ( .A(n447), .Y(n391) );
  INVX1 U369 ( .A(n495), .Y(n395) );
  INVX1 U370 ( .A(n517), .Y(n410) );
  INVX1 U371 ( .A(n523), .Y(n400) );
  INVX1 U372 ( .A(n426), .Y(n392) );
  INVX1 U373 ( .A(n442), .Y(n414) );
  INVX1 U374 ( .A(SH[2]), .Y(n379) );
  INVX1 U375 ( .A(SH[3]), .Y(n382) );
  INVX1 U376 ( .A(SH[1]), .Y(n375) );
  INVX1 U377 ( .A(SH[0]), .Y(n371) );
  INVX1 U378 ( .A(SH[4]), .Y(n386) );
  MUX2X1 U379 ( .B(n389), .A(n419), .S(n385), .Y(B[9]) );
  MUX2X1 U380 ( .B(n421), .A(n422), .S(SH[3]), .Y(n420) );
  MUX2X1 U381 ( .B(n412), .A(n405), .S(n385), .Y(B[8]) );
  MUX2X1 U382 ( .B(n424), .A(n425), .S(SH[3]), .Y(n423) );
  MUX2X1 U383 ( .B(n392), .A(n396), .S(n385), .Y(B[7]) );
  MUX2X1 U384 ( .B(n427), .A(n428), .S(SH[3]), .Y(n426) );
  MUX2X1 U385 ( .B(n429), .A(n430), .S(n378), .Y(n427) );
  MUX2X1 U386 ( .B(n431), .A(n432), .S(n385), .Y(B[6]) );
  MUX2X1 U387 ( .B(n417), .A(n433), .S(n380), .Y(n431) );
  MUX2X1 U388 ( .B(n435), .A(n436), .S(n378), .Y(n434) );
  MUX2X1 U389 ( .B(n437), .A(n438), .S(n385), .Y(B[5]) );
  MUX2X1 U390 ( .B(n390), .A(n402), .S(n380), .Y(n437) );
  MUX2X1 U391 ( .B(n440), .A(n441), .S(n378), .Y(n439) );
  MUX2X1 U392 ( .B(n414), .A(n407), .S(n385), .Y(B[4]) );
  MUX2X1 U393 ( .B(n443), .A(n444), .S(SH[3]), .Y(n442) );
  MUX2X1 U394 ( .B(n445), .A(n446), .S(n378), .Y(n443) );
  MUX2X1 U395 ( .B(n391), .A(n394), .S(n385), .Y(B[3]) );
  MUX2X1 U396 ( .B(n448), .A(n449), .S(SH[3]), .Y(n447) );
  MUX2X1 U397 ( .B(n450), .A(n429), .S(n378), .Y(n448) );
  MUX2X1 U398 ( .B(n451), .A(n452), .S(n374), .Y(n429) );
  MUX2X1 U399 ( .B(n453), .A(n454), .S(n374), .Y(n450) );
  MUX2X1 U400 ( .B(n455), .A(n387), .S(n384), .Y(B[30]) );
  MUX2X1 U401 ( .B(n456), .A(n457), .S(n384), .Y(B[2]) );
  MUX2X1 U402 ( .B(n418), .A(n458), .S(n381), .Y(n456) );
  MUX2X1 U403 ( .B(n460), .A(n435), .S(n378), .Y(n459) );
  MUX2X1 U404 ( .B(n461), .A(n462), .S(n374), .Y(n435) );
  MUX2X1 U405 ( .B(n463), .A(n464), .S(n374), .Y(n460) );
  MUX2X1 U406 ( .B(n465), .A(n387), .S(n384), .Y(B[29]) );
  MUX2X1 U407 ( .B(n406), .A(n387), .S(n384), .Y(B[28]) );
  MUX2X1 U408 ( .B(n393), .A(n387), .S(n384), .Y(B[27]) );
  MUX2X1 U409 ( .B(n466), .A(n387), .S(n384), .Y(B[26]) );
  MUX2X1 U410 ( .B(n419), .A(n387), .S(n384), .Y(B[25]) );
  MUX2X1 U411 ( .B(n467), .A(A[31]), .S(n381), .Y(n419) );
  MUX2X1 U412 ( .B(n405), .A(n387), .S(n384), .Y(B[24]) );
  MUX2X1 U413 ( .B(n469), .A(n387), .S(n381), .Y(n468) );
  MUX2X1 U414 ( .B(n396), .A(n387), .S(n384), .Y(B[23]) );
  MUX2X1 U415 ( .B(n471), .A(n387), .S(n381), .Y(n470) );
  MUX2X1 U416 ( .B(n432), .A(n387), .S(n384), .Y(B[22]) );
  MUX2X1 U417 ( .B(n472), .A(n473), .S(n381), .Y(n432) );
  MUX2X1 U418 ( .B(n438), .A(n387), .S(n384), .Y(B[21]) );
  MUX2X1 U419 ( .B(n398), .A(n474), .S(n381), .Y(n438) );
  MUX2X1 U420 ( .B(n407), .A(n387), .S(n384), .Y(B[20]) );
  MUX2X1 U421 ( .B(n476), .A(n477), .S(n381), .Y(n475) );
  MUX2X1 U422 ( .B(n388), .A(n478), .S(n383), .Y(B[1]) );
  MUX2X1 U423 ( .B(n480), .A(n421), .S(n381), .Y(n479) );
  MUX2X1 U424 ( .B(n441), .A(n481), .S(n378), .Y(n421) );
  MUX2X1 U425 ( .B(n452), .A(n482), .S(n374), .Y(n441) );
  MUX2X1 U426 ( .B(A[9]), .A(A[10]), .S(n370), .Y(n452) );
  MUX2X1 U427 ( .B(n483), .A(n440), .S(n377), .Y(n480) );
  MUX2X1 U428 ( .B(n454), .A(n451), .S(n374), .Y(n440) );
  MUX2X1 U429 ( .B(A[7]), .A(A[8]), .S(n370), .Y(n451) );
  MUX2X1 U430 ( .B(A[5]), .A(A[6]), .S(n370), .Y(n454) );
  MUX2X1 U431 ( .B(n484), .A(n453), .S(n374), .Y(n483) );
  MUX2X1 U432 ( .B(A[3]), .A(A[4]), .S(n370), .Y(n453) );
  MUX2X1 U433 ( .B(A[1]), .A(A[2]), .S(n370), .Y(n484) );
  MUX2X1 U434 ( .B(n394), .A(n387), .S(n383), .Y(B[19]) );
  MUX2X1 U435 ( .B(n486), .A(n487), .S(n381), .Y(n485) );
  MUX2X1 U436 ( .B(n457), .A(n387), .S(n383), .Y(B[18]) );
  MUX2X1 U437 ( .B(n488), .A(n489), .S(n381), .Y(n457) );
  MUX2X1 U438 ( .B(n478), .A(n387), .S(n383), .Y(B[17]) );
  MUX2X1 U439 ( .B(n401), .A(n467), .S(n381), .Y(n478) );
  MUX2X1 U440 ( .B(n399), .A(n397), .S(n377), .Y(n467) );
  MUX2X1 U441 ( .B(n491), .A(n492), .S(n377), .Y(n422) );
  MUX2X1 U442 ( .B(n494), .A(A[31]), .S(n383), .Y(n493) );
  MUX2X1 U443 ( .B(n395), .A(n387), .S(n383), .Y(B[15]) );
  MUX2X1 U444 ( .B(n428), .A(n471), .S(n381), .Y(n495) );
  MUX2X1 U445 ( .B(n496), .A(n497), .S(n377), .Y(n471) );
  MUX2X1 U446 ( .B(n498), .A(n499), .S(n377), .Y(n428) );
  MUX2X1 U447 ( .B(n500), .A(n455), .S(n383), .Y(B[14]) );
  MUX2X1 U448 ( .B(n473), .A(A[31]), .S(n380), .Y(n455) );
  MUX2X1 U449 ( .B(n501), .A(n387), .S(n377), .Y(n473) );
  MUX2X1 U450 ( .B(n433), .A(n472), .S(n380), .Y(n500) );
  MUX2X1 U451 ( .B(n411), .A(n409), .S(n377), .Y(n472) );
  MUX2X1 U452 ( .B(n415), .A(n413), .S(n377), .Y(n433) );
  MUX2X1 U453 ( .B(n502), .A(n465), .S(n383), .Y(B[13]) );
  MUX2X1 U454 ( .B(n474), .A(A[31]), .S(n380), .Y(n465) );
  MUX2X1 U455 ( .B(n397), .A(n387), .S(n377), .Y(n474) );
  MUX2X1 U456 ( .B(n504), .A(n387), .S(n373), .Y(n503) );
  MUX2X1 U457 ( .B(n402), .A(n398), .S(n380), .Y(n502) );
  MUX2X1 U458 ( .B(n492), .A(n490), .S(n377), .Y(n505) );
  MUX2X1 U459 ( .B(n506), .A(n507), .S(n373), .Y(n490) );
  MUX2X1 U460 ( .B(n508), .A(n509), .S(n373), .Y(n492) );
  MUX2X1 U461 ( .B(n481), .A(n491), .S(n377), .Y(n510) );
  MUX2X1 U462 ( .B(n511), .A(n512), .S(n373), .Y(n491) );
  MUX2X1 U463 ( .B(n513), .A(n514), .S(n373), .Y(n481) );
  MUX2X1 U464 ( .B(n410), .A(n406), .S(n383), .Y(B[12]) );
  MUX2X1 U465 ( .B(n477), .A(n387), .S(n380), .Y(n515) );
  MUX2X1 U466 ( .B(n516), .A(A[31]), .S(n377), .Y(n477) );
  MUX2X1 U467 ( .B(n444), .A(n476), .S(n380), .Y(n517) );
  MUX2X1 U468 ( .B(n518), .A(n519), .S(n376), .Y(n476) );
  MUX2X1 U469 ( .B(n520), .A(n521), .S(n376), .Y(n444) );
  MUX2X1 U470 ( .B(n400), .A(n393), .S(n383), .Y(B[11]) );
  MUX2X1 U471 ( .B(n487), .A(n387), .S(n380), .Y(n522) );
  MUX2X1 U472 ( .B(n497), .A(A[31]), .S(n376), .Y(n487) );
  MUX2X1 U473 ( .B(n507), .A(n504), .S(n373), .Y(n497) );
  MUX2X1 U474 ( .B(A[29]), .A(A[30]), .S(n370), .Y(n504) );
  MUX2X1 U475 ( .B(A[27]), .A(A[28]), .S(n370), .Y(n507) );
  MUX2X1 U476 ( .B(n449), .A(n486), .S(n380), .Y(n523) );
  MUX2X1 U477 ( .B(n499), .A(n496), .S(n376), .Y(n486) );
  MUX2X1 U478 ( .B(n509), .A(n506), .S(n373), .Y(n496) );
  MUX2X1 U479 ( .B(A[25]), .A(A[26]), .S(SH[0]), .Y(n506) );
  MUX2X1 U480 ( .B(A[23]), .A(A[24]), .S(SH[0]), .Y(n509) );
  MUX2X1 U481 ( .B(n512), .A(n508), .S(n373), .Y(n499) );
  MUX2X1 U482 ( .B(A[21]), .A(A[22]), .S(SH[0]), .Y(n508) );
  MUX2X1 U483 ( .B(A[19]), .A(A[20]), .S(SH[0]), .Y(n512) );
  MUX2X1 U484 ( .B(n430), .A(n498), .S(n376), .Y(n449) );
  MUX2X1 U485 ( .B(n514), .A(n511), .S(n373), .Y(n498) );
  MUX2X1 U486 ( .B(A[17]), .A(A[18]), .S(SH[0]), .Y(n511) );
  MUX2X1 U487 ( .B(A[15]), .A(A[16]), .S(SH[0]), .Y(n514) );
  MUX2X1 U488 ( .B(n482), .A(n513), .S(n373), .Y(n430) );
  MUX2X1 U489 ( .B(A[13]), .A(A[14]), .S(SH[0]), .Y(n513) );
  MUX2X1 U490 ( .B(A[11]), .A(A[12]), .S(SH[0]), .Y(n482) );
  MUX2X1 U491 ( .B(n524), .A(n466), .S(n383), .Y(B[10]) );
  MUX2X1 U492 ( .B(n489), .A(A[31]), .S(n380), .Y(n466) );
  MUX2X1 U493 ( .B(n409), .A(n501), .S(n376), .Y(n489) );
  MUX2X1 U494 ( .B(n408), .A(A[31]), .S(n373), .Y(n501) );
  MUX2X1 U495 ( .B(n527), .A(n528), .S(n373), .Y(n526) );
  MUX2X1 U496 ( .B(n458), .A(n488), .S(n380), .Y(n524) );
  MUX2X1 U497 ( .B(n413), .A(n411), .S(n376), .Y(n488) );
  MUX2X1 U498 ( .B(n530), .A(n531), .S(n372), .Y(n529) );
  MUX2X1 U499 ( .B(n533), .A(n534), .S(n372), .Y(n532) );
  MUX2X1 U500 ( .B(n416), .A(n415), .S(n376), .Y(n458) );
  MUX2X1 U501 ( .B(n536), .A(n537), .S(n372), .Y(n535) );
  MUX2X1 U502 ( .B(n538), .A(n539), .S(n372), .Y(n436) );
  MUX2X1 U503 ( .B(n541), .A(n494), .S(n383), .Y(n540) );
  MUX2X1 U504 ( .B(n425), .A(n469), .S(n380), .Y(n494) );
  MUX2X1 U505 ( .B(n519), .A(n516), .S(n376), .Y(n469) );
  MUX2X1 U506 ( .B(n528), .A(n525), .S(n372), .Y(n516) );
  MUX2X1 U507 ( .B(A[30]), .A(A[31]), .S(n370), .Y(n525) );
  MUX2X1 U508 ( .B(A[28]), .A(A[29]), .S(n370), .Y(n528) );
  MUX2X1 U509 ( .B(n531), .A(n527), .S(n372), .Y(n519) );
  MUX2X1 U510 ( .B(A[26]), .A(A[27]), .S(n370), .Y(n527) );
  MUX2X1 U511 ( .B(A[24]), .A(A[25]), .S(SH[0]), .Y(n531) );
  MUX2X1 U512 ( .B(n521), .A(n518), .S(n376), .Y(n425) );
  MUX2X1 U513 ( .B(n534), .A(n530), .S(n372), .Y(n518) );
  MUX2X1 U514 ( .B(A[22]), .A(A[23]), .S(n369), .Y(n530) );
  MUX2X1 U515 ( .B(A[20]), .A(A[21]), .S(n369), .Y(n534) );
  MUX2X1 U516 ( .B(n537), .A(n533), .S(n372), .Y(n521) );
  MUX2X1 U517 ( .B(A[18]), .A(A[19]), .S(n369), .Y(n533) );
  MUX2X1 U518 ( .B(A[16]), .A(A[17]), .S(n369), .Y(n537) );
  MUX2X1 U519 ( .B(n542), .A(n424), .S(n380), .Y(n541) );
  MUX2X1 U520 ( .B(n446), .A(n520), .S(n376), .Y(n424) );
  MUX2X1 U521 ( .B(n539), .A(n536), .S(n372), .Y(n520) );
  MUX2X1 U522 ( .B(A[14]), .A(A[15]), .S(n369), .Y(n536) );
  MUX2X1 U523 ( .B(A[12]), .A(A[13]), .S(n369), .Y(n539) );
  MUX2X1 U524 ( .B(n462), .A(n538), .S(n372), .Y(n446) );
  MUX2X1 U525 ( .B(A[10]), .A(A[11]), .S(n369), .Y(n538) );
  MUX2X1 U526 ( .B(A[8]), .A(A[9]), .S(n369), .Y(n462) );
  MUX2X1 U527 ( .B(n543), .A(n445), .S(n376), .Y(n542) );
  MUX2X1 U528 ( .B(n464), .A(n461), .S(n372), .Y(n445) );
  MUX2X1 U529 ( .B(A[6]), .A(A[7]), .S(n369), .Y(n461) );
  MUX2X1 U530 ( .B(A[4]), .A(A[5]), .S(n369), .Y(n464) );
  MUX2X1 U531 ( .B(n544), .A(n463), .S(n372), .Y(n543) );
  MUX2X1 U532 ( .B(A[2]), .A(A[3]), .S(n369), .Y(n463) );
  MUX2X1 U533 ( .B(A[0]), .A(A[1]), .S(n369), .Y(n544) );
endmodule


module alu_DW_rightsh_17 ( A, DATA_TC, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC;
  wire   n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544;

  INVX1 U329 ( .A(n525), .Y(n408) );
  INVX1 U330 ( .A(n422), .Y(n401) );
  INVX1 U331 ( .A(n380), .Y(n379) );
  INVX1 U332 ( .A(n468), .Y(n405) );
  INVX1 U333 ( .A(n470), .Y(n396) );
  INVX1 U334 ( .A(n434), .Y(n417) );
  INVX1 U335 ( .A(n439), .Y(n390) );
  INVX1 U336 ( .A(n485), .Y(n394) );
  INVX1 U337 ( .A(n378), .Y(n376) );
  INVX1 U338 ( .A(n378), .Y(n377) );
  INVX1 U339 ( .A(n515), .Y(n406) );
  INVX1 U340 ( .A(n522), .Y(n393) );
  INVX1 U341 ( .A(n505), .Y(n398) );
  INVX1 U342 ( .A(n475), .Y(n407) );
  INVX1 U343 ( .A(n387), .Y(B[31]) );
  INVX1 U344 ( .A(n387), .Y(n386) );
  INVX1 U345 ( .A(SH[3]), .Y(n380) );
  INVX1 U346 ( .A(n436), .Y(n416) );
  INVX1 U347 ( .A(n493), .Y(B[16]) );
  INVX1 U348 ( .A(n540), .Y(B[0]) );
  INVX1 U349 ( .A(n375), .Y(n374) );
  INVX1 U350 ( .A(n375), .Y(n373) );
  INVX1 U351 ( .A(n384), .Y(n382) );
  INVX1 U352 ( .A(n384), .Y(n381) );
  INVX1 U353 ( .A(A[31]), .Y(n387) );
  INVX1 U354 ( .A(n490), .Y(n399) );
  INVX1 U355 ( .A(n384), .Y(n383) );
  INVX1 U356 ( .A(n529), .Y(n411) );
  INVX1 U357 ( .A(n510), .Y(n402) );
  INVX1 U358 ( .A(SH[2]), .Y(n378) );
  INVX1 U359 ( .A(n479), .Y(n388) );
  INVX1 U360 ( .A(n495), .Y(n395) );
  INVX1 U361 ( .A(n517), .Y(n410) );
  INVX1 U362 ( .A(n523), .Y(n400) );
  INVX1 U363 ( .A(n420), .Y(n389) );
  INVX1 U364 ( .A(n423), .Y(n412) );
  INVX1 U365 ( .A(n426), .Y(n392) );
  INVX1 U366 ( .A(n442), .Y(n414) );
  INVX1 U367 ( .A(n447), .Y(n391) );
  INVX1 U368 ( .A(SH[1]), .Y(n375) );
  INVX1 U369 ( .A(n372), .Y(n370) );
  INVX1 U370 ( .A(n372), .Y(n369) );
  INVX1 U371 ( .A(SH[4]), .Y(n384) );
  INVX1 U372 ( .A(n372), .Y(n371) );
  INVX1 U373 ( .A(n503), .Y(n397) );
  INVX1 U374 ( .A(n526), .Y(n409) );
  INVX1 U375 ( .A(n535), .Y(n415) );
  INVX1 U376 ( .A(n532), .Y(n413) );
  INVX1 U377 ( .A(SH[0]), .Y(n372) );
  INVX1 U378 ( .A(n459), .Y(n418) );
  MUX2X1 U379 ( .B(n389), .A(n419), .S(n383), .Y(B[9]) );
  MUX2X1 U380 ( .B(n421), .A(n422), .S(SH[3]), .Y(n420) );
  MUX2X1 U381 ( .B(n412), .A(n405), .S(n383), .Y(B[8]) );
  MUX2X1 U382 ( .B(n424), .A(n425), .S(SH[3]), .Y(n423) );
  MUX2X1 U383 ( .B(n392), .A(n396), .S(n383), .Y(B[7]) );
  MUX2X1 U384 ( .B(n427), .A(n428), .S(SH[3]), .Y(n426) );
  MUX2X1 U385 ( .B(n429), .A(n430), .S(SH[2]), .Y(n427) );
  MUX2X1 U386 ( .B(n431), .A(n432), .S(n383), .Y(B[6]) );
  MUX2X1 U387 ( .B(n417), .A(n433), .S(SH[3]), .Y(n431) );
  MUX2X1 U388 ( .B(n435), .A(n436), .S(n376), .Y(n434) );
  MUX2X1 U389 ( .B(n437), .A(n438), .S(n383), .Y(B[5]) );
  MUX2X1 U390 ( .B(n390), .A(n402), .S(SH[3]), .Y(n437) );
  MUX2X1 U391 ( .B(n440), .A(n441), .S(n376), .Y(n439) );
  MUX2X1 U392 ( .B(n414), .A(n407), .S(n383), .Y(B[4]) );
  MUX2X1 U393 ( .B(n443), .A(n444), .S(SH[3]), .Y(n442) );
  MUX2X1 U394 ( .B(n445), .A(n446), .S(SH[2]), .Y(n443) );
  MUX2X1 U395 ( .B(n391), .A(n394), .S(n383), .Y(B[3]) );
  MUX2X1 U396 ( .B(n448), .A(n449), .S(SH[3]), .Y(n447) );
  MUX2X1 U397 ( .B(n450), .A(n429), .S(SH[2]), .Y(n448) );
  MUX2X1 U398 ( .B(n451), .A(n452), .S(SH[1]), .Y(n429) );
  MUX2X1 U399 ( .B(n453), .A(n454), .S(SH[1]), .Y(n450) );
  MUX2X1 U400 ( .B(n455), .A(n387), .S(n382), .Y(B[30]) );
  MUX2X1 U401 ( .B(n456), .A(n457), .S(n382), .Y(B[2]) );
  MUX2X1 U402 ( .B(n418), .A(n458), .S(n379), .Y(n456) );
  MUX2X1 U403 ( .B(n460), .A(n435), .S(n376), .Y(n459) );
  MUX2X1 U404 ( .B(n461), .A(n462), .S(SH[1]), .Y(n435) );
  MUX2X1 U405 ( .B(n463), .A(n464), .S(SH[1]), .Y(n460) );
  MUX2X1 U406 ( .B(n465), .A(n387), .S(n382), .Y(B[29]) );
  MUX2X1 U407 ( .B(n406), .A(n387), .S(n382), .Y(B[28]) );
  MUX2X1 U408 ( .B(n393), .A(n387), .S(n382), .Y(B[27]) );
  MUX2X1 U409 ( .B(n466), .A(n387), .S(n382), .Y(B[26]) );
  MUX2X1 U410 ( .B(n419), .A(n387), .S(n382), .Y(B[25]) );
  MUX2X1 U411 ( .B(n467), .A(B[31]), .S(n379), .Y(n419) );
  MUX2X1 U412 ( .B(n405), .A(n387), .S(n382), .Y(B[24]) );
  MUX2X1 U413 ( .B(n469), .A(n387), .S(n379), .Y(n468) );
  MUX2X1 U414 ( .B(n396), .A(n387), .S(n382), .Y(B[23]) );
  MUX2X1 U415 ( .B(n471), .A(n387), .S(n379), .Y(n470) );
  MUX2X1 U416 ( .B(n432), .A(n387), .S(n382), .Y(B[22]) );
  MUX2X1 U417 ( .B(n472), .A(n473), .S(n379), .Y(n432) );
  MUX2X1 U418 ( .B(n438), .A(n387), .S(n382), .Y(B[21]) );
  MUX2X1 U419 ( .B(n398), .A(n474), .S(n379), .Y(n438) );
  MUX2X1 U420 ( .B(n407), .A(n387), .S(n382), .Y(B[20]) );
  MUX2X1 U421 ( .B(n476), .A(n477), .S(n379), .Y(n475) );
  MUX2X1 U422 ( .B(n388), .A(n478), .S(n381), .Y(B[1]) );
  MUX2X1 U423 ( .B(n480), .A(n421), .S(n379), .Y(n479) );
  MUX2X1 U424 ( .B(n441), .A(n481), .S(SH[2]), .Y(n421) );
  MUX2X1 U425 ( .B(n452), .A(n482), .S(SH[1]), .Y(n441) );
  MUX2X1 U426 ( .B(A[9]), .A(A[10]), .S(n371), .Y(n452) );
  MUX2X1 U427 ( .B(n483), .A(n440), .S(n377), .Y(n480) );
  MUX2X1 U428 ( .B(n454), .A(n451), .S(SH[1]), .Y(n440) );
  MUX2X1 U429 ( .B(A[7]), .A(A[8]), .S(n371), .Y(n451) );
  MUX2X1 U430 ( .B(A[5]), .A(A[6]), .S(n371), .Y(n454) );
  MUX2X1 U431 ( .B(n484), .A(n453), .S(SH[1]), .Y(n483) );
  MUX2X1 U432 ( .B(A[3]), .A(A[4]), .S(n371), .Y(n453) );
  MUX2X1 U433 ( .B(A[1]), .A(A[2]), .S(n371), .Y(n484) );
  MUX2X1 U434 ( .B(n394), .A(n387), .S(n381), .Y(B[19]) );
  MUX2X1 U435 ( .B(n486), .A(n487), .S(n379), .Y(n485) );
  MUX2X1 U436 ( .B(n457), .A(n387), .S(n381), .Y(B[18]) );
  MUX2X1 U437 ( .B(n488), .A(n489), .S(n379), .Y(n457) );
  MUX2X1 U438 ( .B(n478), .A(n387), .S(n381), .Y(B[17]) );
  MUX2X1 U439 ( .B(n401), .A(n467), .S(n379), .Y(n478) );
  MUX2X1 U440 ( .B(n399), .A(n397), .S(n377), .Y(n467) );
  MUX2X1 U441 ( .B(n491), .A(n492), .S(n377), .Y(n422) );
  MUX2X1 U442 ( .B(n494), .A(B[31]), .S(n381), .Y(n493) );
  MUX2X1 U443 ( .B(n395), .A(n387), .S(n381), .Y(B[15]) );
  MUX2X1 U444 ( .B(n428), .A(n471), .S(n379), .Y(n495) );
  MUX2X1 U445 ( .B(n496), .A(n497), .S(n377), .Y(n471) );
  MUX2X1 U446 ( .B(n498), .A(n499), .S(n377), .Y(n428) );
  MUX2X1 U447 ( .B(n500), .A(n455), .S(n381), .Y(B[14]) );
  MUX2X1 U448 ( .B(n473), .A(n386), .S(SH[3]), .Y(n455) );
  MUX2X1 U449 ( .B(n501), .A(n387), .S(n377), .Y(n473) );
  MUX2X1 U450 ( .B(n433), .A(n472), .S(SH[3]), .Y(n500) );
  MUX2X1 U451 ( .B(n411), .A(n409), .S(n377), .Y(n472) );
  MUX2X1 U452 ( .B(n415), .A(n413), .S(n377), .Y(n433) );
  MUX2X1 U453 ( .B(n502), .A(n465), .S(n381), .Y(B[13]) );
  MUX2X1 U454 ( .B(n474), .A(n386), .S(SH[3]), .Y(n465) );
  MUX2X1 U455 ( .B(n397), .A(n387), .S(n377), .Y(n474) );
  MUX2X1 U456 ( .B(n504), .A(n387), .S(n374), .Y(n503) );
  MUX2X1 U457 ( .B(n402), .A(n398), .S(SH[3]), .Y(n502) );
  MUX2X1 U458 ( .B(n492), .A(n490), .S(n377), .Y(n505) );
  MUX2X1 U459 ( .B(n506), .A(n507), .S(n374), .Y(n490) );
  MUX2X1 U460 ( .B(n508), .A(n509), .S(n374), .Y(n492) );
  MUX2X1 U461 ( .B(n481), .A(n491), .S(n377), .Y(n510) );
  MUX2X1 U462 ( .B(n511), .A(n512), .S(n374), .Y(n491) );
  MUX2X1 U463 ( .B(n513), .A(n514), .S(n374), .Y(n481) );
  MUX2X1 U464 ( .B(n410), .A(n406), .S(n381), .Y(B[12]) );
  MUX2X1 U465 ( .B(n477), .A(n387), .S(SH[3]), .Y(n515) );
  MUX2X1 U466 ( .B(n516), .A(n386), .S(n377), .Y(n477) );
  MUX2X1 U467 ( .B(n444), .A(n476), .S(SH[3]), .Y(n517) );
  MUX2X1 U468 ( .B(n518), .A(n519), .S(n376), .Y(n476) );
  MUX2X1 U469 ( .B(n520), .A(n521), .S(n376), .Y(n444) );
  MUX2X1 U470 ( .B(n400), .A(n393), .S(n381), .Y(B[11]) );
  MUX2X1 U471 ( .B(n487), .A(n387), .S(SH[3]), .Y(n522) );
  MUX2X1 U472 ( .B(n497), .A(n386), .S(n376), .Y(n487) );
  MUX2X1 U473 ( .B(n507), .A(n504), .S(n374), .Y(n497) );
  MUX2X1 U474 ( .B(A[29]), .A(A[30]), .S(n371), .Y(n504) );
  MUX2X1 U475 ( .B(A[27]), .A(A[28]), .S(n371), .Y(n507) );
  MUX2X1 U476 ( .B(n449), .A(n486), .S(SH[3]), .Y(n523) );
  MUX2X1 U477 ( .B(n499), .A(n496), .S(n376), .Y(n486) );
  MUX2X1 U478 ( .B(n509), .A(n506), .S(n374), .Y(n496) );
  MUX2X1 U479 ( .B(A[25]), .A(A[26]), .S(n370), .Y(n506) );
  MUX2X1 U480 ( .B(A[23]), .A(A[24]), .S(n370), .Y(n509) );
  MUX2X1 U481 ( .B(n512), .A(n508), .S(n374), .Y(n499) );
  MUX2X1 U482 ( .B(A[21]), .A(A[22]), .S(n370), .Y(n508) );
  MUX2X1 U483 ( .B(A[19]), .A(A[20]), .S(n370), .Y(n512) );
  MUX2X1 U484 ( .B(n430), .A(n498), .S(n376), .Y(n449) );
  MUX2X1 U485 ( .B(n514), .A(n511), .S(n374), .Y(n498) );
  MUX2X1 U486 ( .B(A[17]), .A(A[18]), .S(n370), .Y(n511) );
  MUX2X1 U487 ( .B(A[15]), .A(A[16]), .S(n370), .Y(n514) );
  MUX2X1 U488 ( .B(n482), .A(n513), .S(n374), .Y(n430) );
  MUX2X1 U489 ( .B(A[13]), .A(A[14]), .S(n370), .Y(n513) );
  MUX2X1 U490 ( .B(A[11]), .A(A[12]), .S(n370), .Y(n482) );
  MUX2X1 U491 ( .B(n524), .A(n466), .S(n381), .Y(B[10]) );
  MUX2X1 U492 ( .B(n489), .A(n386), .S(SH[3]), .Y(n466) );
  MUX2X1 U493 ( .B(n409), .A(n501), .S(n376), .Y(n489) );
  MUX2X1 U494 ( .B(n408), .A(B[31]), .S(n374), .Y(n501) );
  MUX2X1 U495 ( .B(n527), .A(n528), .S(n374), .Y(n526) );
  MUX2X1 U496 ( .B(n458), .A(n488), .S(SH[3]), .Y(n524) );
  MUX2X1 U497 ( .B(n413), .A(n411), .S(n376), .Y(n488) );
  MUX2X1 U498 ( .B(n530), .A(n531), .S(n373), .Y(n529) );
  MUX2X1 U499 ( .B(n533), .A(n534), .S(n373), .Y(n532) );
  MUX2X1 U500 ( .B(n416), .A(n415), .S(n376), .Y(n458) );
  MUX2X1 U501 ( .B(n536), .A(n537), .S(n373), .Y(n535) );
  MUX2X1 U502 ( .B(n538), .A(n539), .S(n373), .Y(n436) );
  MUX2X1 U503 ( .B(n541), .A(n494), .S(n381), .Y(n540) );
  MUX2X1 U504 ( .B(n425), .A(n469), .S(SH[3]), .Y(n494) );
  MUX2X1 U505 ( .B(n519), .A(n516), .S(n376), .Y(n469) );
  MUX2X1 U506 ( .B(n528), .A(n525), .S(n373), .Y(n516) );
  MUX2X1 U507 ( .B(A[30]), .A(n386), .S(n370), .Y(n525) );
  MUX2X1 U508 ( .B(A[28]), .A(A[29]), .S(n370), .Y(n528) );
  MUX2X1 U509 ( .B(n531), .A(n527), .S(n373), .Y(n519) );
  MUX2X1 U510 ( .B(A[26]), .A(A[27]), .S(n370), .Y(n527) );
  MUX2X1 U511 ( .B(A[24]), .A(A[25]), .S(n370), .Y(n531) );
  MUX2X1 U512 ( .B(n521), .A(n518), .S(n376), .Y(n425) );
  MUX2X1 U513 ( .B(n534), .A(n530), .S(n373), .Y(n518) );
  MUX2X1 U514 ( .B(A[22]), .A(A[23]), .S(n369), .Y(n530) );
  MUX2X1 U515 ( .B(A[20]), .A(A[21]), .S(n369), .Y(n534) );
  MUX2X1 U516 ( .B(n537), .A(n533), .S(n373), .Y(n521) );
  MUX2X1 U517 ( .B(A[18]), .A(A[19]), .S(n369), .Y(n533) );
  MUX2X1 U518 ( .B(A[16]), .A(A[17]), .S(n369), .Y(n537) );
  MUX2X1 U519 ( .B(n542), .A(n424), .S(SH[3]), .Y(n541) );
  MUX2X1 U520 ( .B(n446), .A(n520), .S(n376), .Y(n424) );
  MUX2X1 U521 ( .B(n539), .A(n536), .S(n373), .Y(n520) );
  MUX2X1 U522 ( .B(A[14]), .A(A[15]), .S(n369), .Y(n536) );
  MUX2X1 U523 ( .B(A[12]), .A(A[13]), .S(n369), .Y(n539) );
  MUX2X1 U524 ( .B(n462), .A(n538), .S(n373), .Y(n446) );
  MUX2X1 U525 ( .B(A[10]), .A(A[11]), .S(n369), .Y(n538) );
  MUX2X1 U526 ( .B(A[8]), .A(A[9]), .S(n369), .Y(n462) );
  MUX2X1 U527 ( .B(n543), .A(n445), .S(n376), .Y(n542) );
  MUX2X1 U528 ( .B(n464), .A(n461), .S(n373), .Y(n445) );
  MUX2X1 U529 ( .B(A[6]), .A(A[7]), .S(n369), .Y(n461) );
  MUX2X1 U530 ( .B(A[4]), .A(A[5]), .S(n369), .Y(n464) );
  MUX2X1 U531 ( .B(n544), .A(n463), .S(n373), .Y(n543) );
  MUX2X1 U532 ( .B(A[2]), .A(A[3]), .S(n369), .Y(n463) );
  MUX2X1 U533 ( .B(A[0]), .A(A[1]), .S(n369), .Y(n544) );
endmodule


module alu_DW_rightsh_30 ( A, DATA_TC, SH, B );
  input [63:0] A;
  input [4:0] SH;
  output [63:0] B;
  input DATA_TC;
  wire   n1123, n1122, n1121, n1120, n1119, n1118, n1117, n1116, n1115, n1114,
         n1113, n1112, n1111, n1110, n1109, n1108, n722, n724, n726, n728,
         n729, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n772, n784, n785, n786, n787, n788, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107;

  OR2X1 U638 ( .A(n729), .B(n740), .Y(n899) );
  AND2X1 U639 ( .A(n732), .B(n753), .Y(n874) );
  INVX2 U640 ( .A(SH[0]), .Y(n739) );
  OR2X1 U641 ( .A(n760), .B(n734), .Y(n1108) );
  INVX1 U642 ( .A(n1108), .Y(B[63]) );
  OR2X1 U643 ( .A(n761), .B(n862), .Y(n1119) );
  INVX1 U644 ( .A(n1119), .Y(B[52]) );
  OR2X1 U645 ( .A(n814), .B(n760), .Y(n1121) );
  INVX1 U646 ( .A(n1121), .Y(B[50]) );
  OR2X1 U647 ( .A(n726), .B(n760), .Y(n1110) );
  INVX1 U648 ( .A(n1110), .Y(B[61]) );
  OR2X1 U649 ( .A(n722), .B(n760), .Y(n1113) );
  INVX1 U650 ( .A(n1113), .Y(B[58]) );
  OR2X1 U651 ( .A(n761), .B(n813), .Y(n1122) );
  INVX1 U652 ( .A(n1122), .Y(B[49]) );
  OR2X1 U653 ( .A(n731), .B(n761), .Y(n1109) );
  INVX1 U654 ( .A(n1109), .Y(B[62]) );
  OR2X1 U655 ( .A(n857), .B(n761), .Y(n1114) );
  INVX1 U656 ( .A(n1114), .Y(B[57]) );
  OR2X1 U657 ( .A(n761), .B(n812), .Y(n1123) );
  INVX1 U658 ( .A(n1123), .Y(B[48]) );
  OR2X1 U659 ( .A(n724), .B(n760), .Y(n1111) );
  INVX1 U660 ( .A(n1111), .Y(B[60]) );
  OR2X1 U661 ( .A(n761), .B(n859), .Y(n1116) );
  INVX1 U662 ( .A(n1116), .Y(B[55]) );
  OR2X1 U663 ( .A(n858), .B(n761), .Y(n1115) );
  INVX1 U664 ( .A(n1115), .Y(B[56]) );
  AND2X1 U665 ( .A(n820), .B(n758), .Y(n856) );
  INVX1 U666 ( .A(n856), .Y(n722) );
  OR2X1 U667 ( .A(n815), .B(n761), .Y(n1120) );
  INVX1 U668 ( .A(n1120), .Y(B[51]) );
  AND2X1 U669 ( .A(n880), .B(n758), .Y(n847) );
  INVX1 U670 ( .A(n847), .Y(n724) );
  OR2X1 U671 ( .A(n728), .B(n761), .Y(n1112) );
  INVX1 U672 ( .A(n1112), .Y(B[59]) );
  AND2X1 U673 ( .A(n878), .B(n758), .Y(n846) );
  INVX1 U674 ( .A(n846), .Y(n726) );
  OR2X1 U675 ( .A(n761), .B(n861), .Y(n1118) );
  INVX1 U676 ( .A(n1118), .Y(B[53]) );
  AND2X1 U677 ( .A(n821), .B(n758), .Y(n855) );
  INVX1 U678 ( .A(n855), .Y(n728) );
  AND2X1 U679 ( .A(A[63]), .B(n739), .Y(n911) );
  INVX1 U680 ( .A(n911), .Y(n729) );
  OR2X1 U681 ( .A(n761), .B(n860), .Y(n1117) );
  INVX1 U682 ( .A(n1117), .Y(B[54]) );
  AND2X1 U683 ( .A(n876), .B(n758), .Y(n845) );
  INVX1 U684 ( .A(n845), .Y(n731) );
  AND2X1 U685 ( .A(n733), .B(n753), .Y(n876) );
  INVX1 U686 ( .A(n899), .Y(n732) );
  OR2X1 U687 ( .A(n916), .B(n742), .Y(n901) );
  INVX1 U688 ( .A(n901), .Y(n733) );
  AND2X1 U689 ( .A(n874), .B(n758), .Y(n844) );
  INVX1 U690 ( .A(n844), .Y(n734) );
  INVX1 U691 ( .A(n1018), .Y(B[18]) );
  INVX1 U692 ( .A(n937), .Y(B[2]) );
  INVX1 U693 ( .A(n867), .Y(n784) );
  INVX1 U694 ( .A(n864), .Y(n814) );
  INVX1 U695 ( .A(n906), .Y(n816) );
  INVX1 U696 ( .A(n900), .Y(n819) );
  INVX1 U697 ( .A(n902), .Y(n818) );
  INVX1 U698 ( .A(n904), .Y(n817) );
  INVX1 U699 ( .A(n986), .Y(n802) );
  INVX1 U700 ( .A(n992), .Y(n801) );
  INVX1 U701 ( .A(n973), .Y(n804) );
  INVX1 U702 ( .A(n980), .Y(n803) );
  INVX1 U703 ( .A(n998), .Y(n800) );
  INVX1 U704 ( .A(n977), .Y(n788) );
  INVX1 U705 ( .A(n882), .Y(n821) );
  INVX1 U706 ( .A(n865), .Y(B[4]) );
  INVX1 U707 ( .A(n884), .Y(n820) );
  INVX1 U708 ( .A(n753), .Y(n750) );
  INVX1 U709 ( .A(n753), .Y(n749) );
  INVX1 U710 ( .A(n753), .Y(n752) );
  INVX1 U711 ( .A(n753), .Y(n751) );
  INVX1 U712 ( .A(n741), .Y(n745) );
  INVX1 U713 ( .A(n741), .Y(n746) );
  INVX1 U714 ( .A(n758), .Y(n756) );
  INVX1 U715 ( .A(n758), .Y(n757) );
  INVX1 U716 ( .A(n758), .Y(n755) );
  INVX1 U717 ( .A(n758), .Y(n754) );
  INVX1 U718 ( .A(n881), .Y(n808) );
  INVX1 U719 ( .A(n887), .Y(n805) );
  INVX1 U720 ( .A(n967), .Y(B[25]) );
  INVX1 U721 ( .A(n1076), .Y(B[12]) );
  INVX1 U722 ( .A(n1090), .Y(B[10]) );
  INVX1 U723 ( .A(n922), .Y(B[32]) );
  INVX1 U724 ( .A(n883), .Y(n807) );
  INVX1 U725 ( .A(n875), .Y(n811) );
  INVX1 U726 ( .A(n927), .Y(B[31]) );
  INVX1 U727 ( .A(n1039), .Y(B[15]) );
  INVX1 U728 ( .A(n1049), .Y(B[14]) );
  INVX1 U729 ( .A(n1033), .Y(B[16]) );
  INVX1 U730 ( .A(n889), .Y(B[3]) );
  INVX1 U731 ( .A(n1059), .Y(B[13]) );
  INVX1 U732 ( .A(n822), .Y(B[9]) );
  INVX1 U733 ( .A(n837), .Y(B[6]) );
  INVX1 U734 ( .A(n917), .Y(B[33]) );
  INVX1 U735 ( .A(n872), .Y(n813) );
  INVX1 U736 ( .A(n879), .Y(n809) );
  INVX1 U737 ( .A(n947), .Y(B[29]) );
  INVX1 U738 ( .A(n839), .Y(n786) );
  INVX1 U739 ( .A(n1024), .Y(B[17]) );
  INVX1 U740 ( .A(n877), .Y(n810) );
  INVX1 U741 ( .A(n848), .Y(B[5]) );
  INVX1 U742 ( .A(n850), .Y(n785) );
  INVX1 U743 ( .A(n957), .Y(B[27]) );
  INVX1 U744 ( .A(n1103), .Y(B[0]) );
  INVX1 U745 ( .A(n827), .Y(n772) );
  INVX1 U746 ( .A(n885), .Y(n806) );
  INVX1 U747 ( .A(n830), .Y(B[7]) );
  INVX1 U748 ( .A(n832), .Y(n787) );
  INVX1 U749 ( .A(n1088), .Y(B[11]) );
  INVX1 U750 ( .A(n907), .Y(B[35]) );
  INVX1 U751 ( .A(n932), .Y(B[30]) );
  INVX1 U752 ( .A(n962), .Y(B[26]) );
  INVX1 U753 ( .A(n873), .Y(n812) );
  INVX1 U754 ( .A(n743), .Y(n742) );
  INVX1 U755 ( .A(n743), .Y(n741) );
  INVX1 U756 ( .A(n739), .Y(n735) );
  INVX1 U757 ( .A(n739), .Y(n738) );
  INVX1 U758 ( .A(n739), .Y(n737) );
  INVX1 U759 ( .A(n739), .Y(n736) );
  INVX1 U760 ( .A(n740), .Y(n747) );
  INVX1 U761 ( .A(n740), .Y(n748) );
  INVX1 U762 ( .A(n863), .Y(n815) );
  OR2X1 U763 ( .A(n886), .B(SH[3]), .Y(n857) );
  INVX1 U764 ( .A(SH[2]), .Y(n753) );
  INVX1 U765 ( .A(n1004), .Y(B[1]) );
  INVX1 U766 ( .A(n1012), .Y(B[19]) );
  INVX1 U767 ( .A(n952), .Y(B[28]) );
  INVX1 U768 ( .A(n912), .Y(B[34]) );
  INVX1 U769 ( .A(SH[3]), .Y(n758) );
  INVX1 U770 ( .A(SH[1]), .Y(n743) );
  INVX1 U771 ( .A(n763), .Y(n762) );
  INVX1 U772 ( .A(n763), .Y(n761) );
  INVX1 U773 ( .A(n763), .Y(n760) );
  INVX1 U774 ( .A(n763), .Y(n759) );
  INVX1 U775 ( .A(n744), .Y(n740) );
  INVX1 U776 ( .A(SH[1]), .Y(n744) );
  INVX1 U777 ( .A(SH[4]), .Y(n763) );
  MUX2X1 U778 ( .B(n823), .A(n824), .S(n759), .Y(n822) );
  MUX2X1 U779 ( .B(n825), .A(n826), .S(n754), .Y(n823) );
  MUX2X1 U780 ( .B(n772), .A(n788), .S(n759), .Y(B[8]) );
  MUX2X1 U781 ( .B(n828), .A(n829), .S(n756), .Y(n827) );
  MUX2X1 U782 ( .B(n831), .A(n832), .S(n759), .Y(n830) );
  MUX2X1 U783 ( .B(n833), .A(n834), .S(n755), .Y(n831) );
  MUX2X1 U784 ( .B(n835), .A(n836), .S(n749), .Y(n833) );
  MUX2X1 U785 ( .B(n838), .A(n839), .S(n759), .Y(n837) );
  MUX2X1 U786 ( .B(n840), .A(n841), .S(n756), .Y(n838) );
  MUX2X1 U787 ( .B(n842), .A(n843), .S(n749), .Y(n840) );
  MUX2X1 U788 ( .B(n849), .A(n850), .S(n761), .Y(n848) );
  MUX2X1 U789 ( .B(n851), .A(n852), .S(n755), .Y(n849) );
  MUX2X1 U790 ( .B(n853), .A(n854), .S(n749), .Y(n851) );
  MUX2X1 U791 ( .B(n866), .A(n867), .S(n759), .Y(n865) );
  MUX2X1 U792 ( .B(n868), .A(n869), .S(n756), .Y(n866) );
  MUX2X1 U793 ( .B(n870), .A(n871), .S(n749), .Y(n868) );
  MUX2X1 U794 ( .B(n811), .A(n734), .S(n759), .Y(B[47]) );
  MUX2X1 U795 ( .B(n810), .A(n731), .S(n759), .Y(B[46]) );
  MUX2X1 U796 ( .B(n809), .A(n726), .S(n759), .Y(B[45]) );
  MUX2X1 U797 ( .B(n808), .A(n724), .S(n759), .Y(B[44]) );
  MUX2X1 U798 ( .B(n807), .A(n728), .S(n759), .Y(B[43]) );
  MUX2X1 U799 ( .B(n806), .A(n722), .S(n759), .Y(B[42]) );
  MUX2X1 U800 ( .B(n805), .A(n857), .S(n760), .Y(B[41]) );
  MUX2X1 U801 ( .B(n804), .A(n858), .S(n760), .Y(B[40]) );
  OR2X1 U802 ( .A(n888), .B(n755), .Y(n858) );
  MUX2X1 U803 ( .B(n890), .A(n891), .S(n760), .Y(n889) );
  MUX2X1 U804 ( .B(n892), .A(n893), .S(n755), .Y(n890) );
  MUX2X1 U805 ( .B(n894), .A(n835), .S(n749), .Y(n892) );
  MUX2X1 U806 ( .B(n895), .A(n896), .S(n741), .Y(n835) );
  MUX2X1 U807 ( .B(n897), .A(n898), .S(n741), .Y(n894) );
  MUX2X1 U808 ( .B(n803), .A(n859), .S(n760), .Y(B[39]) );
  MUX2X1 U809 ( .B(n819), .A(n874), .S(n756), .Y(n859) );
  MUX2X1 U810 ( .B(n802), .A(n860), .S(n760), .Y(B[38]) );
  MUX2X1 U811 ( .B(n818), .A(n876), .S(n756), .Y(n860) );
  MUX2X1 U812 ( .B(n801), .A(n861), .S(n760), .Y(B[37]) );
  MUX2X1 U813 ( .B(n817), .A(n878), .S(n757), .Y(n861) );
  AND2X1 U814 ( .A(n903), .B(n753), .Y(n878) );
  MUX2X1 U815 ( .B(n800), .A(n862), .S(n760), .Y(B[36]) );
  MUX2X1 U816 ( .B(n816), .A(n880), .S(n757), .Y(n862) );
  AND2X1 U817 ( .A(n905), .B(n753), .Y(n880) );
  MUX2X1 U818 ( .B(n908), .A(n863), .S(n760), .Y(n907) );
  MUX2X1 U819 ( .B(n909), .A(n882), .S(n757), .Y(n863) );
  MUX2X1 U820 ( .B(n910), .A(n732), .S(n749), .Y(n882) );
  MUX2X1 U821 ( .B(n913), .A(n864), .S(n760), .Y(n912) );
  MUX2X1 U822 ( .B(n914), .A(n884), .S(n757), .Y(n864) );
  MUX2X1 U823 ( .B(n915), .A(n733), .S(n749), .Y(n884) );
  MUX2X1 U824 ( .B(n918), .A(n872), .S(n760), .Y(n917) );
  MUX2X1 U825 ( .B(n919), .A(n886), .S(n757), .Y(n872) );
  MUX2X1 U826 ( .B(n920), .A(n903), .S(n749), .Y(n886) );
  MUX2X1 U827 ( .B(n729), .A(n921), .S(n745), .Y(n903) );
  MUX2X1 U828 ( .B(n923), .A(n873), .S(n760), .Y(n922) );
  MUX2X1 U829 ( .B(n924), .A(n888), .S(n757), .Y(n873) );
  MUX2X1 U830 ( .B(n925), .A(n905), .S(n749), .Y(n888) );
  MUX2X1 U831 ( .B(n916), .A(n926), .S(n745), .Y(n905) );
  MUX2X1 U832 ( .B(A[62]), .A(A[63]), .S(n735), .Y(n916) );
  MUX2X1 U833 ( .B(n928), .A(n875), .S(n760), .Y(n927) );
  MUX2X1 U834 ( .B(n929), .A(n900), .S(n757), .Y(n875) );
  MUX2X1 U835 ( .B(n930), .A(n910), .S(n749), .Y(n900) );
  MUX2X1 U836 ( .B(n921), .A(n931), .S(n745), .Y(n910) );
  MUX2X1 U837 ( .B(A[61]), .A(A[62]), .S(n735), .Y(n921) );
  MUX2X1 U838 ( .B(n933), .A(n877), .S(n761), .Y(n932) );
  MUX2X1 U839 ( .B(n934), .A(n902), .S(n757), .Y(n877) );
  MUX2X1 U840 ( .B(n935), .A(n915), .S(n749), .Y(n902) );
  MUX2X1 U841 ( .B(n926), .A(n936), .S(n745), .Y(n915) );
  MUX2X1 U842 ( .B(A[60]), .A(A[61]), .S(n735), .Y(n926) );
  MUX2X1 U843 ( .B(n938), .A(n939), .S(n761), .Y(n937) );
  MUX2X1 U844 ( .B(n940), .A(n941), .S(n757), .Y(n938) );
  MUX2X1 U845 ( .B(n942), .A(n842), .S(n749), .Y(n940) );
  MUX2X1 U846 ( .B(n943), .A(n944), .S(n742), .Y(n842) );
  MUX2X1 U847 ( .B(n945), .A(n946), .S(n742), .Y(n942) );
  MUX2X1 U848 ( .B(n948), .A(n879), .S(n761), .Y(n947) );
  MUX2X1 U849 ( .B(n949), .A(n904), .S(n757), .Y(n879) );
  MUX2X1 U850 ( .B(n950), .A(n920), .S(n750), .Y(n904) );
  MUX2X1 U851 ( .B(n931), .A(n951), .S(n745), .Y(n920) );
  MUX2X1 U852 ( .B(A[59]), .A(A[60]), .S(n735), .Y(n931) );
  MUX2X1 U853 ( .B(n953), .A(n881), .S(n761), .Y(n952) );
  MUX2X1 U854 ( .B(n954), .A(n906), .S(n757), .Y(n881) );
  MUX2X1 U855 ( .B(n955), .A(n925), .S(n750), .Y(n906) );
  MUX2X1 U856 ( .B(n936), .A(n956), .S(n745), .Y(n925) );
  MUX2X1 U857 ( .B(A[58]), .A(A[59]), .S(n735), .Y(n936) );
  MUX2X1 U858 ( .B(n958), .A(n883), .S(n761), .Y(n957) );
  MUX2X1 U859 ( .B(n959), .A(n909), .S(n757), .Y(n883) );
  MUX2X1 U860 ( .B(n960), .A(n930), .S(n750), .Y(n909) );
  MUX2X1 U861 ( .B(n951), .A(n961), .S(n745), .Y(n930) );
  MUX2X1 U862 ( .B(A[57]), .A(A[58]), .S(n735), .Y(n951) );
  MUX2X1 U863 ( .B(n963), .A(n885), .S(n761), .Y(n962) );
  MUX2X1 U864 ( .B(n964), .A(n914), .S(n756), .Y(n885) );
  MUX2X1 U865 ( .B(n965), .A(n935), .S(n750), .Y(n914) );
  MUX2X1 U866 ( .B(n956), .A(n966), .S(n745), .Y(n935) );
  MUX2X1 U867 ( .B(A[56]), .A(A[57]), .S(n735), .Y(n956) );
  MUX2X1 U868 ( .B(n824), .A(n887), .S(n761), .Y(n967) );
  MUX2X1 U869 ( .B(n968), .A(n919), .S(n756), .Y(n887) );
  MUX2X1 U870 ( .B(n969), .A(n950), .S(n750), .Y(n919) );
  MUX2X1 U871 ( .B(n961), .A(n970), .S(n745), .Y(n950) );
  MUX2X1 U872 ( .B(A[55]), .A(A[56]), .S(n735), .Y(n961) );
  MUX2X1 U873 ( .B(n971), .A(n972), .S(n756), .Y(n824) );
  MUX2X1 U874 ( .B(n788), .A(n804), .S(n761), .Y(B[24]) );
  MUX2X1 U875 ( .B(n974), .A(n924), .S(n756), .Y(n973) );
  MUX2X1 U876 ( .B(n975), .A(n955), .S(n750), .Y(n924) );
  MUX2X1 U877 ( .B(n966), .A(n976), .S(n745), .Y(n955) );
  MUX2X1 U878 ( .B(A[54]), .A(A[55]), .S(n735), .Y(n966) );
  MUX2X1 U879 ( .B(n978), .A(n979), .S(n756), .Y(n977) );
  MUX2X1 U880 ( .B(n787), .A(n803), .S(n761), .Y(B[23]) );
  MUX2X1 U881 ( .B(n981), .A(n929), .S(n756), .Y(n980) );
  MUX2X1 U882 ( .B(n982), .A(n960), .S(n750), .Y(n929) );
  MUX2X1 U883 ( .B(n970), .A(n983), .S(n745), .Y(n960) );
  MUX2X1 U884 ( .B(A[53]), .A(A[54]), .S(n735), .Y(n970) );
  MUX2X1 U885 ( .B(n984), .A(n985), .S(n756), .Y(n832) );
  MUX2X1 U886 ( .B(n786), .A(n802), .S(n761), .Y(B[22]) );
  MUX2X1 U887 ( .B(n987), .A(n934), .S(n756), .Y(n986) );
  MUX2X1 U888 ( .B(n988), .A(n965), .S(n750), .Y(n934) );
  MUX2X1 U889 ( .B(n976), .A(n989), .S(n745), .Y(n965) );
  MUX2X1 U890 ( .B(A[52]), .A(A[53]), .S(n735), .Y(n976) );
  MUX2X1 U891 ( .B(n990), .A(n991), .S(n756), .Y(n839) );
  MUX2X1 U892 ( .B(n785), .A(n801), .S(n761), .Y(B[21]) );
  MUX2X1 U893 ( .B(n993), .A(n949), .S(n756), .Y(n992) );
  MUX2X1 U894 ( .B(n994), .A(n969), .S(n750), .Y(n949) );
  MUX2X1 U895 ( .B(n983), .A(n995), .S(n746), .Y(n969) );
  MUX2X1 U896 ( .B(A[51]), .A(A[52]), .S(n735), .Y(n983) );
  MUX2X1 U897 ( .B(n996), .A(n997), .S(n756), .Y(n850) );
  MUX2X1 U898 ( .B(n784), .A(n800), .S(n762), .Y(B[20]) );
  MUX2X1 U899 ( .B(n999), .A(n954), .S(n755), .Y(n998) );
  MUX2X1 U900 ( .B(n1000), .A(n975), .S(n750), .Y(n954) );
  MUX2X1 U901 ( .B(n989), .A(n1001), .S(n746), .Y(n975) );
  MUX2X1 U902 ( .B(A[50]), .A(A[51]), .S(n736), .Y(n989) );
  MUX2X1 U903 ( .B(n1002), .A(n1003), .S(n755), .Y(n867) );
  MUX2X1 U904 ( .B(n1005), .A(n1006), .S(n762), .Y(n1004) );
  MUX2X1 U905 ( .B(n1007), .A(n825), .S(n755), .Y(n1005) );
  MUX2X1 U906 ( .B(n1008), .A(n854), .S(n753), .Y(n825) );
  MUX2X1 U907 ( .B(n896), .A(n1009), .S(n742), .Y(n854) );
  MUX2X1 U908 ( .B(A[9]), .A(A[10]), .S(n736), .Y(n896) );
  MUX2X1 U909 ( .B(n1010), .A(n853), .S(n750), .Y(n1007) );
  MUX2X1 U910 ( .B(n898), .A(n895), .S(n742), .Y(n853) );
  MUX2X1 U911 ( .B(A[7]), .A(A[8]), .S(n736), .Y(n895) );
  MUX2X1 U912 ( .B(A[5]), .A(A[6]), .S(n736), .Y(n898) );
  MUX2X1 U913 ( .B(n1011), .A(n897), .S(n742), .Y(n1010) );
  MUX2X1 U914 ( .B(A[3]), .A(A[4]), .S(n736), .Y(n897) );
  MUX2X1 U915 ( .B(A[1]), .A(A[2]), .S(n736), .Y(n1011) );
  MUX2X1 U916 ( .B(n891), .A(n908), .S(n762), .Y(n1012) );
  MUX2X1 U917 ( .B(n1013), .A(n959), .S(n755), .Y(n908) );
  MUX2X1 U918 ( .B(n1014), .A(n982), .S(n750), .Y(n959) );
  MUX2X1 U919 ( .B(n995), .A(n1015), .S(n746), .Y(n982) );
  MUX2X1 U920 ( .B(A[49]), .A(A[50]), .S(n736), .Y(n995) );
  MUX2X1 U921 ( .B(n1016), .A(n1017), .S(n755), .Y(n891) );
  MUX2X1 U922 ( .B(n939), .A(n913), .S(n762), .Y(n1018) );
  MUX2X1 U923 ( .B(n1019), .A(n964), .S(n755), .Y(n913) );
  MUX2X1 U924 ( .B(n1020), .A(n988), .S(n751), .Y(n964) );
  MUX2X1 U925 ( .B(n1001), .A(n1021), .S(n746), .Y(n988) );
  MUX2X1 U926 ( .B(A[48]), .A(A[49]), .S(n736), .Y(n1001) );
  MUX2X1 U927 ( .B(n1022), .A(n1023), .S(n755), .Y(n939) );
  MUX2X1 U928 ( .B(n1006), .A(n918), .S(n762), .Y(n1024) );
  MUX2X1 U929 ( .B(n972), .A(n968), .S(n755), .Y(n918) );
  MUX2X1 U930 ( .B(n1025), .A(n994), .S(n751), .Y(n968) );
  MUX2X1 U931 ( .B(n1015), .A(n1026), .S(n746), .Y(n994) );
  MUX2X1 U932 ( .B(A[47]), .A(A[48]), .S(n736), .Y(n1015) );
  MUX2X1 U933 ( .B(n1027), .A(n1028), .S(n751), .Y(n972) );
  MUX2X1 U934 ( .B(n826), .A(n971), .S(n755), .Y(n1006) );
  MUX2X1 U935 ( .B(n1029), .A(n1030), .S(n751), .Y(n971) );
  MUX2X1 U936 ( .B(n1031), .A(n1032), .S(n751), .Y(n826) );
  MUX2X1 U937 ( .B(n1034), .A(n923), .S(n762), .Y(n1033) );
  MUX2X1 U938 ( .B(n979), .A(n974), .S(n755), .Y(n923) );
  MUX2X1 U939 ( .B(n1035), .A(n1000), .S(n751), .Y(n974) );
  MUX2X1 U940 ( .B(n1021), .A(n1036), .S(n746), .Y(n1000) );
  MUX2X1 U941 ( .B(A[46]), .A(A[47]), .S(n736), .Y(n1021) );
  MUX2X1 U942 ( .B(n1037), .A(n1038), .S(n751), .Y(n979) );
  MUX2X1 U943 ( .B(n1040), .A(n928), .S(n762), .Y(n1039) );
  MUX2X1 U944 ( .B(n985), .A(n981), .S(n755), .Y(n928) );
  MUX2X1 U945 ( .B(n1041), .A(n1014), .S(n751), .Y(n981) );
  MUX2X1 U946 ( .B(n1026), .A(n1042), .S(n746), .Y(n1014) );
  MUX2X1 U947 ( .B(A[45]), .A(A[46]), .S(n736), .Y(n1026) );
  MUX2X1 U948 ( .B(n1043), .A(n1044), .S(n751), .Y(n985) );
  MUX2X1 U949 ( .B(n834), .A(n984), .S(n755), .Y(n1040) );
  MUX2X1 U950 ( .B(n1045), .A(n1046), .S(n751), .Y(n984) );
  MUX2X1 U951 ( .B(n1047), .A(n1048), .S(n751), .Y(n834) );
  MUX2X1 U952 ( .B(n1050), .A(n933), .S(n762), .Y(n1049) );
  MUX2X1 U953 ( .B(n991), .A(n987), .S(n754), .Y(n933) );
  MUX2X1 U954 ( .B(n1051), .A(n1020), .S(n751), .Y(n987) );
  MUX2X1 U955 ( .B(n1036), .A(n1052), .S(n746), .Y(n1020) );
  MUX2X1 U956 ( .B(A[44]), .A(A[45]), .S(n736), .Y(n1036) );
  MUX2X1 U957 ( .B(n1053), .A(n1054), .S(n752), .Y(n991) );
  MUX2X1 U958 ( .B(n841), .A(n990), .S(n754), .Y(n1050) );
  MUX2X1 U959 ( .B(n1055), .A(n1056), .S(n752), .Y(n990) );
  MUX2X1 U960 ( .B(n1057), .A(n1058), .S(n752), .Y(n841) );
  MUX2X1 U961 ( .B(n1060), .A(n948), .S(n762), .Y(n1059) );
  MUX2X1 U962 ( .B(n997), .A(n993), .S(n754), .Y(n948) );
  MUX2X1 U963 ( .B(n1028), .A(n1025), .S(n752), .Y(n993) );
  MUX2X1 U964 ( .B(n1042), .A(n1061), .S(n746), .Y(n1025) );
  MUX2X1 U965 ( .B(A[43]), .A(A[44]), .S(n737), .Y(n1042) );
  MUX2X1 U966 ( .B(n1062), .A(n1063), .S(n746), .Y(n1028) );
  MUX2X1 U967 ( .B(n1030), .A(n1027), .S(n752), .Y(n997) );
  MUX2X1 U968 ( .B(n1064), .A(n1065), .S(n746), .Y(n1027) );
  MUX2X1 U969 ( .B(n1066), .A(n1067), .S(n746), .Y(n1030) );
  MUX2X1 U970 ( .B(n852), .A(n996), .S(n754), .Y(n1060) );
  MUX2X1 U971 ( .B(n1032), .A(n1029), .S(n752), .Y(n996) );
  MUX2X1 U972 ( .B(n1068), .A(n1069), .S(n747), .Y(n1029) );
  MUX2X1 U973 ( .B(n1070), .A(n1071), .S(n747), .Y(n1032) );
  MUX2X1 U974 ( .B(n1008), .A(n1031), .S(n752), .Y(n852) );
  MUX2X1 U975 ( .B(n1072), .A(n1073), .S(n747), .Y(n1031) );
  MUX2X1 U976 ( .B(n1074), .A(n1075), .S(n747), .Y(n1008) );
  MUX2X1 U977 ( .B(n1077), .A(n953), .S(n762), .Y(n1076) );
  MUX2X1 U978 ( .B(n1003), .A(n999), .S(n754), .Y(n953) );
  MUX2X1 U979 ( .B(n1038), .A(n1035), .S(n752), .Y(n999) );
  MUX2X1 U980 ( .B(n1052), .A(n1078), .S(n747), .Y(n1035) );
  MUX2X1 U981 ( .B(A[42]), .A(A[43]), .S(n737), .Y(n1052) );
  MUX2X1 U982 ( .B(n1079), .A(n1080), .S(n747), .Y(n1038) );
  MUX2X1 U983 ( .B(n1081), .A(n1037), .S(n752), .Y(n1003) );
  MUX2X1 U984 ( .B(n1082), .A(n1083), .S(n747), .Y(n1037) );
  MUX2X1 U985 ( .B(n869), .A(n1002), .S(n754), .Y(n1077) );
  MUX2X1 U986 ( .B(n1084), .A(n1085), .S(n752), .Y(n1002) );
  MUX2X1 U987 ( .B(n1086), .A(n1087), .S(n752), .Y(n869) );
  MUX2X1 U988 ( .B(n1089), .A(n958), .S(n762), .Y(n1088) );
  MUX2X1 U989 ( .B(n1017), .A(n1013), .S(n754), .Y(n958) );
  MUX2X1 U990 ( .B(n1044), .A(n1041), .S(n752), .Y(n1013) );
  MUX2X1 U991 ( .B(n1061), .A(n1062), .S(n747), .Y(n1041) );
  MUX2X1 U992 ( .B(A[39]), .A(A[40]), .S(n737), .Y(n1062) );
  MUX2X1 U993 ( .B(A[41]), .A(A[42]), .S(n737), .Y(n1061) );
  MUX2X1 U994 ( .B(n1063), .A(n1064), .S(n747), .Y(n1044) );
  MUX2X1 U995 ( .B(A[35]), .A(A[36]), .S(n737), .Y(n1064) );
  MUX2X1 U996 ( .B(A[37]), .A(A[38]), .S(n737), .Y(n1063) );
  MUX2X1 U997 ( .B(n1046), .A(n1043), .S(SH[2]), .Y(n1017) );
  MUX2X1 U998 ( .B(n1065), .A(n1066), .S(n747), .Y(n1043) );
  MUX2X1 U999 ( .B(A[31]), .A(A[32]), .S(n737), .Y(n1066) );
  MUX2X1 U1000 ( .B(A[33]), .A(A[34]), .S(n737), .Y(n1065) );
  MUX2X1 U1001 ( .B(n1067), .A(n1068), .S(n747), .Y(n1046) );
  MUX2X1 U1002 ( .B(A[27]), .A(A[28]), .S(n737), .Y(n1068) );
  MUX2X1 U1003 ( .B(A[29]), .A(A[30]), .S(n737), .Y(n1067) );
  MUX2X1 U1004 ( .B(n893), .A(n1016), .S(n754), .Y(n1089) );
  MUX2X1 U1005 ( .B(n1048), .A(n1045), .S(n751), .Y(n1016) );
  MUX2X1 U1006 ( .B(n1069), .A(n1070), .S(n747), .Y(n1045) );
  MUX2X1 U1007 ( .B(A[23]), .A(A[24]), .S(n737), .Y(n1070) );
  MUX2X1 U1008 ( .B(A[25]), .A(A[26]), .S(n737), .Y(n1069) );
  MUX2X1 U1009 ( .B(n1071), .A(n1072), .S(n748), .Y(n1048) );
  MUX2X1 U1010 ( .B(A[19]), .A(A[20]), .S(n738), .Y(n1072) );
  MUX2X1 U1011 ( .B(A[21]), .A(A[22]), .S(n738), .Y(n1071) );
  MUX2X1 U1012 ( .B(n836), .A(n1047), .S(SH[2]), .Y(n893) );
  MUX2X1 U1013 ( .B(n1073), .A(n1074), .S(n748), .Y(n1047) );
  MUX2X1 U1014 ( .B(A[15]), .A(A[16]), .S(n738), .Y(n1074) );
  MUX2X1 U1015 ( .B(A[17]), .A(A[18]), .S(n738), .Y(n1073) );
  MUX2X1 U1016 ( .B(n1009), .A(n1075), .S(n742), .Y(n836) );
  MUX2X1 U1017 ( .B(A[13]), .A(A[14]), .S(n738), .Y(n1075) );
  MUX2X1 U1018 ( .B(A[11]), .A(A[12]), .S(n738), .Y(n1009) );
  MUX2X1 U1019 ( .B(n1091), .A(n963), .S(n762), .Y(n1090) );
  MUX2X1 U1020 ( .B(n1023), .A(n1019), .S(n754), .Y(n963) );
  MUX2X1 U1021 ( .B(n1054), .A(n1051), .S(SH[2]), .Y(n1019) );
  MUX2X1 U1022 ( .B(n1078), .A(n1079), .S(n748), .Y(n1051) );
  MUX2X1 U1023 ( .B(A[38]), .A(A[39]), .S(n738), .Y(n1079) );
  MUX2X1 U1024 ( .B(A[40]), .A(A[41]), .S(n738), .Y(n1078) );
  MUX2X1 U1025 ( .B(n1080), .A(n1082), .S(n748), .Y(n1054) );
  MUX2X1 U1026 ( .B(A[34]), .A(A[35]), .S(n738), .Y(n1082) );
  MUX2X1 U1027 ( .B(A[36]), .A(A[37]), .S(n738), .Y(n1080) );
  MUX2X1 U1028 ( .B(n1056), .A(n1053), .S(SH[2]), .Y(n1023) );
  MUX2X1 U1029 ( .B(n1083), .A(n1092), .S(n748), .Y(n1053) );
  MUX2X1 U1030 ( .B(A[32]), .A(A[33]), .S(n738), .Y(n1083) );
  MUX2X1 U1031 ( .B(n1093), .A(n1094), .S(n748), .Y(n1056) );
  MUX2X1 U1032 ( .B(n941), .A(n1022), .S(n754), .Y(n1091) );
  MUX2X1 U1033 ( .B(n1058), .A(n1055), .S(SH[2]), .Y(n1022) );
  MUX2X1 U1034 ( .B(n1095), .A(n1096), .S(n748), .Y(n1055) );
  MUX2X1 U1035 ( .B(n1097), .A(n1098), .S(n748), .Y(n1058) );
  MUX2X1 U1036 ( .B(n843), .A(n1057), .S(SH[2]), .Y(n941) );
  MUX2X1 U1037 ( .B(n1099), .A(n1100), .S(n748), .Y(n1057) );
  MUX2X1 U1038 ( .B(n1101), .A(n1102), .S(n742), .Y(n843) );
  MUX2X1 U1039 ( .B(n1104), .A(n1034), .S(n759), .Y(n1103) );
  MUX2X1 U1040 ( .B(n829), .A(n978), .S(n754), .Y(n1034) );
  MUX2X1 U1041 ( .B(n1085), .A(n1081), .S(n752), .Y(n978) );
  MUX2X1 U1042 ( .B(n1092), .A(n1093), .S(n748), .Y(n1081) );
  MUX2X1 U1043 ( .B(A[28]), .A(A[29]), .S(n738), .Y(n1093) );
  MUX2X1 U1044 ( .B(A[30]), .A(A[31]), .S(n737), .Y(n1092) );
  MUX2X1 U1045 ( .B(n1094), .A(n1095), .S(n748), .Y(n1085) );
  MUX2X1 U1046 ( .B(A[24]), .A(A[25]), .S(n737), .Y(n1095) );
  MUX2X1 U1047 ( .B(A[26]), .A(A[27]), .S(n736), .Y(n1094) );
  MUX2X1 U1048 ( .B(n1087), .A(n1084), .S(n749), .Y(n829) );
  MUX2X1 U1049 ( .B(n1096), .A(n1097), .S(n748), .Y(n1084) );
  MUX2X1 U1050 ( .B(A[20]), .A(A[21]), .S(SH[0]), .Y(n1097) );
  MUX2X1 U1051 ( .B(A[22]), .A(A[23]), .S(n738), .Y(n1096) );
  MUX2X1 U1052 ( .B(n1098), .A(n1099), .S(n747), .Y(n1087) );
  MUX2X1 U1053 ( .B(A[16]), .A(A[17]), .S(n738), .Y(n1099) );
  MUX2X1 U1054 ( .B(A[18]), .A(A[19]), .S(n735), .Y(n1098) );
  MUX2X1 U1055 ( .B(n1105), .A(n828), .S(n756), .Y(n1104) );
  MUX2X1 U1056 ( .B(n871), .A(n1086), .S(n751), .Y(n828) );
  MUX2X1 U1057 ( .B(n1100), .A(n1102), .S(n747), .Y(n1086) );
  MUX2X1 U1058 ( .B(A[12]), .A(A[13]), .S(SH[0]), .Y(n1102) );
  MUX2X1 U1059 ( .B(A[14]), .A(A[15]), .S(n738), .Y(n1100) );
  MUX2X1 U1060 ( .B(n944), .A(n1101), .S(n742), .Y(n871) );
  MUX2X1 U1061 ( .B(A[10]), .A(A[11]), .S(SH[0]), .Y(n1101) );
  MUX2X1 U1062 ( .B(A[8]), .A(A[9]), .S(SH[0]), .Y(n944) );
  MUX2X1 U1063 ( .B(n1106), .A(n870), .S(n750), .Y(n1105) );
  MUX2X1 U1064 ( .B(n946), .A(n943), .S(n741), .Y(n870) );
  MUX2X1 U1065 ( .B(A[6]), .A(A[7]), .S(SH[0]), .Y(n943) );
  MUX2X1 U1066 ( .B(A[4]), .A(A[5]), .S(n735), .Y(n946) );
  MUX2X1 U1067 ( .B(n1107), .A(n945), .S(n742), .Y(n1106) );
  MUX2X1 U1068 ( .B(A[2]), .A(A[3]), .S(n736), .Y(n945) );
  MUX2X1 U1069 ( .B(A[0]), .A(A[1]), .S(n737), .Y(n1107) );
endmodule


module alu_DW_rightsh_31 ( A, DATA_TC, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC;
  wire   n544, n543, n542, n541, n540, n539, n538, n537, n536, n535, n534,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n385, n386, n387, n388, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533;

  OR2X1 U308 ( .A(n361), .B(n369), .Y(n487) );
  AND2X1 U309 ( .A(n360), .B(n374), .Y(n464) );
  AND2X2 U310 ( .A(A[31]), .B(n368), .Y(n499) );
  OR2X1 U311 ( .A(n359), .B(n379), .Y(n536) );
  INVX1 U312 ( .A(n536), .Y(B[29]) );
  OR2X1 U313 ( .A(n363), .B(n379), .Y(n537) );
  INVX1 U314 ( .A(n537), .Y(B[28]) );
  OR2X1 U315 ( .A(n458), .B(n379), .Y(n538) );
  INVX1 U316 ( .A(n538), .Y(B[27]) );
  OR2X1 U317 ( .A(n459), .B(n379), .Y(n539) );
  INVX1 U318 ( .A(n539), .Y(B[26]) );
  OR2X1 U319 ( .A(n401), .B(n379), .Y(n540) );
  INVX1 U320 ( .A(n540), .Y(B[25]) );
  OR2X1 U321 ( .A(n379), .B(n410), .Y(n541) );
  INVX1 U322 ( .A(n541), .Y(B[23]) );
  OR2X1 U323 ( .A(n379), .B(n416), .Y(n542) );
  INVX1 U324 ( .A(n542), .Y(B[22]) );
  OR2X1 U325 ( .A(n379), .B(n422), .Y(n543) );
  INVX1 U326 ( .A(n543), .Y(B[21]) );
  OR2X1 U327 ( .A(n379), .B(n428), .Y(n544) );
  INVX1 U328 ( .A(n544), .Y(B[20]) );
  OR2X1 U329 ( .A(n379), .B(n362), .Y(n534) );
  INVX1 U330 ( .A(n534), .Y(B[31]) );
  OR2X1 U331 ( .A(n379), .B(n366), .Y(n535) );
  INVX1 U332 ( .A(n535), .Y(B[30]) );
  AND2X1 U333 ( .A(n364), .B(n380), .Y(B[24]) );
  AND2X1 U334 ( .A(n466), .B(n377), .Y(n456) );
  INVX1 U335 ( .A(n456), .Y(n359) );
  OR2X1 U336 ( .A(n517), .B(n369), .Y(n493) );
  INVX1 U337 ( .A(n493), .Y(n360) );
  INVX1 U338 ( .A(n499), .Y(n361) );
  AND2X1 U339 ( .A(n462), .B(n377), .Y(n444) );
  INVX1 U340 ( .A(n444), .Y(n362) );
  AND2X1 U341 ( .A(n365), .B(n374), .Y(n462) );
  AND2X1 U342 ( .A(n468), .B(n377), .Y(n457) );
  INVX1 U343 ( .A(n457), .Y(n363) );
  OR2X1 U344 ( .A(n461), .B(n375), .Y(n407) );
  INVX1 U345 ( .A(n407), .Y(n364) );
  INVX1 U346 ( .A(n487), .Y(n365) );
  AND2X1 U347 ( .A(n464), .B(n377), .Y(n445) );
  INVX1 U348 ( .A(n445), .Y(n366) );
  INVX1 U349 ( .A(n463), .Y(n400) );
  INVX1 U350 ( .A(n465), .Y(n399) );
  INVX1 U351 ( .A(n467), .Y(n398) );
  INVX1 U352 ( .A(n469), .Y(n397) );
  INVX1 U353 ( .A(n374), .Y(n373) );
  INVX1 U354 ( .A(SH[1]), .Y(n371) );
  INVX1 U355 ( .A(n470), .Y(B[1]) );
  INVX1 U356 ( .A(SH[1]), .Y(n372) );
  INVX1 U357 ( .A(n368), .Y(n367) );
  INVX1 U358 ( .A(n434), .Y(B[3]) );
  INVX1 U359 ( .A(n446), .Y(B[2]) );
  INVX1 U360 ( .A(n423), .Y(n386) );
  INVX1 U361 ( .A(n488), .Y(n396) );
  INVX1 U362 ( .A(n494), .Y(n395) );
  INVX1 U363 ( .A(n501), .Y(n394) );
  INVX1 U364 ( .A(n511), .Y(n393) );
  INVX1 U365 ( .A(n516), .Y(n392) );
  INVX1 U366 ( .A(n520), .Y(n391) );
  INVX1 U367 ( .A(n405), .Y(B[8]) );
  INVX1 U368 ( .A(n411), .Y(n388) );
  INVX1 U369 ( .A(n429), .Y(n385) );
  INVX1 U370 ( .A(n377), .Y(n376) );
  INVX1 U371 ( .A(n377), .Y(n375) );
  INVX1 U372 ( .A(n370), .Y(n369) );
  INVX1 U373 ( .A(SH[0]), .Y(n368) );
  INVX1 U374 ( .A(n402), .Y(n390) );
  INVX1 U375 ( .A(n529), .Y(B[0]) );
  INVX1 U376 ( .A(SH[2]), .Y(n374) );
  INVX1 U377 ( .A(n417), .Y(n387) );
  INVX1 U378 ( .A(SH[1]), .Y(n370) );
  INVX1 U379 ( .A(SH[3]), .Y(n377) );
  INVX1 U380 ( .A(n380), .Y(n378) );
  INVX1 U381 ( .A(n380), .Y(n379) );
  INVX1 U382 ( .A(SH[4]), .Y(n380) );
  MUX2X1 U383 ( .B(n390), .A(n401), .S(n378), .Y(B[9]) );
  MUX2X1 U384 ( .B(n403), .A(n404), .S(n375), .Y(n402) );
  MUX2X1 U385 ( .B(n406), .A(n364), .S(n378), .Y(n405) );
  MUX2X1 U386 ( .B(n408), .A(n409), .S(n376), .Y(n406) );
  MUX2X1 U387 ( .B(n388), .A(n410), .S(n379), .Y(B[7]) );
  MUX2X1 U388 ( .B(n412), .A(n413), .S(n376), .Y(n411) );
  MUX2X1 U389 ( .B(n414), .A(n415), .S(SH[2]), .Y(n412) );
  MUX2X1 U390 ( .B(n387), .A(n416), .S(n379), .Y(B[6]) );
  MUX2X1 U391 ( .B(n418), .A(n419), .S(n376), .Y(n417) );
  MUX2X1 U392 ( .B(n420), .A(n421), .S(SH[2]), .Y(n418) );
  MUX2X1 U393 ( .B(n386), .A(n422), .S(n378), .Y(B[5]) );
  MUX2X1 U394 ( .B(n424), .A(n425), .S(n376), .Y(n423) );
  MUX2X1 U395 ( .B(n426), .A(n427), .S(SH[2]), .Y(n424) );
  MUX2X1 U396 ( .B(n385), .A(n428), .S(n379), .Y(B[4]) );
  MUX2X1 U397 ( .B(n430), .A(n431), .S(n376), .Y(n429) );
  MUX2X1 U398 ( .B(n432), .A(n433), .S(SH[2]), .Y(n430) );
  MUX2X1 U399 ( .B(n435), .A(n436), .S(n379), .Y(n434) );
  MUX2X1 U400 ( .B(n437), .A(n438), .S(n376), .Y(n435) );
  MUX2X1 U401 ( .B(n439), .A(n414), .S(SH[2]), .Y(n437) );
  MUX2X1 U402 ( .B(n440), .A(n441), .S(SH[1]), .Y(n414) );
  MUX2X1 U403 ( .B(n442), .A(n443), .S(SH[1]), .Y(n439) );
  MUX2X1 U404 ( .B(n447), .A(n448), .S(n378), .Y(n446) );
  MUX2X1 U405 ( .B(n449), .A(n450), .S(n376), .Y(n447) );
  MUX2X1 U406 ( .B(n451), .A(n420), .S(SH[2]), .Y(n449) );
  MUX2X1 U407 ( .B(n452), .A(n453), .S(n369), .Y(n420) );
  MUX2X1 U408 ( .B(n454), .A(n455), .S(n369), .Y(n451) );
  OR2X1 U409 ( .A(n460), .B(n376), .Y(n401) );
  MUX2X1 U410 ( .B(n400), .A(n462), .S(n376), .Y(n410) );
  MUX2X1 U411 ( .B(n399), .A(n464), .S(n376), .Y(n416) );
  MUX2X1 U412 ( .B(n398), .A(n466), .S(n376), .Y(n422) );
  MUX2X1 U413 ( .B(n397), .A(n468), .S(n375), .Y(n428) );
  MUX2X1 U414 ( .B(n471), .A(n472), .S(n378), .Y(n470) );
  MUX2X1 U415 ( .B(n473), .A(n403), .S(n375), .Y(n471) );
  MUX2X1 U416 ( .B(n474), .A(n427), .S(n374), .Y(n403) );
  MUX2X1 U417 ( .B(n441), .A(n475), .S(n369), .Y(n427) );
  MUX2X1 U418 ( .B(A[9]), .A(A[10]), .S(n367), .Y(n441) );
  MUX2X1 U419 ( .B(n476), .A(n426), .S(SH[2]), .Y(n473) );
  MUX2X1 U420 ( .B(n443), .A(n440), .S(n369), .Y(n426) );
  MUX2X1 U421 ( .B(A[7]), .A(A[8]), .S(n367), .Y(n440) );
  MUX2X1 U422 ( .B(A[5]), .A(A[6]), .S(n367), .Y(n443) );
  MUX2X1 U423 ( .B(n477), .A(n442), .S(n369), .Y(n476) );
  MUX2X1 U424 ( .B(A[3]), .A(A[4]), .S(n367), .Y(n442) );
  MUX2X1 U425 ( .B(A[1]), .A(A[2]), .S(SH[0]), .Y(n477) );
  AND2X1 U426 ( .A(n436), .B(n380), .Y(B[19]) );
  MUX2X1 U427 ( .B(n478), .A(n479), .S(n375), .Y(n436) );
  AND2X1 U428 ( .A(n448), .B(n380), .Y(B[18]) );
  MUX2X1 U429 ( .B(n480), .A(n481), .S(n375), .Y(n448) );
  AND2X1 U430 ( .A(n380), .B(n472), .Y(B[17]) );
  MUX2X1 U431 ( .B(n404), .A(n460), .S(n375), .Y(n472) );
  MUX2X1 U432 ( .B(n482), .A(n483), .S(SH[2]), .Y(n460) );
  MUX2X1 U433 ( .B(n484), .A(n485), .S(SH[2]), .Y(n404) );
  AND2X1 U434 ( .A(n486), .B(n380), .Y(B[16]) );
  MUX2X1 U435 ( .B(n396), .A(n362), .S(n378), .Y(B[15]) );
  MUX2X1 U436 ( .B(n413), .A(n463), .S(n375), .Y(n488) );
  MUX2X1 U437 ( .B(n489), .A(n490), .S(SH[2]), .Y(n463) );
  MUX2X1 U438 ( .B(n491), .A(n492), .S(SH[2]), .Y(n413) );
  MUX2X1 U439 ( .B(n395), .A(n366), .S(n378), .Y(B[14]) );
  MUX2X1 U440 ( .B(n419), .A(n465), .S(n375), .Y(n494) );
  MUX2X1 U441 ( .B(n495), .A(n496), .S(SH[2]), .Y(n465) );
  MUX2X1 U442 ( .B(n497), .A(n498), .S(n373), .Y(n419) );
  MUX2X1 U443 ( .B(n394), .A(n359), .S(n378), .Y(B[13]) );
  AND2X1 U444 ( .A(n483), .B(n374), .Y(n466) );
  MUX2X1 U445 ( .B(n361), .A(n500), .S(n371), .Y(n483) );
  MUX2X1 U446 ( .B(n425), .A(n467), .S(n375), .Y(n501) );
  MUX2X1 U447 ( .B(n485), .A(n482), .S(n373), .Y(n467) );
  MUX2X1 U448 ( .B(n502), .A(n503), .S(n371), .Y(n482) );
  MUX2X1 U449 ( .B(n504), .A(n505), .S(n371), .Y(n485) );
  MUX2X1 U450 ( .B(n474), .A(n484), .S(n373), .Y(n425) );
  MUX2X1 U451 ( .B(n506), .A(n507), .S(n371), .Y(n484) );
  MUX2X1 U452 ( .B(n508), .A(n509), .S(n371), .Y(n474) );
  MUX2X1 U453 ( .B(n393), .A(n363), .S(n378), .Y(B[12]) );
  AND2X1 U454 ( .A(n510), .B(n374), .Y(n468) );
  MUX2X1 U455 ( .B(n431), .A(n469), .S(n375), .Y(n511) );
  MUX2X1 U456 ( .B(n512), .A(n513), .S(n373), .Y(n469) );
  MUX2X1 U457 ( .B(n514), .A(n515), .S(n373), .Y(n431) );
  MUX2X1 U458 ( .B(n392), .A(n458), .S(n378), .Y(B[11]) );
  OR2X1 U459 ( .A(n479), .B(n376), .Y(n458) );
  MUX2X1 U460 ( .B(n490), .A(n365), .S(n373), .Y(n479) );
  MUX2X1 U461 ( .B(n500), .A(n502), .S(n371), .Y(n490) );
  MUX2X1 U462 ( .B(A[27]), .A(A[28]), .S(n367), .Y(n502) );
  MUX2X1 U463 ( .B(A[29]), .A(A[30]), .S(n367), .Y(n500) );
  MUX2X1 U464 ( .B(n438), .A(n478), .S(n375), .Y(n516) );
  MUX2X1 U465 ( .B(n492), .A(n489), .S(n373), .Y(n478) );
  MUX2X1 U466 ( .B(n503), .A(n504), .S(n371), .Y(n489) );
  MUX2X1 U467 ( .B(A[23]), .A(A[24]), .S(n367), .Y(n504) );
  MUX2X1 U468 ( .B(A[25]), .A(A[26]), .S(n367), .Y(n503) );
  MUX2X1 U469 ( .B(n505), .A(n506), .S(n371), .Y(n492) );
  MUX2X1 U470 ( .B(A[19]), .A(A[20]), .S(n367), .Y(n506) );
  MUX2X1 U471 ( .B(A[21]), .A(A[22]), .S(n367), .Y(n505) );
  MUX2X1 U472 ( .B(n415), .A(n491), .S(n373), .Y(n438) );
  MUX2X1 U473 ( .B(n507), .A(n508), .S(n371), .Y(n491) );
  MUX2X1 U474 ( .B(A[15]), .A(A[16]), .S(n367), .Y(n508) );
  MUX2X1 U475 ( .B(A[17]), .A(A[18]), .S(SH[0]), .Y(n507) );
  MUX2X1 U476 ( .B(n475), .A(n509), .S(n369), .Y(n415) );
  MUX2X1 U477 ( .B(A[13]), .A(A[14]), .S(SH[0]), .Y(n509) );
  MUX2X1 U478 ( .B(A[11]), .A(A[12]), .S(SH[0]), .Y(n475) );
  MUX2X1 U479 ( .B(n391), .A(n459), .S(n378), .Y(B[10]) );
  OR2X1 U480 ( .A(n481), .B(n375), .Y(n459) );
  MUX2X1 U481 ( .B(n496), .A(n360), .S(n373), .Y(n481) );
  MUX2X1 U482 ( .B(n518), .A(n519), .S(n371), .Y(n496) );
  MUX2X1 U483 ( .B(n450), .A(n480), .S(n375), .Y(n520) );
  MUX2X1 U484 ( .B(n498), .A(n495), .S(n373), .Y(n480) );
  MUX2X1 U485 ( .B(n521), .A(n522), .S(n371), .Y(n495) );
  MUX2X1 U486 ( .B(n523), .A(n524), .S(n371), .Y(n498) );
  MUX2X1 U487 ( .B(n421), .A(n497), .S(n373), .Y(n450) );
  MUX2X1 U488 ( .B(n525), .A(n526), .S(n372), .Y(n497) );
  MUX2X1 U489 ( .B(n527), .A(n528), .S(n369), .Y(n421) );
  MUX2X1 U490 ( .B(n530), .A(n486), .S(n378), .Y(n529) );
  MUX2X1 U491 ( .B(n461), .A(n409), .S(n377), .Y(n486) );
  MUX2X1 U492 ( .B(n515), .A(n512), .S(n373), .Y(n409) );
  MUX2X1 U493 ( .B(n522), .A(n523), .S(n372), .Y(n512) );
  MUX2X1 U494 ( .B(A[20]), .A(A[21]), .S(SH[0]), .Y(n523) );
  MUX2X1 U495 ( .B(A[22]), .A(A[23]), .S(SH[0]), .Y(n522) );
  MUX2X1 U496 ( .B(n524), .A(n525), .S(n372), .Y(n515) );
  MUX2X1 U497 ( .B(A[16]), .A(A[17]), .S(SH[0]), .Y(n525) );
  MUX2X1 U498 ( .B(A[18]), .A(A[19]), .S(SH[0]), .Y(n524) );
  MUX2X1 U499 ( .B(n513), .A(n510), .S(n373), .Y(n461) );
  MUX2X1 U500 ( .B(n517), .A(n518), .S(n372), .Y(n510) );
  MUX2X1 U501 ( .B(A[28]), .A(A[29]), .S(SH[0]), .Y(n518) );
  MUX2X1 U502 ( .B(A[30]), .A(A[31]), .S(SH[0]), .Y(n517) );
  MUX2X1 U503 ( .B(n519), .A(n521), .S(n372), .Y(n513) );
  MUX2X1 U504 ( .B(A[24]), .A(A[25]), .S(SH[0]), .Y(n521) );
  MUX2X1 U505 ( .B(A[26]), .A(A[27]), .S(SH[0]), .Y(n519) );
  MUX2X1 U506 ( .B(n531), .A(n408), .S(n376), .Y(n530) );
  MUX2X1 U507 ( .B(n433), .A(n514), .S(n373), .Y(n408) );
  MUX2X1 U508 ( .B(n526), .A(n528), .S(n372), .Y(n514) );
  MUX2X1 U509 ( .B(A[12]), .A(A[13]), .S(SH[0]), .Y(n528) );
  MUX2X1 U510 ( .B(A[14]), .A(A[15]), .S(n367), .Y(n526) );
  MUX2X1 U511 ( .B(n453), .A(n527), .S(n369), .Y(n433) );
  MUX2X1 U512 ( .B(A[10]), .A(A[11]), .S(n367), .Y(n527) );
  MUX2X1 U513 ( .B(A[8]), .A(A[9]), .S(n367), .Y(n453) );
  MUX2X1 U514 ( .B(n532), .A(n432), .S(n373), .Y(n531) );
  MUX2X1 U515 ( .B(n455), .A(n452), .S(n369), .Y(n432) );
  MUX2X1 U516 ( .B(A[6]), .A(A[7]), .S(n367), .Y(n452) );
  MUX2X1 U517 ( .B(A[4]), .A(A[5]), .S(n367), .Y(n455) );
  MUX2X1 U518 ( .B(n533), .A(n454), .S(SH[1]), .Y(n532) );
  MUX2X1 U519 ( .B(A[2]), .A(A[3]), .S(n367), .Y(n454) );
  MUX2X1 U520 ( .B(A[0]), .A(A[1]), .S(n367), .Y(n533) );
endmodule


module alu_DW_rightsh_32 ( A, DATA_TC, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC;
  wire   n543, n542, n541, n540, n539, n538, n537, n536, n535, n534, n533,
         n358, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n384,
         n385, n386, n387, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532;

  AND2X1 U308 ( .A(n365), .B(n374), .Y(n463) );
  AND2X1 U309 ( .A(n360), .B(n374), .Y(n461) );
  AND2X1 U310 ( .A(n364), .B(n379), .Y(B[24]) );
  OR2X1 U311 ( .A(n358), .B(SH[4]), .Y(n535) );
  INVX1 U312 ( .A(n535), .Y(B[29]) );
  OR2X1 U313 ( .A(n363), .B(SH[4]), .Y(n536) );
  INVX1 U314 ( .A(n536), .Y(B[28]) );
  OR2X1 U315 ( .A(n457), .B(SH[4]), .Y(n537) );
  INVX1 U316 ( .A(n537), .Y(B[27]) );
  OR2X1 U317 ( .A(n458), .B(SH[4]), .Y(n538) );
  INVX1 U318 ( .A(n538), .Y(B[26]) );
  OR2X1 U319 ( .A(n400), .B(SH[4]), .Y(n539) );
  INVX1 U320 ( .A(n539), .Y(B[25]) );
  OR2X1 U321 ( .A(SH[4]), .B(n409), .Y(n540) );
  INVX1 U322 ( .A(n540), .Y(B[23]) );
  OR2X1 U323 ( .A(SH[4]), .B(n415), .Y(n541) );
  INVX1 U324 ( .A(n541), .Y(B[22]) );
  OR2X1 U325 ( .A(SH[4]), .B(n421), .Y(n542) );
  INVX1 U326 ( .A(n542), .Y(B[21]) );
  OR2X1 U327 ( .A(SH[4]), .B(n427), .Y(n543) );
  INVX1 U328 ( .A(n543), .Y(B[20]) );
  OR2X1 U329 ( .A(SH[4]), .B(n361), .Y(n533) );
  INVX1 U330 ( .A(n533), .Y(B[31]) );
  AND2X1 U331 ( .A(n465), .B(n377), .Y(n455) );
  INVX1 U332 ( .A(n455), .Y(n358) );
  OR2X1 U333 ( .A(SH[4]), .B(n366), .Y(n534) );
  INVX1 U334 ( .A(n534), .Y(B[30]) );
  OR2X1 U335 ( .A(n362), .B(SH[1]), .Y(n486) );
  INVX1 U336 ( .A(n486), .Y(n360) );
  AND2X1 U337 ( .A(n461), .B(n377), .Y(n443) );
  INVX1 U338 ( .A(n443), .Y(n361) );
  AND2X1 U339 ( .A(A[31]), .B(n368), .Y(n498) );
  INVX1 U340 ( .A(n498), .Y(n362) );
  AND2X1 U341 ( .A(n467), .B(n377), .Y(n456) );
  INVX1 U342 ( .A(n456), .Y(n363) );
  OR2X1 U343 ( .A(n460), .B(n375), .Y(n406) );
  INVX1 U344 ( .A(n406), .Y(n364) );
  OR2X1 U345 ( .A(n516), .B(n369), .Y(n492) );
  INVX1 U346 ( .A(n492), .Y(n365) );
  AND2X1 U347 ( .A(n463), .B(n377), .Y(n444) );
  INVX1 U348 ( .A(n444), .Y(n366) );
  INVX1 U349 ( .A(n445), .Y(B[2]) );
  INVX1 U350 ( .A(n462), .Y(n399) );
  INVX1 U351 ( .A(n464), .Y(n398) );
  INVX1 U352 ( .A(n466), .Y(n397) );
  INVX1 U353 ( .A(n468), .Y(n396) );
  INVX1 U354 ( .A(n374), .Y(n373) );
  INVX1 U355 ( .A(SH[1]), .Y(n371) );
  INVX1 U356 ( .A(n469), .Y(B[1]) );
  INVX1 U357 ( .A(n416), .Y(n386) );
  INVX1 U358 ( .A(SH[1]), .Y(n372) );
  INVX1 U359 ( .A(n433), .Y(B[3]) );
  INVX1 U360 ( .A(n493), .Y(n394) );
  INVX1 U361 ( .A(n487), .Y(n395) );
  INVX1 U362 ( .A(n500), .Y(n393) );
  INVX1 U363 ( .A(n510), .Y(n392) );
  INVX1 U364 ( .A(n515), .Y(n391) );
  INVX1 U365 ( .A(n519), .Y(n390) );
  INVX1 U366 ( .A(n401), .Y(n389) );
  INVX1 U367 ( .A(n422), .Y(n385) );
  INVX1 U368 ( .A(n404), .Y(B[8]) );
  INVX1 U369 ( .A(n410), .Y(n387) );
  INVX1 U370 ( .A(n428), .Y(n384) );
  INVX1 U371 ( .A(n377), .Y(n376) );
  INVX1 U372 ( .A(n377), .Y(n375) );
  INVX1 U373 ( .A(n370), .Y(n369) );
  INVX1 U374 ( .A(SH[0]), .Y(n368) );
  INVX1 U375 ( .A(n368), .Y(n367) );
  INVX1 U376 ( .A(n528), .Y(B[0]) );
  INVX1 U377 ( .A(SH[2]), .Y(n374) );
  INVX1 U378 ( .A(SH[1]), .Y(n370) );
  INVX1 U379 ( .A(SH[3]), .Y(n377) );
  INVX1 U380 ( .A(n379), .Y(n378) );
  INVX1 U381 ( .A(SH[4]), .Y(n379) );
  MUX2X1 U382 ( .B(n389), .A(n400), .S(n378), .Y(B[9]) );
  MUX2X1 U383 ( .B(n402), .A(n403), .S(n375), .Y(n401) );
  MUX2X1 U384 ( .B(n405), .A(n364), .S(n378), .Y(n404) );
  MUX2X1 U385 ( .B(n407), .A(n408), .S(n376), .Y(n405) );
  MUX2X1 U386 ( .B(n387), .A(n409), .S(SH[4]), .Y(B[7]) );
  MUX2X1 U387 ( .B(n411), .A(n412), .S(n376), .Y(n410) );
  MUX2X1 U388 ( .B(n413), .A(n414), .S(SH[2]), .Y(n411) );
  MUX2X1 U389 ( .B(n386), .A(n415), .S(SH[4]), .Y(B[6]) );
  MUX2X1 U390 ( .B(n417), .A(n418), .S(n376), .Y(n416) );
  MUX2X1 U391 ( .B(n419), .A(n420), .S(SH[2]), .Y(n417) );
  MUX2X1 U392 ( .B(n385), .A(n421), .S(n378), .Y(B[5]) );
  MUX2X1 U393 ( .B(n423), .A(n424), .S(n376), .Y(n422) );
  MUX2X1 U394 ( .B(n425), .A(n426), .S(SH[2]), .Y(n423) );
  MUX2X1 U395 ( .B(n384), .A(n427), .S(SH[4]), .Y(B[4]) );
  MUX2X1 U396 ( .B(n429), .A(n430), .S(n376), .Y(n428) );
  MUX2X1 U397 ( .B(n431), .A(n432), .S(SH[2]), .Y(n429) );
  MUX2X1 U398 ( .B(n434), .A(n435), .S(SH[4]), .Y(n433) );
  MUX2X1 U399 ( .B(n436), .A(n437), .S(n376), .Y(n434) );
  MUX2X1 U400 ( .B(n438), .A(n413), .S(SH[2]), .Y(n436) );
  MUX2X1 U401 ( .B(n439), .A(n440), .S(SH[1]), .Y(n413) );
  MUX2X1 U402 ( .B(n441), .A(n442), .S(n369), .Y(n438) );
  MUX2X1 U403 ( .B(n446), .A(n447), .S(n378), .Y(n445) );
  MUX2X1 U404 ( .B(n448), .A(n449), .S(n376), .Y(n446) );
  MUX2X1 U405 ( .B(n450), .A(n419), .S(SH[2]), .Y(n448) );
  MUX2X1 U406 ( .B(n451), .A(n452), .S(n369), .Y(n419) );
  MUX2X1 U407 ( .B(n453), .A(n454), .S(n369), .Y(n450) );
  OR2X1 U408 ( .A(n459), .B(n376), .Y(n400) );
  MUX2X1 U409 ( .B(n399), .A(n461), .S(n376), .Y(n409) );
  MUX2X1 U410 ( .B(n398), .A(n463), .S(n376), .Y(n415) );
  MUX2X1 U411 ( .B(n397), .A(n465), .S(n376), .Y(n421) );
  MUX2X1 U412 ( .B(n396), .A(n467), .S(n375), .Y(n427) );
  MUX2X1 U413 ( .B(n470), .A(n471), .S(n378), .Y(n469) );
  MUX2X1 U414 ( .B(n472), .A(n402), .S(n375), .Y(n470) );
  MUX2X1 U415 ( .B(n473), .A(n426), .S(n374), .Y(n402) );
  MUX2X1 U416 ( .B(n440), .A(n474), .S(n369), .Y(n426) );
  MUX2X1 U417 ( .B(A[9]), .A(A[10]), .S(n367), .Y(n440) );
  MUX2X1 U418 ( .B(n475), .A(n425), .S(SH[2]), .Y(n472) );
  MUX2X1 U419 ( .B(n442), .A(n439), .S(n369), .Y(n425) );
  MUX2X1 U420 ( .B(A[7]), .A(A[8]), .S(n367), .Y(n439) );
  MUX2X1 U421 ( .B(A[5]), .A(A[6]), .S(n367), .Y(n442) );
  MUX2X1 U422 ( .B(n476), .A(n441), .S(n369), .Y(n475) );
  MUX2X1 U423 ( .B(A[3]), .A(A[4]), .S(n367), .Y(n441) );
  MUX2X1 U424 ( .B(A[1]), .A(A[2]), .S(n367), .Y(n476) );
  AND2X1 U425 ( .A(n435), .B(n379), .Y(B[19]) );
  MUX2X1 U426 ( .B(n477), .A(n478), .S(n375), .Y(n435) );
  AND2X1 U427 ( .A(n447), .B(n379), .Y(B[18]) );
  MUX2X1 U428 ( .B(n479), .A(n480), .S(n375), .Y(n447) );
  AND2X1 U429 ( .A(n379), .B(n471), .Y(B[17]) );
  MUX2X1 U430 ( .B(n403), .A(n459), .S(n375), .Y(n471) );
  MUX2X1 U431 ( .B(n481), .A(n482), .S(SH[2]), .Y(n459) );
  MUX2X1 U432 ( .B(n483), .A(n484), .S(SH[2]), .Y(n403) );
  AND2X1 U433 ( .A(n485), .B(n379), .Y(B[16]) );
  MUX2X1 U434 ( .B(n395), .A(n361), .S(n378), .Y(B[15]) );
  MUX2X1 U435 ( .B(n412), .A(n462), .S(n375), .Y(n487) );
  MUX2X1 U436 ( .B(n488), .A(n489), .S(SH[2]), .Y(n462) );
  MUX2X1 U437 ( .B(n490), .A(n491), .S(SH[2]), .Y(n412) );
  MUX2X1 U438 ( .B(n394), .A(n366), .S(n378), .Y(B[14]) );
  MUX2X1 U439 ( .B(n418), .A(n464), .S(n375), .Y(n493) );
  MUX2X1 U440 ( .B(n494), .A(n495), .S(SH[2]), .Y(n464) );
  MUX2X1 U441 ( .B(n496), .A(n497), .S(n373), .Y(n418) );
  MUX2X1 U442 ( .B(n393), .A(n358), .S(n378), .Y(B[13]) );
  AND2X1 U443 ( .A(n482), .B(n374), .Y(n465) );
  MUX2X1 U444 ( .B(n362), .A(n499), .S(n371), .Y(n482) );
  MUX2X1 U445 ( .B(n424), .A(n466), .S(n375), .Y(n500) );
  MUX2X1 U446 ( .B(n484), .A(n481), .S(n373), .Y(n466) );
  MUX2X1 U447 ( .B(n501), .A(n502), .S(n371), .Y(n481) );
  MUX2X1 U448 ( .B(n503), .A(n504), .S(n371), .Y(n484) );
  MUX2X1 U449 ( .B(n473), .A(n483), .S(n373), .Y(n424) );
  MUX2X1 U450 ( .B(n505), .A(n506), .S(n371), .Y(n483) );
  MUX2X1 U451 ( .B(n507), .A(n508), .S(n371), .Y(n473) );
  MUX2X1 U452 ( .B(n392), .A(n363), .S(n378), .Y(B[12]) );
  AND2X1 U453 ( .A(n509), .B(n374), .Y(n467) );
  MUX2X1 U454 ( .B(n430), .A(n468), .S(n375), .Y(n510) );
  MUX2X1 U455 ( .B(n511), .A(n512), .S(n373), .Y(n468) );
  MUX2X1 U456 ( .B(n513), .A(n514), .S(n373), .Y(n430) );
  MUX2X1 U457 ( .B(n391), .A(n457), .S(n378), .Y(B[11]) );
  OR2X1 U458 ( .A(n478), .B(n376), .Y(n457) );
  MUX2X1 U459 ( .B(n489), .A(n360), .S(n373), .Y(n478) );
  MUX2X1 U460 ( .B(n499), .A(n501), .S(n371), .Y(n489) );
  MUX2X1 U461 ( .B(A[27]), .A(A[28]), .S(n367), .Y(n501) );
  MUX2X1 U462 ( .B(A[29]), .A(A[30]), .S(n367), .Y(n499) );
  MUX2X1 U463 ( .B(n437), .A(n477), .S(n375), .Y(n515) );
  MUX2X1 U464 ( .B(n491), .A(n488), .S(n373), .Y(n477) );
  MUX2X1 U465 ( .B(n502), .A(n503), .S(n371), .Y(n488) );
  MUX2X1 U466 ( .B(A[23]), .A(A[24]), .S(n367), .Y(n503) );
  MUX2X1 U467 ( .B(A[25]), .A(A[26]), .S(n367), .Y(n502) );
  MUX2X1 U468 ( .B(n504), .A(n505), .S(n371), .Y(n491) );
  MUX2X1 U469 ( .B(A[19]), .A(A[20]), .S(n367), .Y(n505) );
  MUX2X1 U470 ( .B(A[21]), .A(A[22]), .S(n367), .Y(n504) );
  MUX2X1 U471 ( .B(n414), .A(n490), .S(n373), .Y(n437) );
  MUX2X1 U472 ( .B(n506), .A(n507), .S(n371), .Y(n490) );
  MUX2X1 U473 ( .B(A[15]), .A(A[16]), .S(n367), .Y(n507) );
  MUX2X1 U474 ( .B(A[17]), .A(A[18]), .S(SH[0]), .Y(n506) );
  MUX2X1 U475 ( .B(n474), .A(n508), .S(n369), .Y(n414) );
  MUX2X1 U476 ( .B(A[13]), .A(A[14]), .S(SH[0]), .Y(n508) );
  MUX2X1 U477 ( .B(A[11]), .A(A[12]), .S(SH[0]), .Y(n474) );
  MUX2X1 U478 ( .B(n390), .A(n458), .S(n378), .Y(B[10]) );
  OR2X1 U479 ( .A(n480), .B(n376), .Y(n458) );
  MUX2X1 U480 ( .B(n495), .A(n365), .S(n373), .Y(n480) );
  MUX2X1 U481 ( .B(n517), .A(n518), .S(n371), .Y(n495) );
  MUX2X1 U482 ( .B(n449), .A(n479), .S(n375), .Y(n519) );
  MUX2X1 U483 ( .B(n497), .A(n494), .S(n373), .Y(n479) );
  MUX2X1 U484 ( .B(n520), .A(n521), .S(n371), .Y(n494) );
  MUX2X1 U485 ( .B(n522), .A(n523), .S(n371), .Y(n497) );
  MUX2X1 U486 ( .B(n420), .A(n496), .S(n373), .Y(n449) );
  MUX2X1 U487 ( .B(n524), .A(n525), .S(n372), .Y(n496) );
  MUX2X1 U488 ( .B(n526), .A(n527), .S(n369), .Y(n420) );
  MUX2X1 U489 ( .B(n529), .A(n485), .S(n378), .Y(n528) );
  MUX2X1 U490 ( .B(n460), .A(n408), .S(n377), .Y(n485) );
  MUX2X1 U491 ( .B(n514), .A(n511), .S(n373), .Y(n408) );
  MUX2X1 U492 ( .B(n521), .A(n522), .S(n372), .Y(n511) );
  MUX2X1 U493 ( .B(A[20]), .A(A[21]), .S(SH[0]), .Y(n522) );
  MUX2X1 U494 ( .B(A[22]), .A(A[23]), .S(SH[0]), .Y(n521) );
  MUX2X1 U495 ( .B(n523), .A(n524), .S(n372), .Y(n514) );
  MUX2X1 U496 ( .B(A[16]), .A(A[17]), .S(SH[0]), .Y(n524) );
  MUX2X1 U497 ( .B(A[18]), .A(A[19]), .S(SH[0]), .Y(n523) );
  MUX2X1 U498 ( .B(n512), .A(n509), .S(n373), .Y(n460) );
  MUX2X1 U499 ( .B(n516), .A(n517), .S(n372), .Y(n509) );
  MUX2X1 U500 ( .B(A[28]), .A(A[29]), .S(SH[0]), .Y(n517) );
  MUX2X1 U501 ( .B(A[30]), .A(A[31]), .S(SH[0]), .Y(n516) );
  MUX2X1 U502 ( .B(n518), .A(n520), .S(n372), .Y(n512) );
  MUX2X1 U503 ( .B(A[24]), .A(A[25]), .S(SH[0]), .Y(n520) );
  MUX2X1 U504 ( .B(A[26]), .A(A[27]), .S(SH[0]), .Y(n518) );
  MUX2X1 U505 ( .B(n530), .A(n407), .S(n376), .Y(n529) );
  MUX2X1 U506 ( .B(n432), .A(n513), .S(n373), .Y(n407) );
  MUX2X1 U507 ( .B(n525), .A(n527), .S(n372), .Y(n513) );
  MUX2X1 U508 ( .B(A[12]), .A(A[13]), .S(SH[0]), .Y(n527) );
  MUX2X1 U509 ( .B(A[14]), .A(A[15]), .S(n367), .Y(n525) );
  MUX2X1 U510 ( .B(n452), .A(n526), .S(n369), .Y(n432) );
  MUX2X1 U511 ( .B(A[10]), .A(A[11]), .S(n367), .Y(n526) );
  MUX2X1 U512 ( .B(A[8]), .A(A[9]), .S(n367), .Y(n452) );
  MUX2X1 U513 ( .B(n531), .A(n431), .S(n373), .Y(n530) );
  MUX2X1 U514 ( .B(n454), .A(n451), .S(n369), .Y(n431) );
  MUX2X1 U515 ( .B(A[6]), .A(A[7]), .S(n367), .Y(n451) );
  MUX2X1 U516 ( .B(A[4]), .A(A[5]), .S(n367), .Y(n454) );
  MUX2X1 U517 ( .B(n532), .A(n453), .S(n369), .Y(n531) );
  MUX2X1 U518 ( .B(A[2]), .A(A[3]), .S(SH[0]), .Y(n453) );
  MUX2X1 U519 ( .B(A[0]), .A(A[1]), .S(SH[0]), .Y(n532) );
endmodule


module alu_DW_rightsh_45 ( A, DATA_TC, SH, B );
  input [63:0] A;
  input [5:0] SH;
  output [63:0] B;
  input DATA_TC;
  wire   n1245, n1244, n1243, n1242, n1241, n1240, n1239, n1238, n1237, n1236,
         n1235, n1234, n1233, n1232, n1231, n1230, n1229, n1228, n1227, n1226,
         n1225, n1224, n1223, n1222, n1221, n1220, n1219, n1218, n1217, n1216,
         n1215, n1214, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n845, n846, n849, n850, n852, n853, n854, n858,
         n859, n860, n864, n865, n866, n867, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213;

  AND2X1 U739 ( .A(n839), .B(n889), .Y(n934) );
  OR2X1 U740 ( .A(n891), .B(n831), .Y(n1214) );
  INVX1 U741 ( .A(n1214), .Y(B[63]) );
  OR2X1 U742 ( .A(n890), .B(n832), .Y(n1215) );
  INVX1 U743 ( .A(n1215), .Y(B[62]) );
  OR2X1 U744 ( .A(n835), .B(n892), .Y(n1216) );
  INVX1 U745 ( .A(n1216), .Y(B[61]) );
  OR2X1 U746 ( .A(n837), .B(n892), .Y(n1217) );
  INVX1 U747 ( .A(n1217), .Y(B[60]) );
  OR2X1 U748 ( .A(n836), .B(n892), .Y(n1219) );
  INVX1 U749 ( .A(n1219), .Y(B[58]) );
  OR2X1 U750 ( .A(n838), .B(n892), .Y(n1220) );
  INVX1 U751 ( .A(n1220), .Y(B[57]) );
  OR2X1 U752 ( .A(n833), .B(n892), .Y(n1224) );
  INVX1 U753 ( .A(n1224), .Y(B[53]) );
  OR2X1 U754 ( .A(n842), .B(n892), .Y(n1225) );
  INVX1 U755 ( .A(n1225), .Y(B[52]) );
  OR2X1 U756 ( .A(n834), .B(n891), .Y(n1227) );
  INVX1 U757 ( .A(n1227), .Y(B[50]) );
  OR2X1 U758 ( .A(n840), .B(n892), .Y(n1228) );
  INVX1 U759 ( .A(n1228), .Y(B[49]) );
  OR2X1 U760 ( .A(n892), .B(n954), .Y(n1230) );
  INVX1 U761 ( .A(n1230), .Y(B[47]) );
  OR2X1 U762 ( .A(n892), .B(n956), .Y(n1232) );
  INVX1 U763 ( .A(n1232), .Y(B[45]) );
  OR2X1 U764 ( .A(n892), .B(n957), .Y(n1233) );
  INVX1 U765 ( .A(n1233), .Y(B[44]) );
  OR2X1 U766 ( .A(n892), .B(n958), .Y(n1234) );
  INVX1 U767 ( .A(n1234), .Y(B[43]) );
  OR2X1 U768 ( .A(n892), .B(n959), .Y(n1235) );
  INVX1 U769 ( .A(n1235), .Y(B[42]) );
  OR2X1 U770 ( .A(n892), .B(n895), .Y(n1236) );
  INVX1 U771 ( .A(n1236), .Y(B[41]) );
  OR2X1 U772 ( .A(n892), .B(n985), .Y(n1243) );
  INVX1 U773 ( .A(n1243), .Y(B[34]) );
  OR2X1 U774 ( .A(n850), .B(n892), .Y(n1222) );
  INVX1 U775 ( .A(n1222), .Y(B[55]) );
  OR2X1 U776 ( .A(n846), .B(n892), .Y(n1223) );
  INVX1 U777 ( .A(n1223), .Y(B[54]) );
  AND2X1 U778 ( .A(n845), .B(n889), .Y(n922) );
  INVX1 U779 ( .A(n922), .Y(n831) );
  AND2X1 U780 ( .A(n858), .B(n889), .Y(n923) );
  INVX1 U781 ( .A(n923), .Y(n832) );
  AND2X1 U782 ( .A(n979), .B(n889), .Y(n940) );
  INVX1 U783 ( .A(n940), .Y(n833) );
  AND2X1 U784 ( .A(n997), .B(n889), .Y(n943) );
  INVX1 U785 ( .A(n943), .Y(n834) );
  AND2X1 U786 ( .A(n841), .B(n889), .Y(n924) );
  INVX1 U787 ( .A(n924), .Y(n835) );
  AND2X1 U788 ( .A(n849), .B(n889), .Y(n935) );
  INVX1 U789 ( .A(n935), .Y(n836) );
  AND2X1 U790 ( .A(n852), .B(n889), .Y(n925) );
  INVX1 U791 ( .A(n925), .Y(n837) );
  AND2X1 U792 ( .A(n864), .B(n889), .Y(n936) );
  INVX1 U793 ( .A(n936), .Y(n838) );
  OR2X1 U794 ( .A(n1076), .B(n888), .Y(n1017) );
  INVX1 U795 ( .A(n1017), .Y(n839) );
  AND2X1 U796 ( .A(n1065), .B(n889), .Y(n952) );
  INVX1 U797 ( .A(n952), .Y(n840) );
  OR2X1 U798 ( .A(n859), .B(n888), .Y(n1009) );
  INVX1 U799 ( .A(n1009), .Y(n841) );
  AND2X1 U800 ( .A(n981), .B(n889), .Y(n941) );
  INVX1 U801 ( .A(n941), .Y(n842) );
  OR2X1 U802 ( .A(n945), .B(n891), .Y(n1241) );
  INVX1 U803 ( .A(n1241), .Y(B[36]) );
  OR2X1 U804 ( .A(n854), .B(n892), .Y(n1221) );
  INVX1 U805 ( .A(n1221), .Y(B[56]) );
  OR2X1 U806 ( .A(n853), .B(n887), .Y(n989) );
  INVX1 U807 ( .A(n989), .Y(n845) );
  AND2X1 U808 ( .A(n977), .B(n889), .Y(n939) );
  INVX1 U809 ( .A(n939), .Y(n846) );
  OR2X1 U810 ( .A(n986), .B(n891), .Y(n1244) );
  INVX1 U811 ( .A(n1244), .Y(B[33]) );
  OR2X1 U812 ( .A(n892), .B(n955), .Y(n1231) );
  INVX1 U813 ( .A(n1231), .Y(B[46]) );
  OR2X1 U814 ( .A(n1083), .B(n888), .Y(n1021) );
  INVX1 U815 ( .A(n1021), .Y(n849) );
  AND2X1 U816 ( .A(n975), .B(n889), .Y(n938) );
  INVX1 U817 ( .A(n938), .Y(n850) );
  OR2X1 U818 ( .A(n860), .B(n891), .Y(n1229) );
  INVX1 U819 ( .A(n1229), .Y(B[48]) );
  OR2X1 U820 ( .A(n872), .B(n888), .Y(n1013) );
  INVX1 U821 ( .A(n1013), .Y(n852) );
  AND2X1 U822 ( .A(n865), .B(n882), .Y(n1038) );
  INVX1 U823 ( .A(n1038), .Y(n853) );
  AND2X1 U824 ( .A(n871), .B(n889), .Y(n937) );
  INVX1 U825 ( .A(n937), .Y(n854) );
  OR2X1 U826 ( .A(n892), .B(n965), .Y(n1242) );
  INVX1 U827 ( .A(n1242), .Y(B[35]) );
  OR2X1 U828 ( .A(n891), .B(n867), .Y(n1218) );
  INVX1 U829 ( .A(n1218), .Y(B[59]) );
  OR2X1 U830 ( .A(n907), .B(n890), .Y(n1238) );
  INVX1 U831 ( .A(n1238), .Y(B[39]) );
  OR2X1 U832 ( .A(n866), .B(n887), .Y(n993) );
  INVX1 U833 ( .A(n993), .Y(n858) );
  AND2X1 U834 ( .A(n1089), .B(n883), .Y(n1052) );
  INVX1 U835 ( .A(n1052), .Y(n859) );
  AND2X1 U836 ( .A(n1102), .B(n889), .Y(n953) );
  INVX1 U837 ( .A(n953), .Y(n860) );
  OR2X1 U838 ( .A(n892), .B(n874), .Y(n1226) );
  INVX1 U839 ( .A(n1226), .Y(B[51]) );
  OR2X1 U840 ( .A(n915), .B(n890), .Y(n1239) );
  INVX1 U841 ( .A(n1239), .Y(B[38]) );
  OR2X1 U842 ( .A(n892), .B(n901), .Y(n1237) );
  INVX1 U843 ( .A(n1237), .Y(B[40]) );
  OR2X1 U844 ( .A(n1025), .B(n888), .Y(n960) );
  INVX1 U845 ( .A(n960), .Y(n864) );
  OR2X1 U846 ( .A(n873), .B(SH[1]), .Y(n1110) );
  INVX1 U847 ( .A(n1110), .Y(n865) );
  AND2X1 U848 ( .A(n870), .B(n884), .Y(n1045) );
  INVX1 U849 ( .A(n1045), .Y(n866) );
  INVX1 U850 ( .A(n934), .Y(n867) );
  OR2X1 U851 ( .A(n892), .B(n987), .Y(n1245) );
  INVX1 U852 ( .A(n1245), .Y(B[32]) );
  OR2X1 U853 ( .A(n927), .B(n891), .Y(n1240) );
  INVX1 U854 ( .A(n1240), .Y(B[37]) );
  OR2X1 U855 ( .A(n1191), .B(n878), .Y(n1125) );
  INVX1 U856 ( .A(n1125), .Y(n870) );
  OR2X1 U857 ( .A(n1031), .B(n888), .Y(n962) );
  INVX1 U858 ( .A(n962), .Y(n871) );
  AND2X1 U859 ( .A(n1168), .B(n883), .Y(n1059) );
  INVX1 U860 ( .A(n1059), .Y(n872) );
  AND2X1 U861 ( .A(A[63]), .B(n875), .Y(n1145) );
  INVX1 U862 ( .A(n1145), .Y(n873) );
  AND2X1 U863 ( .A(n983), .B(n889), .Y(n942) );
  INVX1 U864 ( .A(n942), .Y(n874) );
  INVX1 U865 ( .A(n885), .Y(n886) );
  INVX1 U866 ( .A(n885), .Y(n888) );
  INVX1 U867 ( .A(n885), .Y(n887) );
  INVX1 U868 ( .A(SH[0]), .Y(n876) );
  INVX1 U869 ( .A(n881), .Y(n884) );
  INVX1 U870 ( .A(n881), .Y(n883) );
  INVX1 U871 ( .A(SH[4]), .Y(n889) );
  INVX1 U872 ( .A(n880), .Y(n877) );
  INVX1 U873 ( .A(n880), .Y(n878) );
  INVX1 U874 ( .A(n880), .Y(n879) );
  INVX1 U875 ( .A(n882), .Y(n881) );
  INVX1 U876 ( .A(SH[0]), .Y(n875) );
  INVX1 U877 ( .A(SH[1]), .Y(n880) );
  INVX1 U878 ( .A(SH[2]), .Y(n882) );
  INVX1 U879 ( .A(SH[3]), .Y(n885) );
  INVX1 U880 ( .A(n893), .Y(n892) );
  INVX1 U881 ( .A(n893), .Y(n891) );
  INVX1 U882 ( .A(n893), .Y(n890) );
  INVX1 U883 ( .A(SH[5]), .Y(n893) );
  MUX2X1 U884 ( .B(n894), .A(n895), .S(n890), .Y(B[9]) );
  MUX2X1 U885 ( .B(n896), .A(n897), .S(n889), .Y(n894) );
  MUX2X1 U886 ( .B(n898), .A(n899), .S(n885), .Y(n897) );
  MUX2X1 U887 ( .B(n900), .A(n901), .S(n890), .Y(B[8]) );
  MUX2X1 U888 ( .B(n902), .A(n903), .S(n889), .Y(n900) );
  MUX2X1 U889 ( .B(n904), .A(n905), .S(n885), .Y(n903) );
  MUX2X1 U890 ( .B(n906), .A(n907), .S(n890), .Y(B[7]) );
  MUX2X1 U891 ( .B(n908), .A(n909), .S(n889), .Y(n906) );
  MUX2X1 U892 ( .B(n910), .A(n911), .S(n885), .Y(n909) );
  MUX2X1 U893 ( .B(n912), .A(n913), .S(n883), .Y(n911) );
  MUX2X1 U894 ( .B(n914), .A(n915), .S(n890), .Y(B[6]) );
  MUX2X1 U895 ( .B(n916), .A(n917), .S(n889), .Y(n914) );
  MUX2X1 U896 ( .B(n918), .A(n919), .S(n885), .Y(n917) );
  MUX2X1 U897 ( .B(n920), .A(n921), .S(n882), .Y(n919) );
  MUX2X1 U898 ( .B(n926), .A(n927), .S(n891), .Y(B[5]) );
  MUX2X1 U899 ( .B(n928), .A(n929), .S(n889), .Y(n926) );
  MUX2X1 U900 ( .B(n930), .A(n931), .S(n885), .Y(n929) );
  MUX2X1 U901 ( .B(n932), .A(n933), .S(n882), .Y(n931) );
  MUX2X1 U902 ( .B(n944), .A(n945), .S(n890), .Y(B[4]) );
  MUX2X1 U903 ( .B(n946), .A(n947), .S(n889), .Y(n944) );
  MUX2X1 U904 ( .B(n948), .A(n949), .S(n885), .Y(n947) );
  MUX2X1 U905 ( .B(n950), .A(n951), .S(n882), .Y(n949) );
  MUX2X1 U906 ( .B(n864), .A(n961), .S(n889), .Y(n895) );
  MUX2X1 U907 ( .B(n871), .A(n963), .S(n889), .Y(n901) );
  MUX2X1 U908 ( .B(n964), .A(n965), .S(n890), .Y(B[3]) );
  MUX2X1 U909 ( .B(n966), .A(n967), .S(n889), .Y(n964) );
  MUX2X1 U910 ( .B(n968), .A(n969), .S(n885), .Y(n967) );
  MUX2X1 U911 ( .B(n913), .A(n970), .S(n882), .Y(n969) );
  MUX2X1 U912 ( .B(n971), .A(n972), .S(SH[1]), .Y(n970) );
  MUX2X1 U913 ( .B(n973), .A(n974), .S(n879), .Y(n913) );
  MUX2X1 U914 ( .B(n975), .A(n976), .S(n889), .Y(n907) );
  MUX2X1 U915 ( .B(n977), .A(n978), .S(n889), .Y(n915) );
  MUX2X1 U916 ( .B(n979), .A(n980), .S(n889), .Y(n927) );
  MUX2X1 U917 ( .B(n981), .A(n982), .S(n889), .Y(n945) );
  MUX2X1 U918 ( .B(n983), .A(n984), .S(n889), .Y(n965) );
  MUX2X1 U919 ( .B(n988), .A(n831), .S(n890), .Y(B[31]) );
  MUX2X1 U920 ( .B(n990), .A(n991), .S(n889), .Y(n988) );
  MUX2X1 U921 ( .B(n992), .A(n832), .S(n890), .Y(B[30]) );
  MUX2X1 U922 ( .B(n994), .A(n995), .S(n889), .Y(n992) );
  MUX2X1 U923 ( .B(n996), .A(n985), .S(n890), .Y(B[2]) );
  MUX2X1 U924 ( .B(n997), .A(n998), .S(n889), .Y(n985) );
  MUX2X1 U925 ( .B(n999), .A(n1000), .S(n889), .Y(n996) );
  MUX2X1 U926 ( .B(n1001), .A(n1002), .S(n885), .Y(n1000) );
  MUX2X1 U927 ( .B(n921), .A(n1003), .S(n882), .Y(n1002) );
  MUX2X1 U928 ( .B(n1004), .A(n1005), .S(n879), .Y(n1003) );
  MUX2X1 U929 ( .B(n1006), .A(n1007), .S(n879), .Y(n921) );
  MUX2X1 U930 ( .B(n1008), .A(n835), .S(n890), .Y(B[29]) );
  MUX2X1 U931 ( .B(n1010), .A(n1011), .S(n889), .Y(n1008) );
  MUX2X1 U932 ( .B(n1012), .A(n837), .S(n890), .Y(B[28]) );
  MUX2X1 U933 ( .B(n1014), .A(n1015), .S(n889), .Y(n1012) );
  MUX2X1 U934 ( .B(n1016), .A(n867), .S(n891), .Y(B[27]) );
  MUX2X1 U935 ( .B(n1018), .A(n1019), .S(n889), .Y(n1016) );
  MUX2X1 U936 ( .B(n1020), .A(n836), .S(n891), .Y(B[26]) );
  MUX2X1 U937 ( .B(n1022), .A(n1023), .S(n889), .Y(n1020) );
  MUX2X1 U938 ( .B(n1024), .A(n838), .S(n891), .Y(B[25]) );
  MUX2X1 U939 ( .B(n961), .A(n896), .S(n889), .Y(n1024) );
  MUX2X1 U940 ( .B(n1026), .A(n1027), .S(n888), .Y(n896) );
  MUX2X1 U941 ( .B(n1028), .A(n1029), .S(n888), .Y(n961) );
  MUX2X1 U942 ( .B(n1030), .A(n854), .S(n891), .Y(B[24]) );
  MUX2X1 U943 ( .B(n963), .A(n902), .S(n889), .Y(n1030) );
  MUX2X1 U944 ( .B(n1032), .A(n1033), .S(n888), .Y(n902) );
  MUX2X1 U945 ( .B(n1034), .A(n1035), .S(n887), .Y(n963) );
  MUX2X1 U946 ( .B(n1036), .A(n850), .S(n891), .Y(B[23]) );
  MUX2X1 U947 ( .B(n1037), .A(n853), .S(n888), .Y(n975) );
  MUX2X1 U948 ( .B(n976), .A(n908), .S(n889), .Y(n1036) );
  MUX2X1 U949 ( .B(n1039), .A(n1040), .S(n888), .Y(n908) );
  MUX2X1 U950 ( .B(n1041), .A(n1042), .S(n888), .Y(n976) );
  MUX2X1 U951 ( .B(n1043), .A(n846), .S(n891), .Y(B[22]) );
  MUX2X1 U952 ( .B(n1044), .A(n866), .S(n888), .Y(n977) );
  MUX2X1 U953 ( .B(n978), .A(n916), .S(n889), .Y(n1043) );
  MUX2X1 U954 ( .B(n1046), .A(n1047), .S(n888), .Y(n916) );
  MUX2X1 U955 ( .B(n1048), .A(n1049), .S(n888), .Y(n978) );
  MUX2X1 U956 ( .B(n1050), .A(n833), .S(n891), .Y(B[21]) );
  MUX2X1 U957 ( .B(n1051), .A(n859), .S(n888), .Y(n979) );
  MUX2X1 U958 ( .B(n980), .A(n928), .S(n889), .Y(n1050) );
  MUX2X1 U959 ( .B(n1053), .A(n1054), .S(n888), .Y(n928) );
  MUX2X1 U960 ( .B(n1055), .A(n1056), .S(n888), .Y(n980) );
  MUX2X1 U961 ( .B(n1057), .A(n842), .S(n891), .Y(B[20]) );
  MUX2X1 U962 ( .B(n1058), .A(n872), .S(n888), .Y(n981) );
  MUX2X1 U963 ( .B(n982), .A(n946), .S(n889), .Y(n1057) );
  MUX2X1 U964 ( .B(n1060), .A(n1061), .S(n888), .Y(n946) );
  MUX2X1 U965 ( .B(n1062), .A(n1063), .S(n888), .Y(n982) );
  MUX2X1 U966 ( .B(n1064), .A(n986), .S(n891), .Y(B[1]) );
  MUX2X1 U967 ( .B(n1065), .A(n1066), .S(n889), .Y(n986) );
  MUX2X1 U968 ( .B(n1067), .A(n1068), .S(n889), .Y(n1064) );
  MUX2X1 U969 ( .B(n899), .A(n1069), .S(n885), .Y(n1068) );
  MUX2X1 U970 ( .B(n933), .A(n1070), .S(n882), .Y(n1069) );
  MUX2X1 U971 ( .B(n1071), .A(n971), .S(n878), .Y(n1070) );
  MUX2X1 U972 ( .B(A[4]), .A(A[3]), .S(n876), .Y(n971) );
  MUX2X1 U973 ( .B(A[2]), .A(A[1]), .S(n876), .Y(n1071) );
  MUX2X1 U974 ( .B(n972), .A(n973), .S(n878), .Y(n933) );
  MUX2X1 U975 ( .B(A[8]), .A(A[7]), .S(n875), .Y(n973) );
  MUX2X1 U976 ( .B(A[6]), .A(A[5]), .S(n876), .Y(n972) );
  MUX2X1 U977 ( .B(n1072), .A(n932), .S(n884), .Y(n899) );
  MUX2X1 U978 ( .B(n974), .A(n1073), .S(n879), .Y(n932) );
  MUX2X1 U979 ( .B(A[10]), .A(A[9]), .S(n875), .Y(n974) );
  MUX2X1 U980 ( .B(n1074), .A(n874), .S(n891), .Y(B[19]) );
  MUX2X1 U981 ( .B(n1075), .A(n1076), .S(n887), .Y(n983) );
  MUX2X1 U982 ( .B(n984), .A(n966), .S(n889), .Y(n1074) );
  MUX2X1 U983 ( .B(n1077), .A(n1078), .S(n887), .Y(n966) );
  MUX2X1 U984 ( .B(n1079), .A(n1080), .S(n887), .Y(n984) );
  MUX2X1 U985 ( .B(n1081), .A(n834), .S(n891), .Y(B[18]) );
  MUX2X1 U986 ( .B(n1082), .A(n1083), .S(n887), .Y(n997) );
  MUX2X1 U987 ( .B(n998), .A(n999), .S(n889), .Y(n1081) );
  MUX2X1 U988 ( .B(n1084), .A(n1085), .S(n887), .Y(n999) );
  MUX2X1 U989 ( .B(n1086), .A(n1087), .S(n887), .Y(n998) );
  MUX2X1 U990 ( .B(n1088), .A(n840), .S(n891), .Y(B[17]) );
  MUX2X1 U991 ( .B(n1029), .A(n1025), .S(n887), .Y(n1065) );
  MUX2X1 U992 ( .B(n1089), .A(n1090), .S(n884), .Y(n1025) );
  MUX2X1 U993 ( .B(n1091), .A(n1092), .S(n882), .Y(n1029) );
  MUX2X1 U994 ( .B(n1066), .A(n1067), .S(n889), .Y(n1088) );
  MUX2X1 U995 ( .B(n898), .A(n1026), .S(n887), .Y(n1067) );
  MUX2X1 U996 ( .B(n1093), .A(n1094), .S(n882), .Y(n1026) );
  MUX2X1 U997 ( .B(n1095), .A(n1096), .S(n882), .Y(n898) );
  MUX2X1 U998 ( .B(n1027), .A(n1028), .S(n887), .Y(n1066) );
  MUX2X1 U999 ( .B(n1097), .A(n1098), .S(n882), .Y(n1028) );
  MUX2X1 U1000 ( .B(n1099), .A(n1100), .S(n884), .Y(n1027) );
  MUX2X1 U1001 ( .B(n1101), .A(n860), .S(n891), .Y(B[16]) );
  MUX2X1 U1002 ( .B(n1103), .A(n1104), .S(n889), .Y(n1101) );
  MUX2X1 U1003 ( .B(n1105), .A(n954), .S(n891), .Y(B[15]) );
  MUX2X1 U1004 ( .B(n845), .A(n990), .S(n889), .Y(n954) );
  MUX2X1 U1005 ( .B(n1042), .A(n1037), .S(n887), .Y(n990) );
  MUX2X1 U1006 ( .B(n1106), .A(n1107), .S(n882), .Y(n1037) );
  MUX2X1 U1007 ( .B(n1108), .A(n1109), .S(n882), .Y(n1042) );
  MUX2X1 U1008 ( .B(n991), .A(n1111), .S(n889), .Y(n1105) );
  MUX2X1 U1009 ( .B(n1039), .A(n910), .S(n885), .Y(n1111) );
  MUX2X1 U1010 ( .B(n1112), .A(n1113), .S(n882), .Y(n910) );
  MUX2X1 U1011 ( .B(n1114), .A(n1115), .S(n882), .Y(n1039) );
  MUX2X1 U1012 ( .B(n1040), .A(n1041), .S(n887), .Y(n991) );
  MUX2X1 U1013 ( .B(n1116), .A(n1117), .S(n882), .Y(n1041) );
  MUX2X1 U1014 ( .B(n1118), .A(n1119), .S(n882), .Y(n1040) );
  MUX2X1 U1015 ( .B(n1120), .A(n955), .S(n890), .Y(B[14]) );
  MUX2X1 U1016 ( .B(n858), .A(n994), .S(n889), .Y(n955) );
  MUX2X1 U1017 ( .B(n1049), .A(n1044), .S(n886), .Y(n994) );
  MUX2X1 U1018 ( .B(n1121), .A(n1122), .S(n884), .Y(n1044) );
  MUX2X1 U1019 ( .B(n1123), .A(n1124), .S(n884), .Y(n1049) );
  MUX2X1 U1020 ( .B(n995), .A(n1126), .S(n889), .Y(n1120) );
  MUX2X1 U1021 ( .B(n1046), .A(n918), .S(n885), .Y(n1126) );
  MUX2X1 U1022 ( .B(n1127), .A(n1128), .S(n884), .Y(n918) );
  MUX2X1 U1023 ( .B(n1129), .A(n1130), .S(n884), .Y(n1046) );
  MUX2X1 U1024 ( .B(n1047), .A(n1048), .S(n886), .Y(n995) );
  MUX2X1 U1025 ( .B(n1131), .A(n1132), .S(n884), .Y(n1048) );
  MUX2X1 U1026 ( .B(n1133), .A(n1134), .S(n884), .Y(n1047) );
  MUX2X1 U1027 ( .B(n1135), .A(n956), .S(n891), .Y(B[13]) );
  MUX2X1 U1028 ( .B(n841), .A(n1010), .S(n889), .Y(n956) );
  MUX2X1 U1029 ( .B(n1056), .A(n1051), .S(n886), .Y(n1010) );
  MUX2X1 U1030 ( .B(n1090), .A(n1091), .S(n884), .Y(n1051) );
  MUX2X1 U1031 ( .B(n1136), .A(n1137), .S(n879), .Y(n1091) );
  MUX2X1 U1032 ( .B(n1138), .A(n1139), .S(n879), .Y(n1090) );
  MUX2X1 U1033 ( .B(n1092), .A(n1097), .S(n884), .Y(n1056) );
  MUX2X1 U1034 ( .B(n1140), .A(n1141), .S(n879), .Y(n1097) );
  MUX2X1 U1035 ( .B(n1142), .A(n1143), .S(n879), .Y(n1092) );
  MUX2X1 U1036 ( .B(n1144), .A(n873), .S(n879), .Y(n1089) );
  MUX2X1 U1037 ( .B(n1011), .A(n1146), .S(n889), .Y(n1135) );
  MUX2X1 U1038 ( .B(n1053), .A(n930), .S(n885), .Y(n1146) );
  MUX2X1 U1039 ( .B(n1096), .A(n1072), .S(n884), .Y(n930) );
  MUX2X1 U1040 ( .B(n1147), .A(n1148), .S(n877), .Y(n1072) );
  MUX2X1 U1041 ( .B(n1149), .A(n1150), .S(n877), .Y(n1096) );
  MUX2X1 U1042 ( .B(n1094), .A(n1095), .S(n884), .Y(n1053) );
  MUX2X1 U1043 ( .B(n1151), .A(n1152), .S(n877), .Y(n1095) );
  MUX2X1 U1044 ( .B(n1153), .A(n1154), .S(n877), .Y(n1094) );
  MUX2X1 U1045 ( .B(n1054), .A(n1055), .S(n886), .Y(n1011) );
  MUX2X1 U1046 ( .B(n1098), .A(n1099), .S(n884), .Y(n1055) );
  MUX2X1 U1047 ( .B(n1155), .A(n1156), .S(n877), .Y(n1099) );
  MUX2X1 U1048 ( .B(n1157), .A(n1158), .S(n877), .Y(n1098) );
  MUX2X1 U1049 ( .B(n1100), .A(n1093), .S(n884), .Y(n1054) );
  MUX2X1 U1050 ( .B(n1159), .A(n1160), .S(n877), .Y(n1093) );
  MUX2X1 U1051 ( .B(n1161), .A(n1162), .S(n877), .Y(n1100) );
  MUX2X1 U1052 ( .B(n1163), .A(n957), .S(n890), .Y(B[12]) );
  MUX2X1 U1053 ( .B(n852), .A(n1014), .S(n889), .Y(n957) );
  MUX2X1 U1054 ( .B(n1063), .A(n1058), .S(n886), .Y(n1014) );
  MUX2X1 U1055 ( .B(n1164), .A(n1165), .S(n884), .Y(n1058) );
  MUX2X1 U1056 ( .B(n1166), .A(n1167), .S(n884), .Y(n1063) );
  MUX2X1 U1057 ( .B(n1015), .A(n1169), .S(n889), .Y(n1163) );
  MUX2X1 U1058 ( .B(n1060), .A(n948), .S(n885), .Y(n1169) );
  MUX2X1 U1059 ( .B(n1170), .A(n1171), .S(n884), .Y(n948) );
  MUX2X1 U1060 ( .B(n1172), .A(n1173), .S(n884), .Y(n1060) );
  MUX2X1 U1061 ( .B(n1061), .A(n1062), .S(n886), .Y(n1015) );
  MUX2X1 U1062 ( .B(n1174), .A(n1175), .S(n883), .Y(n1062) );
  MUX2X1 U1063 ( .B(n1176), .A(n1177), .S(n883), .Y(n1061) );
  MUX2X1 U1064 ( .B(n1178), .A(n958), .S(n891), .Y(B[11]) );
  MUX2X1 U1065 ( .B(n839), .A(n1018), .S(n889), .Y(n958) );
  MUX2X1 U1066 ( .B(n1080), .A(n1075), .S(n886), .Y(n1018) );
  MUX2X1 U1067 ( .B(n1107), .A(n1108), .S(n883), .Y(n1075) );
  MUX2X1 U1068 ( .B(n1143), .A(n1136), .S(n877), .Y(n1108) );
  MUX2X1 U1069 ( .B(A[54]), .A(A[53]), .S(n875), .Y(n1136) );
  MUX2X1 U1070 ( .B(A[52]), .A(A[51]), .S(n875), .Y(n1143) );
  MUX2X1 U1071 ( .B(n1137), .A(n1138), .S(n877), .Y(n1107) );
  MUX2X1 U1072 ( .B(A[58]), .A(A[57]), .S(n875), .Y(n1138) );
  MUX2X1 U1073 ( .B(A[56]), .A(A[55]), .S(n875), .Y(n1137) );
  MUX2X1 U1074 ( .B(n1109), .A(n1116), .S(n883), .Y(n1080) );
  MUX2X1 U1075 ( .B(n1158), .A(n1140), .S(n877), .Y(n1116) );
  MUX2X1 U1076 ( .B(A[46]), .A(A[45]), .S(n875), .Y(n1140) );
  MUX2X1 U1077 ( .B(A[44]), .A(A[43]), .S(n876), .Y(n1158) );
  MUX2X1 U1078 ( .B(n1141), .A(n1142), .S(n877), .Y(n1109) );
  MUX2X1 U1079 ( .B(A[50]), .A(A[49]), .S(n875), .Y(n1142) );
  MUX2X1 U1080 ( .B(A[48]), .A(A[47]), .S(n875), .Y(n1141) );
  MUX2X1 U1081 ( .B(n865), .A(n1106), .S(n883), .Y(n1076) );
  MUX2X1 U1082 ( .B(n1139), .A(n1144), .S(SH[1]), .Y(n1106) );
  MUX2X1 U1083 ( .B(A[62]), .A(A[61]), .S(n875), .Y(n1144) );
  MUX2X1 U1084 ( .B(A[60]), .A(A[59]), .S(n875), .Y(n1139) );
  MUX2X1 U1085 ( .B(n1019), .A(n1179), .S(n889), .Y(n1178) );
  MUX2X1 U1086 ( .B(n1077), .A(n968), .S(n885), .Y(n1179) );
  MUX2X1 U1087 ( .B(n1113), .A(n912), .S(n883), .Y(n968) );
  MUX2X1 U1088 ( .B(n1073), .A(n1147), .S(SH[1]), .Y(n912) );
  MUX2X1 U1089 ( .B(A[14]), .A(A[13]), .S(n876), .Y(n1147) );
  MUX2X1 U1090 ( .B(A[12]), .A(A[11]), .S(n876), .Y(n1073) );
  MUX2X1 U1091 ( .B(n1148), .A(n1149), .S(SH[1]), .Y(n1113) );
  MUX2X1 U1092 ( .B(A[18]), .A(A[17]), .S(n876), .Y(n1149) );
  MUX2X1 U1093 ( .B(A[16]), .A(A[15]), .S(n875), .Y(n1148) );
  MUX2X1 U1094 ( .B(n1115), .A(n1112), .S(n883), .Y(n1077) );
  MUX2X1 U1095 ( .B(n1150), .A(n1151), .S(n879), .Y(n1112) );
  MUX2X1 U1096 ( .B(A[22]), .A(A[21]), .S(n876), .Y(n1151) );
  MUX2X1 U1097 ( .B(A[20]), .A(A[19]), .S(n875), .Y(n1150) );
  MUX2X1 U1098 ( .B(n1152), .A(n1153), .S(n878), .Y(n1115) );
  MUX2X1 U1099 ( .B(A[26]), .A(A[25]), .S(n875), .Y(n1153) );
  MUX2X1 U1100 ( .B(A[24]), .A(A[23]), .S(n876), .Y(n1152) );
  MUX2X1 U1101 ( .B(n1078), .A(n1079), .S(n886), .Y(n1019) );
  MUX2X1 U1102 ( .B(n1117), .A(n1118), .S(n883), .Y(n1079) );
  MUX2X1 U1103 ( .B(n1162), .A(n1155), .S(n879), .Y(n1118) );
  MUX2X1 U1104 ( .B(A[38]), .A(A[37]), .S(n876), .Y(n1155) );
  MUX2X1 U1105 ( .B(A[36]), .A(A[35]), .S(n875), .Y(n1162) );
  MUX2X1 U1106 ( .B(n1156), .A(n1157), .S(n878), .Y(n1117) );
  MUX2X1 U1107 ( .B(A[42]), .A(A[41]), .S(n876), .Y(n1157) );
  MUX2X1 U1108 ( .B(A[40]), .A(A[39]), .S(n875), .Y(n1156) );
  MUX2X1 U1109 ( .B(n1119), .A(n1114), .S(n883), .Y(n1078) );
  MUX2X1 U1110 ( .B(n1154), .A(n1159), .S(n878), .Y(n1114) );
  MUX2X1 U1111 ( .B(A[30]), .A(A[29]), .S(n875), .Y(n1159) );
  MUX2X1 U1112 ( .B(A[28]), .A(A[27]), .S(n876), .Y(n1154) );
  MUX2X1 U1113 ( .B(n1160), .A(n1161), .S(n878), .Y(n1119) );
  MUX2X1 U1114 ( .B(A[34]), .A(A[33]), .S(n876), .Y(n1161) );
  MUX2X1 U1115 ( .B(A[32]), .A(A[31]), .S(n876), .Y(n1160) );
  MUX2X1 U1116 ( .B(n1180), .A(n959), .S(n891), .Y(B[10]) );
  MUX2X1 U1117 ( .B(n849), .A(n1022), .S(n889), .Y(n959) );
  MUX2X1 U1118 ( .B(n1087), .A(n1082), .S(n886), .Y(n1022) );
  MUX2X1 U1119 ( .B(n1122), .A(n1123), .S(n883), .Y(n1082) );
  MUX2X1 U1120 ( .B(n1181), .A(n1182), .S(n878), .Y(n1123) );
  MUX2X1 U1121 ( .B(n1183), .A(n1184), .S(n878), .Y(n1122) );
  MUX2X1 U1122 ( .B(n1124), .A(n1131), .S(n883), .Y(n1087) );
  MUX2X1 U1123 ( .B(n1185), .A(n1186), .S(n878), .Y(n1131) );
  MUX2X1 U1124 ( .B(n1187), .A(n1188), .S(n878), .Y(n1124) );
  MUX2X1 U1125 ( .B(n870), .A(n1121), .S(n883), .Y(n1083) );
  MUX2X1 U1126 ( .B(n1189), .A(n1190), .S(n878), .Y(n1121) );
  MUX2X1 U1127 ( .B(n1023), .A(n1192), .S(n889), .Y(n1180) );
  MUX2X1 U1128 ( .B(n1084), .A(n1001), .S(n885), .Y(n1192) );
  MUX2X1 U1129 ( .B(n1128), .A(n920), .S(n883), .Y(n1001) );
  MUX2X1 U1130 ( .B(n1193), .A(n1194), .S(n878), .Y(n920) );
  MUX2X1 U1131 ( .B(n1195), .A(n1196), .S(n878), .Y(n1128) );
  MUX2X1 U1132 ( .B(n1130), .A(n1127), .S(n883), .Y(n1084) );
  MUX2X1 U1133 ( .B(n1197), .A(n1198), .S(n878), .Y(n1127) );
  MUX2X1 U1134 ( .B(n1199), .A(n1200), .S(n878), .Y(n1130) );
  MUX2X1 U1135 ( .B(n1085), .A(n1086), .S(n886), .Y(n1023) );
  MUX2X1 U1136 ( .B(n1132), .A(n1133), .S(n883), .Y(n1086) );
  MUX2X1 U1137 ( .B(n1201), .A(n1202), .S(n878), .Y(n1133) );
  MUX2X1 U1138 ( .B(n1203), .A(n1204), .S(n878), .Y(n1132) );
  MUX2X1 U1139 ( .B(n1134), .A(n1129), .S(n883), .Y(n1085) );
  MUX2X1 U1140 ( .B(n1205), .A(n1206), .S(n878), .Y(n1129) );
  MUX2X1 U1141 ( .B(n1207), .A(n1208), .S(n878), .Y(n1134) );
  MUX2X1 U1142 ( .B(n1209), .A(n987), .S(n890), .Y(B[0]) );
  MUX2X1 U1143 ( .B(n1102), .A(n1103), .S(n889), .Y(n987) );
  MUX2X1 U1144 ( .B(n1033), .A(n1034), .S(n886), .Y(n1103) );
  MUX2X1 U1145 ( .B(n1167), .A(n1174), .S(n883), .Y(n1034) );
  MUX2X1 U1146 ( .B(n1204), .A(n1185), .S(n878), .Y(n1174) );
  MUX2X1 U1147 ( .B(A[43]), .A(A[42]), .S(n876), .Y(n1185) );
  MUX2X1 U1148 ( .B(A[41]), .A(A[40]), .S(n876), .Y(n1204) );
  MUX2X1 U1149 ( .B(n1186), .A(n1187), .S(n879), .Y(n1167) );
  MUX2X1 U1150 ( .B(A[47]), .A(A[46]), .S(n876), .Y(n1187) );
  MUX2X1 U1151 ( .B(A[45]), .A(A[44]), .S(n876), .Y(n1186) );
  MUX2X1 U1152 ( .B(n1175), .A(n1176), .S(n883), .Y(n1033) );
  MUX2X1 U1153 ( .B(n1208), .A(n1201), .S(n879), .Y(n1176) );
  MUX2X1 U1154 ( .B(A[35]), .A(A[34]), .S(n876), .Y(n1201) );
  MUX2X1 U1155 ( .B(A[33]), .A(A[32]), .S(n876), .Y(n1208) );
  MUX2X1 U1156 ( .B(n1202), .A(n1203), .S(n879), .Y(n1175) );
  MUX2X1 U1157 ( .B(A[39]), .A(A[38]), .S(n876), .Y(n1203) );
  MUX2X1 U1158 ( .B(A[37]), .A(A[36]), .S(n876), .Y(n1202) );
  MUX2X1 U1159 ( .B(n1035), .A(n1031), .S(n886), .Y(n1102) );
  MUX2X1 U1160 ( .B(n1168), .A(n1164), .S(n883), .Y(n1031) );
  MUX2X1 U1161 ( .B(n1184), .A(n1189), .S(n879), .Y(n1164) );
  MUX2X1 U1162 ( .B(A[59]), .A(A[58]), .S(n875), .Y(n1189) );
  MUX2X1 U1163 ( .B(A[57]), .A(A[56]), .S(n876), .Y(n1184) );
  MUX2X1 U1164 ( .B(n1190), .A(n1191), .S(n879), .Y(n1168) );
  MUX2X1 U1165 ( .B(A[63]), .A(A[62]), .S(n876), .Y(n1191) );
  MUX2X1 U1166 ( .B(A[61]), .A(A[60]), .S(n875), .Y(n1190) );
  MUX2X1 U1167 ( .B(n1165), .A(n1166), .S(n883), .Y(n1035) );
  MUX2X1 U1168 ( .B(n1188), .A(n1181), .S(n879), .Y(n1166) );
  MUX2X1 U1169 ( .B(A[51]), .A(A[50]), .S(n876), .Y(n1181) );
  MUX2X1 U1170 ( .B(A[49]), .A(A[48]), .S(n875), .Y(n1188) );
  MUX2X1 U1171 ( .B(n1182), .A(n1183), .S(n879), .Y(n1165) );
  MUX2X1 U1172 ( .B(A[55]), .A(A[54]), .S(n875), .Y(n1183) );
  MUX2X1 U1173 ( .B(A[53]), .A(A[52]), .S(n876), .Y(n1182) );
  MUX2X1 U1174 ( .B(n1104), .A(n1210), .S(n889), .Y(n1209) );
  MUX2X1 U1175 ( .B(n905), .A(n1211), .S(n885), .Y(n1210) );
  MUX2X1 U1176 ( .B(n951), .A(n1212), .S(n883), .Y(n1211) );
  MUX2X1 U1177 ( .B(n1213), .A(n1004), .S(n879), .Y(n1212) );
  MUX2X1 U1178 ( .B(A[3]), .A(A[2]), .S(n876), .Y(n1004) );
  MUX2X1 U1179 ( .B(A[1]), .A(A[0]), .S(n875), .Y(n1213) );
  MUX2X1 U1180 ( .B(n1005), .A(n1006), .S(n879), .Y(n951) );
  MUX2X1 U1181 ( .B(A[7]), .A(A[6]), .S(n876), .Y(n1006) );
  MUX2X1 U1182 ( .B(A[5]), .A(A[4]), .S(n875), .Y(n1005) );
  MUX2X1 U1183 ( .B(n1171), .A(n950), .S(n883), .Y(n905) );
  MUX2X1 U1184 ( .B(n1007), .A(n1193), .S(n879), .Y(n950) );
  MUX2X1 U1185 ( .B(A[11]), .A(A[10]), .S(n876), .Y(n1193) );
  MUX2X1 U1186 ( .B(A[9]), .A(A[8]), .S(n875), .Y(n1007) );
  MUX2X1 U1187 ( .B(n1194), .A(n1195), .S(n879), .Y(n1171) );
  MUX2X1 U1188 ( .B(A[15]), .A(A[14]), .S(n876), .Y(n1195) );
  MUX2X1 U1189 ( .B(A[13]), .A(A[12]), .S(n875), .Y(n1194) );
  MUX2X1 U1190 ( .B(n904), .A(n1032), .S(n887), .Y(n1104) );
  MUX2X1 U1191 ( .B(n1177), .A(n1172), .S(n883), .Y(n1032) );
  MUX2X1 U1192 ( .B(n1200), .A(n1205), .S(n879), .Y(n1172) );
  MUX2X1 U1193 ( .B(A[27]), .A(A[26]), .S(n876), .Y(n1205) );
  MUX2X1 U1194 ( .B(A[25]), .A(A[24]), .S(n875), .Y(n1200) );
  MUX2X1 U1195 ( .B(n1206), .A(n1207), .S(n879), .Y(n1177) );
  MUX2X1 U1196 ( .B(A[31]), .A(A[30]), .S(n876), .Y(n1207) );
  MUX2X1 U1197 ( .B(A[29]), .A(A[28]), .S(n876), .Y(n1206) );
  MUX2X1 U1198 ( .B(n1173), .A(n1170), .S(n884), .Y(n904) );
  MUX2X1 U1199 ( .B(n1196), .A(n1197), .S(n879), .Y(n1170) );
  MUX2X1 U1200 ( .B(A[19]), .A(A[18]), .S(n876), .Y(n1197) );
  MUX2X1 U1201 ( .B(A[17]), .A(A[16]), .S(n875), .Y(n1196) );
  MUX2X1 U1202 ( .B(n1198), .A(n1199), .S(n879), .Y(n1173) );
  MUX2X1 U1203 ( .B(A[23]), .A(A[22]), .S(n876), .Y(n1199) );
  MUX2X1 U1204 ( .B(A[21]), .A(A[20]), .S(n876), .Y(n1198) );
endmodule


module alu_DW_rightsh_46 ( A, DATA_TC, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC;
  wire   n542, n541, n540, n539, n538, n537, n536, n535, n534, n533, n532,
         n357, n359, n360, n361, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n380, n381,
         n383, n384, n385, n386, n387, n388, n391, n392, n393, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531;

  OR2X1 U308 ( .A(n359), .B(n369), .Y(n485) );
  AND2X1 U309 ( .A(n360), .B(n373), .Y(n462) );
  AND2X1 U310 ( .A(n365), .B(n373), .Y(n460) );
  AND2X1 U311 ( .A(n364), .B(n378), .Y(B[24]) );
  OR2X1 U312 ( .A(n377), .B(n366), .Y(n532) );
  INVX1 U313 ( .A(n532), .Y(B[31]) );
  OR2X1 U314 ( .A(n357), .B(n377), .Y(n534) );
  INVX1 U315 ( .A(n534), .Y(B[29]) );
  OR2X1 U316 ( .A(n377), .B(n426), .Y(n542) );
  INVX1 U317 ( .A(n542), .Y(B[20]) );
  OR2X1 U318 ( .A(n377), .B(n420), .Y(n541) );
  INVX1 U319 ( .A(n541), .Y(B[21]) );
  OR2X1 U320 ( .A(n377), .B(n414), .Y(n540) );
  INVX1 U321 ( .A(n540), .Y(B[22]) );
  OR2X1 U322 ( .A(n377), .B(n408), .Y(n539) );
  INVX1 U323 ( .A(n539), .Y(B[23]) );
  OR2X1 U324 ( .A(n399), .B(n377), .Y(n538) );
  INVX1 U325 ( .A(n538), .Y(B[25]) );
  OR2X1 U326 ( .A(n457), .B(n377), .Y(n537) );
  INVX1 U327 ( .A(n537), .Y(B[26]) );
  OR2X1 U328 ( .A(n377), .B(n361), .Y(n533) );
  INVX1 U329 ( .A(n533), .Y(B[30]) );
  AND2X1 U330 ( .A(n464), .B(n375), .Y(n454) );
  INVX1 U331 ( .A(n454), .Y(n357) );
  OR2X1 U332 ( .A(n363), .B(n377), .Y(n535) );
  INVX1 U333 ( .A(n535), .Y(B[28]) );
  AND2X1 U334 ( .A(A[31]), .B(n368), .Y(n497) );
  INVX1 U335 ( .A(n497), .Y(n359) );
  OR2X1 U336 ( .A(n515), .B(n369), .Y(n491) );
  INVX1 U337 ( .A(n491), .Y(n360) );
  AND2X1 U338 ( .A(n462), .B(n375), .Y(n443) );
  INVX1 U339 ( .A(n443), .Y(n361) );
  OR2X1 U340 ( .A(n456), .B(n377), .Y(n536) );
  INVX1 U341 ( .A(n536), .Y(B[27]) );
  AND2X1 U342 ( .A(n466), .B(n375), .Y(n455) );
  INVX1 U343 ( .A(n455), .Y(n363) );
  OR2X1 U344 ( .A(n459), .B(n374), .Y(n405) );
  INVX1 U345 ( .A(n405), .Y(n364) );
  INVX1 U346 ( .A(n485), .Y(n365) );
  AND2X1 U347 ( .A(n460), .B(n375), .Y(n442) );
  INVX1 U348 ( .A(n442), .Y(n366) );
  INVX1 U349 ( .A(n461), .Y(n385) );
  INVX1 U350 ( .A(n463), .Y(n397) );
  INVX1 U351 ( .A(n465), .Y(n387) );
  INVX1 U352 ( .A(n467), .Y(n392) );
  INVX1 U353 ( .A(n514), .Y(n388) );
  INVX1 U354 ( .A(n518), .Y(n393) );
  INVX1 U355 ( .A(n400), .Y(n380) );
  INVX1 U356 ( .A(n409), .Y(n383) );
  INVX1 U357 ( .A(n427), .Y(n398) );
  INVX1 U358 ( .A(n421), .Y(n381) );
  INVX1 U359 ( .A(n403), .Y(B[8]) );
  INVX1 U360 ( .A(n486), .Y(n384) );
  INVX1 U361 ( .A(n492), .Y(n395) );
  INVX1 U362 ( .A(n499), .Y(n386) );
  INVX1 U363 ( .A(n509), .Y(n391) );
  INVX1 U364 ( .A(SH[1]), .Y(n370) );
  INVX1 U365 ( .A(n432), .Y(B[3]) );
  INVX1 U366 ( .A(n444), .Y(B[2]) );
  INVX1 U367 ( .A(n373), .Y(n371) );
  INVX1 U368 ( .A(n373), .Y(n372) );
  INVX1 U369 ( .A(n375), .Y(n374) );
  INVX1 U370 ( .A(n378), .Y(n376) );
  INVX1 U371 ( .A(n378), .Y(n377) );
  INVX1 U372 ( .A(n527), .Y(B[0]) );
  INVX1 U373 ( .A(n370), .Y(n369) );
  INVX1 U374 ( .A(n368), .Y(n367) );
  INVX1 U375 ( .A(SH[0]), .Y(n368) );
  INVX1 U376 ( .A(SH[2]), .Y(n373) );
  INVX1 U377 ( .A(SH[4]), .Y(n378) );
  INVX1 U378 ( .A(SH[3]), .Y(n375) );
  INVX1 U379 ( .A(n415), .Y(n396) );
  INVX1 U380 ( .A(n468), .Y(B[1]) );
  MUX2X1 U381 ( .B(n380), .A(n399), .S(n376), .Y(B[9]) );
  MUX2X1 U382 ( .B(n401), .A(n402), .S(n374), .Y(n400) );
  MUX2X1 U383 ( .B(n404), .A(n364), .S(n376), .Y(n403) );
  MUX2X1 U384 ( .B(n406), .A(n407), .S(SH[3]), .Y(n404) );
  MUX2X1 U385 ( .B(n383), .A(n408), .S(n377), .Y(B[7]) );
  MUX2X1 U386 ( .B(n410), .A(n411), .S(SH[3]), .Y(n409) );
  MUX2X1 U387 ( .B(n412), .A(n413), .S(n371), .Y(n410) );
  MUX2X1 U388 ( .B(n396), .A(n414), .S(n377), .Y(B[6]) );
  MUX2X1 U389 ( .B(n416), .A(n417), .S(SH[3]), .Y(n415) );
  MUX2X1 U390 ( .B(n418), .A(n419), .S(n371), .Y(n416) );
  MUX2X1 U391 ( .B(n381), .A(n420), .S(n376), .Y(B[5]) );
  MUX2X1 U392 ( .B(n422), .A(n423), .S(SH[3]), .Y(n421) );
  MUX2X1 U393 ( .B(n424), .A(n425), .S(n371), .Y(n422) );
  MUX2X1 U394 ( .B(n398), .A(n426), .S(n377), .Y(B[4]) );
  MUX2X1 U395 ( .B(n428), .A(n429), .S(SH[3]), .Y(n427) );
  MUX2X1 U396 ( .B(n430), .A(n431), .S(n371), .Y(n428) );
  MUX2X1 U397 ( .B(n433), .A(n434), .S(n377), .Y(n432) );
  MUX2X1 U398 ( .B(n435), .A(n436), .S(SH[3]), .Y(n433) );
  MUX2X1 U399 ( .B(n437), .A(n412), .S(n371), .Y(n435) );
  MUX2X1 U400 ( .B(n438), .A(n439), .S(SH[1]), .Y(n412) );
  MUX2X1 U401 ( .B(n440), .A(n441), .S(SH[1]), .Y(n437) );
  MUX2X1 U402 ( .B(n445), .A(n446), .S(n376), .Y(n444) );
  MUX2X1 U403 ( .B(n447), .A(n448), .S(SH[3]), .Y(n445) );
  MUX2X1 U404 ( .B(n449), .A(n418), .S(n371), .Y(n447) );
  MUX2X1 U405 ( .B(n450), .A(n451), .S(n369), .Y(n418) );
  MUX2X1 U406 ( .B(n452), .A(n453), .S(n369), .Y(n449) );
  OR2X1 U407 ( .A(n458), .B(SH[3]), .Y(n399) );
  MUX2X1 U408 ( .B(n385), .A(n460), .S(SH[3]), .Y(n408) );
  MUX2X1 U409 ( .B(n397), .A(n462), .S(SH[3]), .Y(n414) );
  MUX2X1 U410 ( .B(n387), .A(n464), .S(SH[3]), .Y(n420) );
  MUX2X1 U411 ( .B(n392), .A(n466), .S(n374), .Y(n426) );
  MUX2X1 U412 ( .B(n469), .A(n470), .S(n376), .Y(n468) );
  MUX2X1 U413 ( .B(n471), .A(n401), .S(n374), .Y(n469) );
  MUX2X1 U414 ( .B(n472), .A(n425), .S(n373), .Y(n401) );
  MUX2X1 U415 ( .B(n439), .A(n473), .S(n369), .Y(n425) );
  MUX2X1 U416 ( .B(A[9]), .A(A[10]), .S(n367), .Y(n439) );
  MUX2X1 U417 ( .B(n474), .A(n424), .S(n371), .Y(n471) );
  MUX2X1 U418 ( .B(n441), .A(n438), .S(n369), .Y(n424) );
  MUX2X1 U419 ( .B(A[7]), .A(A[8]), .S(n367), .Y(n438) );
  MUX2X1 U420 ( .B(A[5]), .A(A[6]), .S(n367), .Y(n441) );
  MUX2X1 U421 ( .B(n475), .A(n440), .S(n369), .Y(n474) );
  MUX2X1 U422 ( .B(A[3]), .A(A[4]), .S(n367), .Y(n440) );
  MUX2X1 U423 ( .B(A[1]), .A(A[2]), .S(n367), .Y(n475) );
  AND2X1 U424 ( .A(n434), .B(n378), .Y(B[19]) );
  MUX2X1 U425 ( .B(n476), .A(n477), .S(n374), .Y(n434) );
  AND2X1 U426 ( .A(n446), .B(n378), .Y(B[18]) );
  MUX2X1 U427 ( .B(n478), .A(n479), .S(n374), .Y(n446) );
  AND2X1 U428 ( .A(n378), .B(n470), .Y(B[17]) );
  MUX2X1 U429 ( .B(n402), .A(n458), .S(n374), .Y(n470) );
  MUX2X1 U430 ( .B(n480), .A(n481), .S(n371), .Y(n458) );
  MUX2X1 U431 ( .B(n482), .A(n483), .S(n371), .Y(n402) );
  AND2X1 U432 ( .A(n484), .B(n378), .Y(B[16]) );
  MUX2X1 U433 ( .B(n384), .A(n366), .S(n376), .Y(B[15]) );
  MUX2X1 U434 ( .B(n411), .A(n461), .S(n374), .Y(n486) );
  MUX2X1 U435 ( .B(n487), .A(n488), .S(n371), .Y(n461) );
  MUX2X1 U436 ( .B(n489), .A(n490), .S(n371), .Y(n411) );
  MUX2X1 U437 ( .B(n395), .A(n361), .S(n376), .Y(B[14]) );
  MUX2X1 U438 ( .B(n417), .A(n463), .S(n374), .Y(n492) );
  MUX2X1 U439 ( .B(n493), .A(n494), .S(n371), .Y(n463) );
  MUX2X1 U440 ( .B(n495), .A(n496), .S(n372), .Y(n417) );
  MUX2X1 U441 ( .B(n386), .A(n357), .S(n376), .Y(B[13]) );
  AND2X1 U442 ( .A(n481), .B(n373), .Y(n464) );
  MUX2X1 U443 ( .B(n359), .A(n498), .S(n370), .Y(n481) );
  MUX2X1 U444 ( .B(n423), .A(n465), .S(n374), .Y(n499) );
  MUX2X1 U445 ( .B(n483), .A(n480), .S(n372), .Y(n465) );
  MUX2X1 U446 ( .B(n500), .A(n501), .S(n370), .Y(n480) );
  MUX2X1 U447 ( .B(n502), .A(n503), .S(n370), .Y(n483) );
  MUX2X1 U448 ( .B(n472), .A(n482), .S(n372), .Y(n423) );
  MUX2X1 U449 ( .B(n504), .A(n505), .S(n370), .Y(n482) );
  MUX2X1 U450 ( .B(n506), .A(n507), .S(n370), .Y(n472) );
  MUX2X1 U451 ( .B(n391), .A(n363), .S(n376), .Y(B[12]) );
  AND2X1 U452 ( .A(n508), .B(n373), .Y(n466) );
  MUX2X1 U453 ( .B(n429), .A(n467), .S(n374), .Y(n509) );
  MUX2X1 U454 ( .B(n510), .A(n511), .S(n372), .Y(n467) );
  MUX2X1 U455 ( .B(n512), .A(n513), .S(n372), .Y(n429) );
  MUX2X1 U456 ( .B(n388), .A(n456), .S(n376), .Y(B[11]) );
  OR2X1 U457 ( .A(n477), .B(SH[3]), .Y(n456) );
  MUX2X1 U458 ( .B(n488), .A(n365), .S(n372), .Y(n477) );
  MUX2X1 U459 ( .B(n498), .A(n500), .S(n370), .Y(n488) );
  MUX2X1 U460 ( .B(A[27]), .A(A[28]), .S(n367), .Y(n500) );
  MUX2X1 U461 ( .B(A[29]), .A(A[30]), .S(n367), .Y(n498) );
  MUX2X1 U462 ( .B(n436), .A(n476), .S(n374), .Y(n514) );
  MUX2X1 U463 ( .B(n490), .A(n487), .S(n372), .Y(n476) );
  MUX2X1 U464 ( .B(n501), .A(n502), .S(n370), .Y(n487) );
  MUX2X1 U465 ( .B(A[23]), .A(A[24]), .S(n367), .Y(n502) );
  MUX2X1 U466 ( .B(A[25]), .A(A[26]), .S(n367), .Y(n501) );
  MUX2X1 U467 ( .B(n503), .A(n504), .S(n370), .Y(n490) );
  MUX2X1 U468 ( .B(A[19]), .A(A[20]), .S(n367), .Y(n504) );
  MUX2X1 U469 ( .B(A[21]), .A(A[22]), .S(n367), .Y(n503) );
  MUX2X1 U470 ( .B(n413), .A(n489), .S(n372), .Y(n436) );
  MUX2X1 U471 ( .B(n505), .A(n506), .S(n370), .Y(n489) );
  MUX2X1 U472 ( .B(A[15]), .A(A[16]), .S(n367), .Y(n506) );
  MUX2X1 U473 ( .B(A[17]), .A(A[18]), .S(SH[0]), .Y(n505) );
  MUX2X1 U474 ( .B(n473), .A(n507), .S(n369), .Y(n413) );
  MUX2X1 U475 ( .B(A[13]), .A(A[14]), .S(SH[0]), .Y(n507) );
  MUX2X1 U476 ( .B(A[11]), .A(A[12]), .S(SH[0]), .Y(n473) );
  MUX2X1 U477 ( .B(n393), .A(n457), .S(n376), .Y(B[10]) );
  OR2X1 U478 ( .A(n479), .B(n374), .Y(n457) );
  MUX2X1 U479 ( .B(n494), .A(n360), .S(n372), .Y(n479) );
  MUX2X1 U480 ( .B(n516), .A(n517), .S(n370), .Y(n494) );
  MUX2X1 U481 ( .B(n448), .A(n478), .S(n374), .Y(n518) );
  MUX2X1 U482 ( .B(n496), .A(n493), .S(n372), .Y(n478) );
  MUX2X1 U483 ( .B(n519), .A(n520), .S(n370), .Y(n493) );
  MUX2X1 U484 ( .B(n521), .A(n522), .S(n370), .Y(n496) );
  MUX2X1 U485 ( .B(n419), .A(n495), .S(n372), .Y(n448) );
  MUX2X1 U486 ( .B(n523), .A(n524), .S(n370), .Y(n495) );
  MUX2X1 U487 ( .B(n525), .A(n526), .S(n369), .Y(n419) );
  MUX2X1 U488 ( .B(n528), .A(n484), .S(n376), .Y(n527) );
  MUX2X1 U489 ( .B(n459), .A(n407), .S(n375), .Y(n484) );
  MUX2X1 U490 ( .B(n513), .A(n510), .S(n372), .Y(n407) );
  MUX2X1 U491 ( .B(n520), .A(n521), .S(n370), .Y(n510) );
  MUX2X1 U492 ( .B(A[20]), .A(A[21]), .S(SH[0]), .Y(n521) );
  MUX2X1 U493 ( .B(A[22]), .A(A[23]), .S(SH[0]), .Y(n520) );
  MUX2X1 U494 ( .B(n522), .A(n523), .S(n370), .Y(n513) );
  MUX2X1 U495 ( .B(A[16]), .A(A[17]), .S(SH[0]), .Y(n523) );
  MUX2X1 U496 ( .B(A[18]), .A(A[19]), .S(SH[0]), .Y(n522) );
  MUX2X1 U497 ( .B(n511), .A(n508), .S(n372), .Y(n459) );
  MUX2X1 U498 ( .B(n515), .A(n516), .S(n370), .Y(n508) );
  MUX2X1 U499 ( .B(A[28]), .A(A[29]), .S(SH[0]), .Y(n516) );
  MUX2X1 U500 ( .B(A[30]), .A(A[31]), .S(SH[0]), .Y(n515) );
  MUX2X1 U501 ( .B(n517), .A(n519), .S(n370), .Y(n511) );
  MUX2X1 U502 ( .B(A[24]), .A(A[25]), .S(SH[0]), .Y(n519) );
  MUX2X1 U503 ( .B(A[26]), .A(A[27]), .S(SH[0]), .Y(n517) );
  MUX2X1 U504 ( .B(n529), .A(n406), .S(SH[3]), .Y(n528) );
  MUX2X1 U505 ( .B(n431), .A(n512), .S(n372), .Y(n406) );
  MUX2X1 U506 ( .B(n524), .A(n526), .S(n370), .Y(n512) );
  MUX2X1 U507 ( .B(A[12]), .A(A[13]), .S(SH[0]), .Y(n526) );
  MUX2X1 U508 ( .B(A[14]), .A(A[15]), .S(n367), .Y(n524) );
  MUX2X1 U509 ( .B(n451), .A(n525), .S(n369), .Y(n431) );
  MUX2X1 U510 ( .B(A[10]), .A(A[11]), .S(n367), .Y(n525) );
  MUX2X1 U511 ( .B(A[8]), .A(A[9]), .S(n367), .Y(n451) );
  MUX2X1 U512 ( .B(n530), .A(n430), .S(n372), .Y(n529) );
  MUX2X1 U513 ( .B(n453), .A(n450), .S(n369), .Y(n430) );
  MUX2X1 U514 ( .B(A[6]), .A(A[7]), .S(SH[0]), .Y(n450) );
  MUX2X1 U515 ( .B(A[4]), .A(A[5]), .S(SH[0]), .Y(n453) );
  MUX2X1 U516 ( .B(n531), .A(n452), .S(SH[1]), .Y(n530) );
  MUX2X1 U517 ( .B(A[2]), .A(A[3]), .S(SH[0]), .Y(n452) );
  MUX2X1 U518 ( .B(A[0]), .A(A[1]), .S(SH[0]), .Y(n531) );
endmodule


module alu_DW_rightsh_47 ( A, DATA_TC, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC;
  wire   n546, n545, n544, n543, n542, n541, n540, n539, n538, n537, n536,
         n357, n359, n360, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n384, n385, n387, n388, n389, n390, n391, n392, n395,
         n396, n397, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535;

  AND2X1 U308 ( .A(n359), .B(n376), .Y(n464) );
  AND2X1 U309 ( .A(n364), .B(n382), .Y(B[24]) );
  OR2X1 U310 ( .A(n357), .B(n381), .Y(n538) );
  INVX1 U311 ( .A(n538), .Y(B[29]) );
  OR2X1 U312 ( .A(n381), .B(n366), .Y(n536) );
  INVX1 U313 ( .A(n536), .Y(B[31]) );
  OR2X1 U314 ( .A(n381), .B(n360), .Y(n537) );
  INVX1 U315 ( .A(n537), .Y(B[30]) );
  OR2X1 U316 ( .A(n381), .B(n430), .Y(n546) );
  INVX1 U317 ( .A(n546), .Y(B[20]) );
  OR2X1 U318 ( .A(n381), .B(n424), .Y(n545) );
  INVX1 U319 ( .A(n545), .Y(B[21]) );
  OR2X1 U320 ( .A(n381), .B(n418), .Y(n544) );
  INVX1 U321 ( .A(n544), .Y(B[22]) );
  OR2X1 U322 ( .A(n381), .B(n412), .Y(n543) );
  INVX1 U323 ( .A(n543), .Y(B[23]) );
  OR2X1 U324 ( .A(n403), .B(n381), .Y(n542) );
  INVX1 U325 ( .A(n542), .Y(B[25]) );
  OR2X1 U326 ( .A(n461), .B(n381), .Y(n541) );
  INVX1 U327 ( .A(n541), .Y(B[26]) );
  AND2X1 U328 ( .A(n468), .B(n379), .Y(n458) );
  INVX1 U329 ( .A(n458), .Y(n357) );
  OR2X1 U330 ( .A(n363), .B(n381), .Y(n539) );
  INVX1 U331 ( .A(n539), .Y(B[28]) );
  OR2X1 U332 ( .A(n362), .B(n372), .Y(n489) );
  INVX1 U333 ( .A(n489), .Y(n359) );
  AND2X1 U334 ( .A(n466), .B(n379), .Y(n447) );
  INVX1 U335 ( .A(n447), .Y(n360) );
  AND2X1 U336 ( .A(n365), .B(n376), .Y(n466) );
  OR2X1 U337 ( .A(n460), .B(n381), .Y(n540) );
  INVX1 U338 ( .A(n540), .Y(B[27]) );
  AND2X1 U339 ( .A(A[31]), .B(n369), .Y(n501) );
  INVX1 U340 ( .A(n501), .Y(n362) );
  AND2X1 U341 ( .A(n470), .B(n379), .Y(n459) );
  INVX1 U342 ( .A(n459), .Y(n363) );
  OR2X1 U343 ( .A(n463), .B(n377), .Y(n409) );
  INVX1 U344 ( .A(n409), .Y(n364) );
  OR2X1 U345 ( .A(n519), .B(n372), .Y(n495) );
  INVX1 U346 ( .A(n495), .Y(n365) );
  AND2X1 U347 ( .A(n464), .B(n379), .Y(n446) );
  INVX1 U348 ( .A(n446), .Y(n366) );
  INVX1 U349 ( .A(n465), .Y(n389) );
  INVX1 U350 ( .A(n467), .Y(n401) );
  INVX1 U351 ( .A(n469), .Y(n391) );
  INVX1 U352 ( .A(n471), .Y(n396) );
  INVX1 U353 ( .A(n379), .Y(n378) );
  INVX1 U354 ( .A(n379), .Y(n377) );
  INVX1 U355 ( .A(n496), .Y(n399) );
  INVX1 U356 ( .A(n490), .Y(n388) );
  INVX1 U357 ( .A(n503), .Y(n390) );
  INVX1 U358 ( .A(n518), .Y(n392) );
  INVX1 U359 ( .A(n522), .Y(n397) );
  INVX1 U360 ( .A(n404), .Y(n384) );
  INVX1 U361 ( .A(n413), .Y(n387) );
  INVX1 U362 ( .A(n425), .Y(n385) );
  INVX1 U363 ( .A(n431), .Y(n402) );
  INVX1 U364 ( .A(n513), .Y(n395) );
  INVX1 U365 ( .A(n376), .Y(n374) );
  INVX1 U366 ( .A(n376), .Y(n375) );
  INVX1 U367 ( .A(n436), .Y(B[3]) );
  INVX1 U368 ( .A(n407), .Y(B[8]) );
  INVX1 U369 ( .A(SH[3]), .Y(n379) );
  INVX1 U370 ( .A(n382), .Y(n380) );
  INVX1 U371 ( .A(n382), .Y(n381) );
  INVX1 U372 ( .A(n373), .Y(n371) );
  INVX1 U373 ( .A(n373), .Y(n370) );
  INVX1 U374 ( .A(SH[2]), .Y(n376) );
  INVX1 U375 ( .A(n531), .Y(B[0]) );
  INVX1 U376 ( .A(n373), .Y(n372) );
  INVX1 U377 ( .A(SH[1]), .Y(n373) );
  INVX1 U378 ( .A(SH[4]), .Y(n382) );
  INVX1 U379 ( .A(n419), .Y(n400) );
  INVX1 U380 ( .A(n369), .Y(n368) );
  INVX1 U381 ( .A(SH[0]), .Y(n369) );
  INVX1 U382 ( .A(n369), .Y(n367) );
  INVX1 U383 ( .A(n448), .Y(B[2]) );
  INVX1 U384 ( .A(n472), .Y(B[1]) );
  MUX2X1 U385 ( .B(n384), .A(n403), .S(n380), .Y(B[9]) );
  MUX2X1 U386 ( .B(n405), .A(n406), .S(n377), .Y(n404) );
  MUX2X1 U387 ( .B(n408), .A(n364), .S(n380), .Y(n407) );
  MUX2X1 U388 ( .B(n410), .A(n411), .S(n378), .Y(n408) );
  MUX2X1 U389 ( .B(n387), .A(n412), .S(n381), .Y(B[7]) );
  MUX2X1 U390 ( .B(n414), .A(n415), .S(n378), .Y(n413) );
  MUX2X1 U391 ( .B(n416), .A(n417), .S(n374), .Y(n414) );
  MUX2X1 U392 ( .B(n400), .A(n418), .S(n381), .Y(B[6]) );
  MUX2X1 U393 ( .B(n420), .A(n421), .S(n378), .Y(n419) );
  MUX2X1 U394 ( .B(n422), .A(n423), .S(n374), .Y(n420) );
  MUX2X1 U395 ( .B(n385), .A(n424), .S(n380), .Y(B[5]) );
  MUX2X1 U396 ( .B(n426), .A(n427), .S(n378), .Y(n425) );
  MUX2X1 U397 ( .B(n428), .A(n429), .S(n374), .Y(n426) );
  MUX2X1 U398 ( .B(n402), .A(n430), .S(n381), .Y(B[4]) );
  MUX2X1 U399 ( .B(n432), .A(n433), .S(n378), .Y(n431) );
  MUX2X1 U400 ( .B(n434), .A(n435), .S(n374), .Y(n432) );
  MUX2X1 U401 ( .B(n437), .A(n438), .S(n381), .Y(n436) );
  MUX2X1 U402 ( .B(n439), .A(n440), .S(n378), .Y(n437) );
  MUX2X1 U403 ( .B(n441), .A(n416), .S(n374), .Y(n439) );
  MUX2X1 U404 ( .B(n442), .A(n443), .S(n370), .Y(n416) );
  MUX2X1 U405 ( .B(n444), .A(n445), .S(n370), .Y(n441) );
  MUX2X1 U406 ( .B(n449), .A(n450), .S(n380), .Y(n448) );
  MUX2X1 U407 ( .B(n451), .A(n452), .S(n378), .Y(n449) );
  MUX2X1 U408 ( .B(n453), .A(n422), .S(n374), .Y(n451) );
  MUX2X1 U409 ( .B(n454), .A(n455), .S(n371), .Y(n422) );
  MUX2X1 U410 ( .B(n456), .A(n457), .S(n371), .Y(n453) );
  OR2X1 U411 ( .A(n462), .B(n378), .Y(n403) );
  MUX2X1 U412 ( .B(n389), .A(n464), .S(n378), .Y(n412) );
  MUX2X1 U413 ( .B(n401), .A(n466), .S(n378), .Y(n418) );
  MUX2X1 U414 ( .B(n391), .A(n468), .S(n378), .Y(n424) );
  MUX2X1 U415 ( .B(n396), .A(n470), .S(n377), .Y(n430) );
  MUX2X1 U416 ( .B(n473), .A(n474), .S(n380), .Y(n472) );
  MUX2X1 U417 ( .B(n475), .A(n405), .S(n377), .Y(n473) );
  MUX2X1 U418 ( .B(n476), .A(n429), .S(n376), .Y(n405) );
  MUX2X1 U419 ( .B(n443), .A(n477), .S(n371), .Y(n429) );
  MUX2X1 U420 ( .B(A[9]), .A(A[10]), .S(n367), .Y(n443) );
  MUX2X1 U421 ( .B(n478), .A(n428), .S(n374), .Y(n475) );
  MUX2X1 U422 ( .B(n445), .A(n442), .S(n371), .Y(n428) );
  MUX2X1 U423 ( .B(A[7]), .A(A[8]), .S(n367), .Y(n442) );
  MUX2X1 U424 ( .B(A[5]), .A(A[6]), .S(n367), .Y(n445) );
  MUX2X1 U425 ( .B(n479), .A(n444), .S(n371), .Y(n478) );
  MUX2X1 U426 ( .B(A[3]), .A(A[4]), .S(n367), .Y(n444) );
  MUX2X1 U427 ( .B(A[1]), .A(A[2]), .S(n367), .Y(n479) );
  AND2X1 U428 ( .A(n438), .B(n382), .Y(B[19]) );
  MUX2X1 U429 ( .B(n480), .A(n481), .S(n377), .Y(n438) );
  AND2X1 U430 ( .A(n450), .B(n382), .Y(B[18]) );
  MUX2X1 U431 ( .B(n482), .A(n483), .S(n377), .Y(n450) );
  AND2X1 U432 ( .A(n382), .B(n474), .Y(B[17]) );
  MUX2X1 U433 ( .B(n406), .A(n462), .S(n377), .Y(n474) );
  MUX2X1 U434 ( .B(n484), .A(n485), .S(n374), .Y(n462) );
  MUX2X1 U435 ( .B(n486), .A(n487), .S(n374), .Y(n406) );
  AND2X1 U436 ( .A(n488), .B(n382), .Y(B[16]) );
  MUX2X1 U437 ( .B(n388), .A(n366), .S(n380), .Y(B[15]) );
  MUX2X1 U438 ( .B(n415), .A(n465), .S(n377), .Y(n490) );
  MUX2X1 U439 ( .B(n491), .A(n492), .S(n374), .Y(n465) );
  MUX2X1 U440 ( .B(n493), .A(n494), .S(n374), .Y(n415) );
  MUX2X1 U441 ( .B(n399), .A(n360), .S(n380), .Y(B[14]) );
  MUX2X1 U442 ( .B(n421), .A(n467), .S(n377), .Y(n496) );
  MUX2X1 U443 ( .B(n497), .A(n498), .S(n374), .Y(n467) );
  MUX2X1 U444 ( .B(n499), .A(n500), .S(n375), .Y(n421) );
  MUX2X1 U445 ( .B(n390), .A(n357), .S(n380), .Y(B[13]) );
  AND2X1 U446 ( .A(n485), .B(n376), .Y(n468) );
  MUX2X1 U447 ( .B(n362), .A(n502), .S(n373), .Y(n485) );
  MUX2X1 U448 ( .B(n427), .A(n469), .S(n377), .Y(n503) );
  MUX2X1 U449 ( .B(n487), .A(n484), .S(n375), .Y(n469) );
  MUX2X1 U450 ( .B(n504), .A(n505), .S(n373), .Y(n484) );
  MUX2X1 U451 ( .B(n506), .A(n507), .S(n373), .Y(n487) );
  MUX2X1 U452 ( .B(n476), .A(n486), .S(n375), .Y(n427) );
  MUX2X1 U453 ( .B(n508), .A(n509), .S(n373), .Y(n486) );
  MUX2X1 U454 ( .B(n510), .A(n511), .S(n373), .Y(n476) );
  MUX2X1 U455 ( .B(n395), .A(n363), .S(n380), .Y(B[12]) );
  AND2X1 U456 ( .A(n512), .B(n376), .Y(n470) );
  MUX2X1 U457 ( .B(n433), .A(n471), .S(n377), .Y(n513) );
  MUX2X1 U458 ( .B(n514), .A(n515), .S(n375), .Y(n471) );
  MUX2X1 U459 ( .B(n516), .A(n517), .S(n375), .Y(n433) );
  MUX2X1 U460 ( .B(n392), .A(n460), .S(n380), .Y(B[11]) );
  OR2X1 U461 ( .A(n481), .B(n378), .Y(n460) );
  MUX2X1 U462 ( .B(n492), .A(n359), .S(n375), .Y(n481) );
  MUX2X1 U463 ( .B(n502), .A(n504), .S(n373), .Y(n492) );
  MUX2X1 U464 ( .B(A[27]), .A(A[28]), .S(n367), .Y(n504) );
  MUX2X1 U465 ( .B(A[29]), .A(A[30]), .S(n367), .Y(n502) );
  MUX2X1 U466 ( .B(n440), .A(n480), .S(n377), .Y(n518) );
  MUX2X1 U467 ( .B(n494), .A(n491), .S(n375), .Y(n480) );
  MUX2X1 U468 ( .B(n505), .A(n506), .S(n373), .Y(n491) );
  MUX2X1 U469 ( .B(A[23]), .A(A[24]), .S(n367), .Y(n506) );
  MUX2X1 U470 ( .B(A[25]), .A(A[26]), .S(n367), .Y(n505) );
  MUX2X1 U471 ( .B(n507), .A(n508), .S(n373), .Y(n494) );
  MUX2X1 U472 ( .B(A[19]), .A(A[20]), .S(n367), .Y(n508) );
  MUX2X1 U473 ( .B(A[21]), .A(A[22]), .S(n367), .Y(n507) );
  MUX2X1 U474 ( .B(n417), .A(n493), .S(n375), .Y(n440) );
  MUX2X1 U475 ( .B(n509), .A(n510), .S(n373), .Y(n493) );
  MUX2X1 U476 ( .B(A[15]), .A(A[16]), .S(n367), .Y(n510) );
  MUX2X1 U477 ( .B(A[17]), .A(A[18]), .S(n368), .Y(n509) );
  MUX2X1 U478 ( .B(n477), .A(n511), .S(n371), .Y(n417) );
  MUX2X1 U479 ( .B(A[13]), .A(A[14]), .S(n368), .Y(n511) );
  MUX2X1 U480 ( .B(A[11]), .A(A[12]), .S(n368), .Y(n477) );
  MUX2X1 U481 ( .B(n397), .A(n461), .S(n380), .Y(B[10]) );
  OR2X1 U482 ( .A(n483), .B(n378), .Y(n461) );
  MUX2X1 U483 ( .B(n498), .A(n365), .S(n375), .Y(n483) );
  MUX2X1 U484 ( .B(n520), .A(n521), .S(n373), .Y(n498) );
  MUX2X1 U485 ( .B(n452), .A(n482), .S(n377), .Y(n522) );
  MUX2X1 U486 ( .B(n500), .A(n497), .S(n375), .Y(n482) );
  MUX2X1 U487 ( .B(n523), .A(n524), .S(n373), .Y(n497) );
  MUX2X1 U488 ( .B(n525), .A(n526), .S(n373), .Y(n500) );
  MUX2X1 U489 ( .B(n423), .A(n499), .S(n375), .Y(n452) );
  MUX2X1 U490 ( .B(n527), .A(n528), .S(n373), .Y(n499) );
  MUX2X1 U491 ( .B(n529), .A(n530), .S(n371), .Y(n423) );
  MUX2X1 U492 ( .B(n532), .A(n488), .S(n380), .Y(n531) );
  MUX2X1 U493 ( .B(n463), .A(n411), .S(n379), .Y(n488) );
  MUX2X1 U494 ( .B(n517), .A(n514), .S(n375), .Y(n411) );
  MUX2X1 U495 ( .B(n524), .A(n525), .S(n373), .Y(n514) );
  MUX2X1 U496 ( .B(A[20]), .A(A[21]), .S(n368), .Y(n525) );
  MUX2X1 U497 ( .B(A[22]), .A(A[23]), .S(n368), .Y(n524) );
  MUX2X1 U498 ( .B(n526), .A(n527), .S(n373), .Y(n517) );
  MUX2X1 U499 ( .B(A[16]), .A(A[17]), .S(n368), .Y(n527) );
  MUX2X1 U500 ( .B(A[18]), .A(A[19]), .S(n368), .Y(n526) );
  MUX2X1 U501 ( .B(n515), .A(n512), .S(n375), .Y(n463) );
  MUX2X1 U502 ( .B(n519), .A(n520), .S(n373), .Y(n512) );
  MUX2X1 U503 ( .B(A[28]), .A(A[29]), .S(n368), .Y(n520) );
  MUX2X1 U504 ( .B(A[30]), .A(A[31]), .S(n368), .Y(n519) );
  MUX2X1 U505 ( .B(n521), .A(n523), .S(n373), .Y(n515) );
  MUX2X1 U506 ( .B(A[24]), .A(A[25]), .S(n368), .Y(n523) );
  MUX2X1 U507 ( .B(A[26]), .A(A[27]), .S(n368), .Y(n521) );
  MUX2X1 U508 ( .B(n533), .A(n410), .S(n378), .Y(n532) );
  MUX2X1 U509 ( .B(n435), .A(n516), .S(n374), .Y(n410) );
  MUX2X1 U510 ( .B(n528), .A(n530), .S(n373), .Y(n516) );
  MUX2X1 U511 ( .B(A[12]), .A(A[13]), .S(n368), .Y(n530) );
  MUX2X1 U512 ( .B(A[14]), .A(A[15]), .S(n367), .Y(n528) );
  MUX2X1 U513 ( .B(n455), .A(n529), .S(n372), .Y(n435) );
  MUX2X1 U514 ( .B(A[10]), .A(A[11]), .S(n367), .Y(n529) );
  MUX2X1 U515 ( .B(A[8]), .A(A[9]), .S(n368), .Y(n455) );
  MUX2X1 U516 ( .B(n534), .A(n434), .S(n375), .Y(n533) );
  MUX2X1 U517 ( .B(n457), .A(n454), .S(n371), .Y(n434) );
  MUX2X1 U518 ( .B(A[6]), .A(A[7]), .S(n368), .Y(n454) );
  MUX2X1 U519 ( .B(A[4]), .A(A[5]), .S(n367), .Y(n457) );
  MUX2X1 U520 ( .B(n535), .A(n456), .S(n370), .Y(n534) );
  MUX2X1 U521 ( .B(A[2]), .A(A[3]), .S(n367), .Y(n456) );
  MUX2X1 U522 ( .B(A[0]), .A(A[1]), .S(n367), .Y(n535) );
endmodule


module alu_DW_leftsh_0 ( A, SH, B );
  input [63:0] A;
  input [4:0] SH;
  output [63:0] B;
  wire   n1141, n1140, n1139, n1138, n1137, n1136, n1135, n1134, n1133, n1132,
         n1131, n1130, n749, n751, n752, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n790, n792, n793, n795, n796, n797, n799,
         n800, n802, n804, n806, n808, n810, n812, n814, n816, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129;

  OR2X1 U668 ( .A(n752), .B(n765), .Y(n1123) );
  AND2X1 U669 ( .A(n756), .B(n774), .Y(n1069) );
  OR2X1 U670 ( .A(n749), .B(n784), .Y(n1139) );
  INVX1 U671 ( .A(n1139), .Y(B[2]) );
  OR2X1 U672 ( .A(n941), .B(n783), .Y(n1137) );
  INVX1 U673 ( .A(n1137), .Y(B[4]) );
  OR2X1 U674 ( .A(n754), .B(n784), .Y(n1138) );
  INVX1 U675 ( .A(n1138), .Y(B[3]) );
  OR2X1 U676 ( .A(n783), .B(n1056), .Y(n1130) );
  INVX1 U677 ( .A(n1130), .Y(B[11]) );
  OR2X1 U678 ( .A(n876), .B(n784), .Y(n1136) );
  INVX1 U679 ( .A(n1136), .Y(B[5]) );
  OR2X1 U680 ( .A(n783), .B(n1060), .Y(n1131) );
  INVX1 U681 ( .A(n1131), .Y(B[10]) );
  OR2X1 U682 ( .A(n840), .B(n783), .Y(n1134) );
  INVX1 U683 ( .A(n1134), .Y(B[7]) );
  OR2X1 U684 ( .A(n841), .B(n783), .Y(n1135) );
  INVX1 U685 ( .A(n1135), .Y(B[6]) );
  OR2X1 U686 ( .A(n751), .B(n784), .Y(n1140) );
  INVX1 U687 ( .A(n1140), .Y(B[1]) );
  OR2X1 U688 ( .A(n784), .B(n839), .Y(n1133) );
  INVX1 U689 ( .A(n1133), .Y(B[8]) );
  AND2X1 U690 ( .A(n1095), .B(n780), .Y(n1045) );
  INVX1 U691 ( .A(n1045), .Y(n749) );
  OR2X1 U692 ( .A(n784), .B(n757), .Y(n1141) );
  INVX1 U693 ( .A(n1141), .Y(B[0]) );
  AND2X1 U694 ( .A(n1064), .B(n780), .Y(n1090) );
  INVX1 U695 ( .A(n1090), .Y(n751) );
  AND2X1 U696 ( .A(n755), .B(n774), .Y(n1064) );
  AND2X1 U697 ( .A(A[0]), .B(n762), .Y(n1129) );
  INVX1 U698 ( .A(n1129), .Y(n752) );
  OR2X1 U699 ( .A(n784), .B(n838), .Y(n1132) );
  INVX1 U700 ( .A(n1132), .Y(B[9]) );
  AND2X1 U701 ( .A(n1091), .B(n780), .Y(n994) );
  INVX1 U702 ( .A(n994), .Y(n754) );
  OR2X1 U703 ( .A(n1117), .B(n763), .Y(n1099) );
  INVX1 U704 ( .A(n1099), .Y(n755) );
  INVX1 U705 ( .A(n1123), .Y(n756) );
  AND2X1 U706 ( .A(n1069), .B(n780), .Y(n1104) );
  INVX1 U707 ( .A(n1104), .Y(n757) );
  INVX1 U708 ( .A(n1096), .Y(n796) );
  INVX1 U709 ( .A(n1065), .Y(n795) );
  INVX1 U710 ( .A(n1070), .Y(n792) );
  INVX1 U711 ( .A(n774), .Y(n773) );
  INVX1 U712 ( .A(n774), .Y(n772) );
  INVX1 U713 ( .A(n764), .Y(n768) );
  INVX1 U714 ( .A(n764), .Y(n769) );
  INVX1 U715 ( .A(n1092), .Y(n799) );
  INVX1 U716 ( .A(n1001), .Y(n806) );
  INVX1 U717 ( .A(n884), .Y(B[58]) );
  INVX1 U718 ( .A(n860), .Y(B[61]) );
  INVX1 U719 ( .A(n935), .Y(B[50]) );
  INVX1 U720 ( .A(n1035), .Y(B[31]) );
  INVX1 U721 ( .A(n954), .Y(B[47]) );
  INVX1 U722 ( .A(n942), .Y(B[49]) );
  INVX1 U723 ( .A(n1025), .Y(B[33]) );
  INVX1 U724 ( .A(n979), .Y(B[42]) );
  INVX1 U725 ( .A(n964), .Y(B[45]) );
  INVX1 U726 ( .A(n1016), .Y(n800) );
  INVX1 U727 ( .A(n1031), .Y(n790) );
  INVX1 U728 ( .A(n974), .Y(B[43]) );
  INVX1 U729 ( .A(n1015), .Y(B[35]) );
  INVX1 U730 ( .A(n959), .Y(B[46]) );
  INVX1 U731 ( .A(n923), .Y(B[52]) );
  INVX1 U732 ( .A(n989), .Y(B[40]) );
  INVX1 U733 ( .A(n995), .Y(B[39]) );
  INVX1 U734 ( .A(n905), .Y(B[55]) );
  INVX1 U735 ( .A(n990), .Y(n810) );
  INVX1 U736 ( .A(n996), .Y(n808) );
  INVX1 U737 ( .A(n877), .Y(B[59]) );
  INVX1 U738 ( .A(n929), .Y(B[51]) );
  INVX1 U739 ( .A(n1010), .Y(B[36]) );
  INVX1 U740 ( .A(n975), .Y(n816) );
  INVX1 U741 ( .A(n868), .Y(B[60]) );
  INVX1 U742 ( .A(n911), .Y(B[54]) );
  INVX1 U743 ( .A(n948), .Y(B[48]) );
  INVX1 U744 ( .A(n1046), .Y(B[29]) );
  INVX1 U745 ( .A(n1051), .Y(B[28]) );
  INVX1 U746 ( .A(n980), .Y(n814) );
  INVX1 U747 ( .A(n985), .Y(n812) );
  INVX1 U748 ( .A(n1021), .Y(n797) );
  INVX1 U749 ( .A(n780), .Y(n777) );
  INVX1 U750 ( .A(n780), .Y(n778) );
  INVX1 U751 ( .A(n780), .Y(n776) );
  INVX1 U752 ( .A(n780), .Y(n775) );
  INVX1 U753 ( .A(n1020), .Y(B[34]) );
  INVX1 U754 ( .A(n780), .Y(n779) );
  INVX1 U755 ( .A(n1011), .Y(n802) );
  INVX1 U756 ( .A(n766), .Y(n765) );
  INVX1 U757 ( .A(n766), .Y(n764) );
  INVX1 U758 ( .A(n762), .Y(n761) );
  INVX1 U759 ( .A(n762), .Y(n758) );
  INVX1 U760 ( .A(n762), .Y(n759) );
  INVX1 U761 ( .A(n762), .Y(n760) );
  INVX1 U762 ( .A(SH[0]), .Y(n762) );
  INVX1 U763 ( .A(n763), .Y(n771) );
  INVX1 U764 ( .A(n763), .Y(n770) );
  INVX1 U765 ( .A(n1026), .Y(n793) );
  INVX1 U766 ( .A(n1006), .Y(n804) );
  INVX1 U767 ( .A(SH[2]), .Y(n774) );
  INVX1 U768 ( .A(n898), .Y(B[56]) );
  INVX1 U769 ( .A(n851), .Y(B[62]) );
  INVX1 U770 ( .A(n1040), .Y(B[30]) );
  INVX1 U771 ( .A(n1030), .Y(B[32]) );
  INVX1 U772 ( .A(n1000), .Y(B[38]) );
  INVX1 U773 ( .A(n891), .Y(B[57]) );
  INVX1 U774 ( .A(n917), .Y(B[53]) );
  INVX1 U775 ( .A(n984), .Y(B[41]) );
  INVX1 U776 ( .A(n1005), .Y(B[37]) );
  INVX1 U777 ( .A(n969), .Y(B[44]) );
  INVX1 U778 ( .A(n842), .Y(B[63]) );
  INVX1 U779 ( .A(SH[3]), .Y(n780) );
  INVX1 U780 ( .A(SH[1]), .Y(n766) );
  INVX1 U781 ( .A(n785), .Y(n784) );
  INVX1 U782 ( .A(n785), .Y(n781) );
  INVX1 U783 ( .A(n785), .Y(n782) );
  INVX1 U784 ( .A(n785), .Y(n783) );
  INVX1 U785 ( .A(n767), .Y(n763) );
  INVX1 U786 ( .A(SH[1]), .Y(n767) );
  INVX1 U787 ( .A(SH[4]), .Y(n785) );
  MUX2X1 U788 ( .B(n843), .A(n844), .S(n785), .Y(n842) );
  MUX2X1 U789 ( .B(n845), .A(n846), .S(n775), .Y(n844) );
  MUX2X1 U790 ( .B(n847), .A(n848), .S(n772), .Y(n845) );
  MUX2X1 U791 ( .B(n849), .A(n850), .S(n764), .Y(n847) );
  MUX2X1 U792 ( .B(A[63]), .A(A[62]), .S(n758), .Y(n849) );
  MUX2X1 U793 ( .B(n852), .A(n853), .S(n781), .Y(n851) );
  MUX2X1 U794 ( .B(n854), .A(n855), .S(n779), .Y(n852) );
  MUX2X1 U795 ( .B(n856), .A(n857), .S(n772), .Y(n854) );
  MUX2X1 U796 ( .B(n858), .A(n859), .S(n764), .Y(n856) );
  MUX2X1 U797 ( .B(A[62]), .A(A[61]), .S(n758), .Y(n858) );
  MUX2X1 U798 ( .B(n861), .A(n862), .S(n781), .Y(n860) );
  MUX2X1 U799 ( .B(n863), .A(n864), .S(n779), .Y(n861) );
  MUX2X1 U800 ( .B(n865), .A(n866), .S(n772), .Y(n863) );
  MUX2X1 U801 ( .B(n850), .A(n867), .S(n764), .Y(n865) );
  MUX2X1 U802 ( .B(A[61]), .A(A[60]), .S(n758), .Y(n850) );
  MUX2X1 U803 ( .B(n869), .A(n870), .S(n781), .Y(n868) );
  MUX2X1 U804 ( .B(n871), .A(n872), .S(n779), .Y(n869) );
  MUX2X1 U805 ( .B(n873), .A(n874), .S(n772), .Y(n871) );
  MUX2X1 U806 ( .B(n859), .A(n875), .S(n765), .Y(n873) );
  MUX2X1 U807 ( .B(A[60]), .A(A[59]), .S(n758), .Y(n859) );
  MUX2X1 U808 ( .B(n878), .A(n879), .S(n781), .Y(n877) );
  MUX2X1 U809 ( .B(n880), .A(n881), .S(n779), .Y(n878) );
  MUX2X1 U810 ( .B(n848), .A(n882), .S(n772), .Y(n880) );
  MUX2X1 U811 ( .B(n867), .A(n883), .S(n765), .Y(n848) );
  MUX2X1 U812 ( .B(A[59]), .A(A[58]), .S(n758), .Y(n867) );
  MUX2X1 U813 ( .B(n885), .A(n886), .S(n781), .Y(n884) );
  MUX2X1 U814 ( .B(n887), .A(n888), .S(n779), .Y(n885) );
  MUX2X1 U815 ( .B(n857), .A(n889), .S(n772), .Y(n887) );
  MUX2X1 U816 ( .B(n875), .A(n890), .S(n765), .Y(n857) );
  MUX2X1 U817 ( .B(A[58]), .A(A[57]), .S(n758), .Y(n875) );
  MUX2X1 U818 ( .B(n892), .A(n893), .S(n781), .Y(n891) );
  MUX2X1 U819 ( .B(n894), .A(n895), .S(n779), .Y(n892) );
  MUX2X1 U820 ( .B(n866), .A(n896), .S(n772), .Y(n894) );
  MUX2X1 U821 ( .B(n883), .A(n897), .S(n765), .Y(n866) );
  MUX2X1 U822 ( .B(A[57]), .A(A[56]), .S(n758), .Y(n883) );
  MUX2X1 U823 ( .B(n899), .A(n900), .S(n781), .Y(n898) );
  MUX2X1 U824 ( .B(n901), .A(n902), .S(n779), .Y(n899) );
  MUX2X1 U825 ( .B(n874), .A(n903), .S(n772), .Y(n901) );
  MUX2X1 U826 ( .B(n890), .A(n904), .S(n765), .Y(n874) );
  MUX2X1 U827 ( .B(A[56]), .A(A[55]), .S(n758), .Y(n890) );
  MUX2X1 U828 ( .B(n906), .A(n907), .S(n782), .Y(n905) );
  MUX2X1 U829 ( .B(n846), .A(n908), .S(n779), .Y(n906) );
  MUX2X1 U830 ( .B(n882), .A(n909), .S(n772), .Y(n846) );
  MUX2X1 U831 ( .B(n897), .A(n910), .S(n765), .Y(n882) );
  MUX2X1 U832 ( .B(A[55]), .A(A[54]), .S(n758), .Y(n897) );
  MUX2X1 U833 ( .B(n912), .A(n913), .S(n782), .Y(n911) );
  MUX2X1 U834 ( .B(n855), .A(n914), .S(n778), .Y(n912) );
  MUX2X1 U835 ( .B(n915), .A(n889), .S(n774), .Y(n855) );
  MUX2X1 U836 ( .B(n904), .A(n916), .S(n765), .Y(n889) );
  MUX2X1 U837 ( .B(A[54]), .A(A[53]), .S(n758), .Y(n904) );
  MUX2X1 U838 ( .B(n918), .A(n919), .S(n782), .Y(n917) );
  MUX2X1 U839 ( .B(n864), .A(n920), .S(n778), .Y(n918) );
  MUX2X1 U840 ( .B(n896), .A(n921), .S(n772), .Y(n864) );
  MUX2X1 U841 ( .B(n910), .A(n922), .S(n765), .Y(n896) );
  MUX2X1 U842 ( .B(A[53]), .A(A[52]), .S(n758), .Y(n910) );
  MUX2X1 U843 ( .B(n924), .A(n925), .S(n782), .Y(n923) );
  MUX2X1 U844 ( .B(n872), .A(n926), .S(n778), .Y(n924) );
  MUX2X1 U845 ( .B(n903), .A(n927), .S(n772), .Y(n872) );
  MUX2X1 U846 ( .B(n916), .A(n928), .S(n765), .Y(n903) );
  MUX2X1 U847 ( .B(A[52]), .A(A[51]), .S(n758), .Y(n916) );
  MUX2X1 U848 ( .B(n930), .A(n931), .S(n782), .Y(n929) );
  MUX2X1 U849 ( .B(n881), .A(n932), .S(n778), .Y(n930) );
  MUX2X1 U850 ( .B(n909), .A(n933), .S(n772), .Y(n881) );
  MUX2X1 U851 ( .B(n934), .A(n922), .S(n768), .Y(n909) );
  MUX2X1 U852 ( .B(A[51]), .A(A[50]), .S(n759), .Y(n922) );
  MUX2X1 U853 ( .B(n936), .A(n937), .S(n782), .Y(n935) );
  MUX2X1 U854 ( .B(n888), .A(n938), .S(n778), .Y(n936) );
  MUX2X1 U855 ( .B(n915), .A(n939), .S(SH[2]), .Y(n888) );
  MUX2X1 U856 ( .B(n940), .A(n928), .S(n768), .Y(n915) );
  MUX2X1 U857 ( .B(A[50]), .A(A[49]), .S(n759), .Y(n928) );
  MUX2X1 U858 ( .B(n943), .A(n944), .S(n782), .Y(n942) );
  MUX2X1 U859 ( .B(n895), .A(n945), .S(n778), .Y(n943) );
  MUX2X1 U860 ( .B(n921), .A(n946), .S(SH[2]), .Y(n895) );
  MUX2X1 U861 ( .B(n947), .A(n934), .S(n768), .Y(n921) );
  MUX2X1 U862 ( .B(A[49]), .A(A[48]), .S(n759), .Y(n934) );
  MUX2X1 U863 ( .B(n949), .A(n950), .S(n782), .Y(n948) );
  MUX2X1 U864 ( .B(n902), .A(n951), .S(n778), .Y(n949) );
  MUX2X1 U865 ( .B(n927), .A(n952), .S(SH[2]), .Y(n902) );
  MUX2X1 U866 ( .B(n953), .A(n940), .S(n768), .Y(n927) );
  MUX2X1 U867 ( .B(A[48]), .A(A[47]), .S(n759), .Y(n940) );
  MUX2X1 U868 ( .B(n843), .A(n955), .S(n782), .Y(n954) );
  MUX2X1 U869 ( .B(n908), .A(n956), .S(n778), .Y(n843) );
  MUX2X1 U870 ( .B(n933), .A(n957), .S(n773), .Y(n908) );
  MUX2X1 U871 ( .B(n958), .A(n947), .S(n768), .Y(n933) );
  MUX2X1 U872 ( .B(A[47]), .A(A[46]), .S(n759), .Y(n947) );
  MUX2X1 U873 ( .B(n853), .A(n960), .S(n782), .Y(n959) );
  MUX2X1 U874 ( .B(n914), .A(n961), .S(n778), .Y(n853) );
  MUX2X1 U875 ( .B(n939), .A(n962), .S(SH[2]), .Y(n914) );
  MUX2X1 U876 ( .B(n963), .A(n953), .S(n768), .Y(n939) );
  MUX2X1 U877 ( .B(A[46]), .A(A[45]), .S(n759), .Y(n953) );
  MUX2X1 U878 ( .B(n862), .A(n965), .S(n782), .Y(n964) );
  MUX2X1 U879 ( .B(n920), .A(n966), .S(n778), .Y(n862) );
  MUX2X1 U880 ( .B(n946), .A(n967), .S(SH[2]), .Y(n920) );
  MUX2X1 U881 ( .B(n968), .A(n958), .S(n768), .Y(n946) );
  MUX2X1 U882 ( .B(A[45]), .A(A[44]), .S(n759), .Y(n958) );
  MUX2X1 U883 ( .B(n870), .A(n970), .S(n783), .Y(n969) );
  MUX2X1 U884 ( .B(n926), .A(n971), .S(n778), .Y(n870) );
  MUX2X1 U885 ( .B(n952), .A(n972), .S(SH[2]), .Y(n926) );
  MUX2X1 U886 ( .B(n973), .A(n963), .S(n768), .Y(n952) );
  MUX2X1 U887 ( .B(A[44]), .A(A[43]), .S(n759), .Y(n963) );
  MUX2X1 U888 ( .B(n879), .A(n975), .S(n783), .Y(n974) );
  MUX2X1 U889 ( .B(n932), .A(n976), .S(n778), .Y(n879) );
  MUX2X1 U890 ( .B(n957), .A(n977), .S(SH[2]), .Y(n932) );
  MUX2X1 U891 ( .B(n978), .A(n968), .S(n768), .Y(n957) );
  MUX2X1 U892 ( .B(A[43]), .A(A[42]), .S(n759), .Y(n968) );
  MUX2X1 U893 ( .B(n886), .A(n980), .S(n783), .Y(n979) );
  MUX2X1 U894 ( .B(n938), .A(n981), .S(n777), .Y(n886) );
  MUX2X1 U895 ( .B(n962), .A(n982), .S(SH[2]), .Y(n938) );
  MUX2X1 U896 ( .B(n983), .A(n973), .S(n768), .Y(n962) );
  MUX2X1 U897 ( .B(A[42]), .A(A[41]), .S(n759), .Y(n973) );
  MUX2X1 U898 ( .B(n893), .A(n985), .S(n783), .Y(n984) );
  MUX2X1 U899 ( .B(n945), .A(n986), .S(n777), .Y(n893) );
  MUX2X1 U900 ( .B(n967), .A(n987), .S(SH[2]), .Y(n945) );
  MUX2X1 U901 ( .B(n988), .A(n978), .S(n768), .Y(n967) );
  MUX2X1 U902 ( .B(A[41]), .A(A[40]), .S(n759), .Y(n978) );
  MUX2X1 U903 ( .B(n900), .A(n990), .S(n783), .Y(n989) );
  MUX2X1 U904 ( .B(n951), .A(n991), .S(n777), .Y(n900) );
  MUX2X1 U905 ( .B(n972), .A(n992), .S(SH[2]), .Y(n951) );
  MUX2X1 U906 ( .B(n993), .A(n983), .S(n768), .Y(n972) );
  MUX2X1 U907 ( .B(A[40]), .A(A[39]), .S(n759), .Y(n983) );
  MUX2X1 U908 ( .B(n907), .A(n996), .S(n783), .Y(n995) );
  MUX2X1 U909 ( .B(n956), .A(n997), .S(n777), .Y(n907) );
  MUX2X1 U910 ( .B(n977), .A(n998), .S(SH[2]), .Y(n956) );
  MUX2X1 U911 ( .B(n999), .A(n988), .S(n769), .Y(n977) );
  MUX2X1 U912 ( .B(A[39]), .A(A[38]), .S(n760), .Y(n988) );
  MUX2X1 U913 ( .B(n913), .A(n1001), .S(n783), .Y(n1000) );
  MUX2X1 U914 ( .B(n961), .A(n1002), .S(n777), .Y(n913) );
  MUX2X1 U915 ( .B(n982), .A(n1003), .S(n773), .Y(n961) );
  MUX2X1 U916 ( .B(n1004), .A(n993), .S(n769), .Y(n982) );
  MUX2X1 U917 ( .B(A[38]), .A(A[37]), .S(n760), .Y(n993) );
  MUX2X1 U918 ( .B(n919), .A(n1006), .S(n783), .Y(n1005) );
  MUX2X1 U919 ( .B(n966), .A(n1007), .S(n777), .Y(n919) );
  MUX2X1 U920 ( .B(n987), .A(n1008), .S(n773), .Y(n966) );
  MUX2X1 U921 ( .B(n1009), .A(n999), .S(n769), .Y(n987) );
  MUX2X1 U922 ( .B(A[37]), .A(A[36]), .S(n760), .Y(n999) );
  MUX2X1 U923 ( .B(n925), .A(n1011), .S(n783), .Y(n1010) );
  MUX2X1 U924 ( .B(n971), .A(n1012), .S(n777), .Y(n925) );
  MUX2X1 U925 ( .B(n992), .A(n1013), .S(n773), .Y(n971) );
  MUX2X1 U926 ( .B(n1014), .A(n1004), .S(n769), .Y(n992) );
  MUX2X1 U927 ( .B(A[36]), .A(A[35]), .S(n760), .Y(n1004) );
  MUX2X1 U928 ( .B(n931), .A(n1016), .S(n783), .Y(n1015) );
  MUX2X1 U929 ( .B(n976), .A(n1017), .S(n777), .Y(n931) );
  MUX2X1 U930 ( .B(n998), .A(n1018), .S(n773), .Y(n976) );
  MUX2X1 U931 ( .B(n1019), .A(n1009), .S(n769), .Y(n998) );
  MUX2X1 U932 ( .B(A[35]), .A(A[34]), .S(n760), .Y(n1009) );
  MUX2X1 U933 ( .B(n937), .A(n1021), .S(n783), .Y(n1020) );
  MUX2X1 U934 ( .B(n981), .A(n1022), .S(n777), .Y(n937) );
  MUX2X1 U935 ( .B(n1003), .A(n1023), .S(n773), .Y(n981) );
  MUX2X1 U936 ( .B(n1024), .A(n1014), .S(n769), .Y(n1003) );
  MUX2X1 U937 ( .B(A[34]), .A(A[33]), .S(n760), .Y(n1014) );
  MUX2X1 U938 ( .B(n944), .A(n1026), .S(n784), .Y(n1025) );
  MUX2X1 U939 ( .B(n986), .A(n1027), .S(n777), .Y(n944) );
  MUX2X1 U940 ( .B(n1008), .A(n1028), .S(n773), .Y(n986) );
  MUX2X1 U941 ( .B(n1029), .A(n1019), .S(n769), .Y(n1008) );
  MUX2X1 U942 ( .B(A[33]), .A(A[32]), .S(n760), .Y(n1019) );
  MUX2X1 U943 ( .B(n950), .A(n1031), .S(n784), .Y(n1030) );
  MUX2X1 U944 ( .B(n991), .A(n1032), .S(n777), .Y(n950) );
  MUX2X1 U945 ( .B(n1013), .A(n1033), .S(n773), .Y(n991) );
  MUX2X1 U946 ( .B(n1034), .A(n1024), .S(n769), .Y(n1013) );
  MUX2X1 U947 ( .B(A[32]), .A(A[31]), .S(n760), .Y(n1024) );
  MUX2X1 U948 ( .B(n955), .A(n1036), .S(n784), .Y(n1035) );
  MUX2X1 U949 ( .B(n997), .A(n1037), .S(n776), .Y(n955) );
  MUX2X1 U950 ( .B(n1018), .A(n1038), .S(n773), .Y(n997) );
  MUX2X1 U951 ( .B(n1039), .A(n1029), .S(n769), .Y(n1018) );
  MUX2X1 U952 ( .B(A[31]), .A(A[30]), .S(n760), .Y(n1029) );
  MUX2X1 U953 ( .B(n960), .A(n1041), .S(n784), .Y(n1040) );
  MUX2X1 U954 ( .B(n1002), .A(n1042), .S(n776), .Y(n960) );
  MUX2X1 U955 ( .B(n1023), .A(n1043), .S(n773), .Y(n1002) );
  MUX2X1 U956 ( .B(n1044), .A(n1034), .S(n769), .Y(n1023) );
  MUX2X1 U957 ( .B(A[30]), .A(A[29]), .S(n760), .Y(n1034) );
  MUX2X1 U958 ( .B(n965), .A(n1047), .S(n784), .Y(n1046) );
  MUX2X1 U959 ( .B(n1007), .A(n1048), .S(n776), .Y(n965) );
  MUX2X1 U960 ( .B(n1028), .A(n1049), .S(n773), .Y(n1007) );
  MUX2X1 U961 ( .B(n1050), .A(n1039), .S(n769), .Y(n1028) );
  MUX2X1 U962 ( .B(A[29]), .A(A[28]), .S(n760), .Y(n1039) );
  MUX2X1 U963 ( .B(n970), .A(n1052), .S(n784), .Y(n1051) );
  MUX2X1 U964 ( .B(n1012), .A(n1053), .S(n776), .Y(n970) );
  MUX2X1 U965 ( .B(n1033), .A(n1054), .S(n773), .Y(n1012) );
  MUX2X1 U966 ( .B(n1055), .A(n1044), .S(n769), .Y(n1033) );
  MUX2X1 U967 ( .B(A[28]), .A(A[27]), .S(n760), .Y(n1044) );
  MUX2X1 U968 ( .B(n816), .A(n1056), .S(n784), .Y(B[27]) );
  MUX2X1 U969 ( .B(n1017), .A(n1057), .S(n776), .Y(n975) );
  MUX2X1 U970 ( .B(n1038), .A(n1058), .S(n773), .Y(n1017) );
  MUX2X1 U971 ( .B(n1059), .A(n1050), .S(n770), .Y(n1038) );
  MUX2X1 U972 ( .B(A[27]), .A(A[26]), .S(n758), .Y(n1050) );
  MUX2X1 U973 ( .B(n814), .A(n1060), .S(n784), .Y(B[26]) );
  MUX2X1 U974 ( .B(n1022), .A(n1061), .S(n776), .Y(n980) );
  MUX2X1 U975 ( .B(n1043), .A(n1062), .S(SH[2]), .Y(n1022) );
  MUX2X1 U976 ( .B(n1063), .A(n1055), .S(n770), .Y(n1043) );
  MUX2X1 U977 ( .B(A[26]), .A(A[25]), .S(SH[0]), .Y(n1055) );
  MUX2X1 U978 ( .B(n812), .A(n838), .S(n784), .Y(B[25]) );
  MUX2X1 U979 ( .B(n795), .A(n1064), .S(n776), .Y(n838) );
  MUX2X1 U980 ( .B(n1027), .A(n1066), .S(n776), .Y(n985) );
  MUX2X1 U981 ( .B(n1049), .A(n1067), .S(SH[2]), .Y(n1027) );
  MUX2X1 U982 ( .B(n1068), .A(n1059), .S(n770), .Y(n1049) );
  MUX2X1 U983 ( .B(A[25]), .A(A[24]), .S(SH[0]), .Y(n1059) );
  MUX2X1 U984 ( .B(n810), .A(n839), .S(n784), .Y(B[24]) );
  MUX2X1 U985 ( .B(n792), .A(n1069), .S(n776), .Y(n839) );
  MUX2X1 U986 ( .B(n1032), .A(n1071), .S(n776), .Y(n990) );
  MUX2X1 U987 ( .B(n1054), .A(n1072), .S(SH[2]), .Y(n1032) );
  MUX2X1 U988 ( .B(n1073), .A(n1063), .S(n770), .Y(n1054) );
  MUX2X1 U989 ( .B(A[24]), .A(A[23]), .S(SH[0]), .Y(n1063) );
  MUX2X1 U990 ( .B(n808), .A(n840), .S(n784), .Y(B[23]) );
  OR2X1 U991 ( .A(n1074), .B(n779), .Y(n840) );
  MUX2X1 U992 ( .B(n1037), .A(n1075), .S(n776), .Y(n996) );
  MUX2X1 U993 ( .B(n1058), .A(n1076), .S(SH[2]), .Y(n1037) );
  MUX2X1 U994 ( .B(n1077), .A(n1068), .S(n770), .Y(n1058) );
  MUX2X1 U995 ( .B(A[23]), .A(A[22]), .S(n759), .Y(n1068) );
  MUX2X1 U996 ( .B(n806), .A(n841), .S(n783), .Y(B[22]) );
  OR2X1 U997 ( .A(n1078), .B(n779), .Y(n841) );
  MUX2X1 U998 ( .B(n1042), .A(n1079), .S(n776), .Y(n1001) );
  MUX2X1 U999 ( .B(n1062), .A(n1080), .S(SH[2]), .Y(n1042) );
  MUX2X1 U1000 ( .B(n1081), .A(n1073), .S(n770), .Y(n1062) );
  MUX2X1 U1001 ( .B(A[22]), .A(A[21]), .S(SH[0]), .Y(n1073) );
  MUX2X1 U1002 ( .B(n804), .A(n876), .S(n782), .Y(B[21]) );
  OR2X1 U1003 ( .A(n1082), .B(n779), .Y(n876) );
  MUX2X1 U1004 ( .B(n1048), .A(n1083), .S(n775), .Y(n1006) );
  MUX2X1 U1005 ( .B(n1067), .A(n1084), .S(SH[2]), .Y(n1048) );
  MUX2X1 U1006 ( .B(n1085), .A(n1077), .S(n770), .Y(n1067) );
  MUX2X1 U1007 ( .B(A[21]), .A(A[20]), .S(n760), .Y(n1077) );
  MUX2X1 U1008 ( .B(n802), .A(n941), .S(n781), .Y(B[20]) );
  OR2X1 U1009 ( .A(n1086), .B(n779), .Y(n941) );
  MUX2X1 U1010 ( .B(n1053), .A(n1087), .S(n775), .Y(n1011) );
  MUX2X1 U1011 ( .B(n1072), .A(n1088), .S(SH[2]), .Y(n1053) );
  MUX2X1 U1012 ( .B(n1089), .A(n1081), .S(n770), .Y(n1072) );
  MUX2X1 U1013 ( .B(A[20]), .A(A[19]), .S(SH[0]), .Y(n1081) );
  MUX2X1 U1014 ( .B(n800), .A(n754), .S(n781), .Y(B[19]) );
  MUX2X1 U1015 ( .B(n1057), .A(n1092), .S(n775), .Y(n1016) );
  MUX2X1 U1016 ( .B(n1076), .A(n1093), .S(SH[2]), .Y(n1057) );
  MUX2X1 U1017 ( .B(n1094), .A(n1085), .S(n770), .Y(n1076) );
  MUX2X1 U1018 ( .B(A[19]), .A(A[18]), .S(n761), .Y(n1085) );
  MUX2X1 U1019 ( .B(n797), .A(n749), .S(n781), .Y(B[18]) );
  MUX2X1 U1020 ( .B(n1061), .A(n1096), .S(n775), .Y(n1021) );
  MUX2X1 U1021 ( .B(n1080), .A(n1097), .S(SH[2]), .Y(n1061) );
  MUX2X1 U1022 ( .B(n1098), .A(n1089), .S(n770), .Y(n1080) );
  MUX2X1 U1023 ( .B(A[18]), .A(A[17]), .S(SH[0]), .Y(n1089) );
  MUX2X1 U1024 ( .B(n793), .A(n751), .S(n781), .Y(B[17]) );
  MUX2X1 U1025 ( .B(n1066), .A(n1065), .S(n775), .Y(n1026) );
  MUX2X1 U1026 ( .B(n1100), .A(n1101), .S(SH[2]), .Y(n1065) );
  MUX2X1 U1027 ( .B(n1084), .A(n1102), .S(SH[2]), .Y(n1066) );
  MUX2X1 U1028 ( .B(n1103), .A(n1094), .S(n770), .Y(n1084) );
  MUX2X1 U1029 ( .B(A[17]), .A(A[16]), .S(SH[0]), .Y(n1094) );
  MUX2X1 U1030 ( .B(n790), .A(n757), .S(n781), .Y(B[16]) );
  MUX2X1 U1031 ( .B(n1071), .A(n1070), .S(n775), .Y(n1031) );
  MUX2X1 U1032 ( .B(n1105), .A(n1106), .S(SH[2]), .Y(n1070) );
  MUX2X1 U1033 ( .B(n1088), .A(n1107), .S(SH[2]), .Y(n1071) );
  MUX2X1 U1034 ( .B(n1108), .A(n1098), .S(n770), .Y(n1088) );
  MUX2X1 U1035 ( .B(A[16]), .A(A[15]), .S(SH[0]), .Y(n1098) );
  AND2X1 U1036 ( .A(n785), .B(n1036), .Y(B[15]) );
  MUX2X1 U1037 ( .B(n1075), .A(n1074), .S(n775), .Y(n1036) );
  MUX2X1 U1038 ( .B(n1109), .A(n1110), .S(n772), .Y(n1074) );
  MUX2X1 U1039 ( .B(n1093), .A(n1111), .S(n772), .Y(n1075) );
  MUX2X1 U1040 ( .B(n1112), .A(n1103), .S(n771), .Y(n1093) );
  MUX2X1 U1041 ( .B(A[15]), .A(A[14]), .S(n761), .Y(n1103) );
  AND2X1 U1042 ( .A(n785), .B(n1041), .Y(B[14]) );
  MUX2X1 U1043 ( .B(n1079), .A(n1078), .S(n775), .Y(n1041) );
  MUX2X1 U1044 ( .B(n1113), .A(n1114), .S(n772), .Y(n1078) );
  MUX2X1 U1045 ( .B(n1097), .A(n1115), .S(n772), .Y(n1079) );
  MUX2X1 U1046 ( .B(n1116), .A(n1108), .S(n771), .Y(n1097) );
  MUX2X1 U1047 ( .B(A[14]), .A(A[13]), .S(n761), .Y(n1108) );
  AND2X1 U1048 ( .A(n1047), .B(n785), .Y(B[13]) );
  MUX2X1 U1049 ( .B(n1083), .A(n1082), .S(n775), .Y(n1047) );
  MUX2X1 U1050 ( .B(n1101), .A(n755), .S(n772), .Y(n1082) );
  MUX2X1 U1051 ( .B(n1118), .A(n1119), .S(n771), .Y(n1101) );
  MUX2X1 U1052 ( .B(n1102), .A(n1100), .S(n773), .Y(n1083) );
  MUX2X1 U1053 ( .B(n1120), .A(n1121), .S(n771), .Y(n1100) );
  MUX2X1 U1054 ( .B(n1122), .A(n1112), .S(n771), .Y(n1102) );
  MUX2X1 U1055 ( .B(A[13]), .A(A[12]), .S(n761), .Y(n1112) );
  AND2X1 U1056 ( .A(n1052), .B(n785), .Y(B[12]) );
  MUX2X1 U1057 ( .B(n1087), .A(n1086), .S(n775), .Y(n1052) );
  MUX2X1 U1058 ( .B(n1106), .A(n756), .S(n773), .Y(n1086) );
  MUX2X1 U1059 ( .B(n1124), .A(n1125), .S(n771), .Y(n1106) );
  MUX2X1 U1060 ( .B(n1107), .A(n1105), .S(SH[2]), .Y(n1087) );
  MUX2X1 U1061 ( .B(n1126), .A(n1127), .S(n771), .Y(n1105) );
  MUX2X1 U1062 ( .B(n1128), .A(n1116), .S(n771), .Y(n1107) );
  MUX2X1 U1063 ( .B(A[12]), .A(A[11]), .S(n761), .Y(n1116) );
  MUX2X1 U1064 ( .B(n799), .A(n1091), .S(n775), .Y(n1056) );
  AND2X1 U1065 ( .A(n1110), .B(n774), .Y(n1091) );
  MUX2X1 U1066 ( .B(n1117), .A(n1118), .S(n771), .Y(n1110) );
  MUX2X1 U1067 ( .B(A[3]), .A(A[2]), .S(n761), .Y(n1118) );
  MUX2X1 U1068 ( .B(A[1]), .A(A[0]), .S(n761), .Y(n1117) );
  MUX2X1 U1069 ( .B(n1111), .A(n1109), .S(n772), .Y(n1092) );
  MUX2X1 U1070 ( .B(n1119), .A(n1120), .S(n771), .Y(n1109) );
  MUX2X1 U1071 ( .B(A[7]), .A(A[6]), .S(n761), .Y(n1120) );
  MUX2X1 U1072 ( .B(A[5]), .A(A[4]), .S(n761), .Y(n1119) );
  MUX2X1 U1073 ( .B(n1121), .A(n1122), .S(n771), .Y(n1111) );
  MUX2X1 U1074 ( .B(A[11]), .A(A[10]), .S(n761), .Y(n1122) );
  MUX2X1 U1075 ( .B(A[9]), .A(A[8]), .S(n761), .Y(n1121) );
  MUX2X1 U1076 ( .B(n796), .A(n1095), .S(n777), .Y(n1060) );
  AND2X1 U1077 ( .A(n1114), .B(n774), .Y(n1095) );
  MUX2X1 U1078 ( .B(n752), .A(n1124), .S(n771), .Y(n1114) );
  MUX2X1 U1079 ( .B(A[2]), .A(A[1]), .S(n761), .Y(n1124) );
  MUX2X1 U1080 ( .B(n1115), .A(n1113), .S(n772), .Y(n1096) );
  MUX2X1 U1081 ( .B(n1125), .A(n1126), .S(n771), .Y(n1113) );
  MUX2X1 U1082 ( .B(A[6]), .A(A[5]), .S(n761), .Y(n1126) );
  MUX2X1 U1083 ( .B(A[4]), .A(A[3]), .S(n758), .Y(n1125) );
  MUX2X1 U1084 ( .B(n1127), .A(n1128), .S(n771), .Y(n1115) );
  MUX2X1 U1085 ( .B(A[10]), .A(A[9]), .S(n761), .Y(n1128) );
  MUX2X1 U1086 ( .B(A[8]), .A(A[7]), .S(n758), .Y(n1127) );
endmodule


module alu_DW_leftsh_1 ( A, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  wire   n570, n569, n568, n567, n566, n565, n564, n563, n562, n561, n560,
         n559, n385, n388, n389, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558;

  AND2X1 U338 ( .A(n388), .B(n401), .Y(n493) );
  OR2X1 U339 ( .A(n430), .B(SH[4]), .Y(n564) );
  INVX1 U340 ( .A(n564), .Y(B[6]) );
  OR2X1 U341 ( .A(SH[4]), .B(n389), .Y(n569) );
  INVX1 U342 ( .A(n569), .Y(B[1]) );
  OR2X1 U343 ( .A(SH[4]), .B(n395), .Y(n570) );
  INVX1 U344 ( .A(n570), .Y(B[0]) );
  OR2X1 U345 ( .A(n385), .B(SH[4]), .Y(n568) );
  INVX1 U346 ( .A(n568), .Y(B[2]) );
  OR2X1 U347 ( .A(n392), .B(SH[4]), .Y(n567) );
  INVX1 U348 ( .A(n567), .Y(B[3]) );
  OR2X1 U349 ( .A(SH[4]), .B(n428), .Y(n562) );
  INVX1 U350 ( .A(n562), .Y(B[8]) );
  OR2X1 U351 ( .A(n432), .B(SH[4]), .Y(n566) );
  INVX1 U352 ( .A(n566), .Y(B[4]) );
  OR2X1 U353 ( .A(SH[4]), .B(n427), .Y(n561) );
  INVX1 U354 ( .A(n561), .Y(B[9]) );
  AND2X1 U355 ( .A(n525), .B(n404), .Y(n452) );
  INVX1 U356 ( .A(n452), .Y(n385) );
  OR2X1 U357 ( .A(n431), .B(SH[4]), .Y(n565) );
  INVX1 U358 ( .A(n565), .Y(B[5]) );
  OR2X1 U359 ( .A(SH[4]), .B(n475), .Y(n560) );
  INVX1 U360 ( .A(n560), .Y(B[10]) );
  OR2X1 U361 ( .A(n393), .B(n397), .Y(n552) );
  INVX1 U362 ( .A(n552), .Y(n388) );
  AND2X1 U363 ( .A(n486), .B(n404), .Y(n515) );
  INVX1 U364 ( .A(n515), .Y(n389) );
  AND2X1 U365 ( .A(n394), .B(n401), .Y(n486) );
  OR2X1 U366 ( .A(n429), .B(SH[4]), .Y(n563) );
  INVX1 U367 ( .A(n563), .Y(B[7]) );
  OR2X1 U368 ( .A(SH[4]), .B(n469), .Y(n559) );
  INVX1 U369 ( .A(n559), .Y(B[11]) );
  AND2X1 U370 ( .A(n520), .B(n404), .Y(n433) );
  INVX1 U371 ( .A(n433), .Y(n392) );
  AND2X1 U372 ( .A(A[0]), .B(n396), .Y(n558) );
  INVX1 U373 ( .A(n558), .Y(n393) );
  OR2X1 U374 ( .A(n546), .B(n397), .Y(n531) );
  INVX1 U375 ( .A(n531), .Y(n394) );
  AND2X1 U376 ( .A(n493), .B(n404), .Y(n532) );
  INVX1 U377 ( .A(n532), .Y(n395) );
  INVX1 U378 ( .A(n487), .Y(n414) );
  INVX1 U379 ( .A(n517), .Y(n417) );
  INVX1 U380 ( .A(n522), .Y(n415) );
  INVX1 U381 ( .A(n494), .Y(n412) );
  INVX1 U382 ( .A(n461), .Y(B[28]) );
  INVX1 U383 ( .A(n470), .Y(n426) );
  INVX1 U384 ( .A(n476), .Y(n425) );
  INVX1 U385 ( .A(n481), .Y(n424) );
  INVX1 U386 ( .A(n488), .Y(n423) );
  INVX1 U387 ( .A(n495), .Y(n422) );
  INVX1 U388 ( .A(n500), .Y(n421) );
  INVX1 U389 ( .A(n510), .Y(n419) );
  INVX1 U390 ( .A(n533), .Y(n411) );
  INVX1 U391 ( .A(n443), .Y(B[30]) );
  INVX1 U392 ( .A(n453), .Y(B[29]) );
  INVX1 U393 ( .A(n516), .Y(n418) );
  INVX1 U394 ( .A(n521), .Y(n416) );
  INVX1 U395 ( .A(n526), .Y(n413) );
  INVX1 U396 ( .A(n505), .Y(n420) );
  INVX1 U397 ( .A(SH[1]), .Y(n399) );
  INVX1 U398 ( .A(n434), .Y(B[31]) );
  INVX1 U399 ( .A(SH[1]), .Y(n400) );
  INVX1 U400 ( .A(n404), .Y(n403) );
  INVX1 U401 ( .A(n404), .Y(n402) );
  INVX1 U402 ( .A(n398), .Y(n397) );
  INVX1 U403 ( .A(SH[0]), .Y(n396) );
  INVX1 U404 ( .A(SH[4]), .Y(n406) );
  INVX1 U405 ( .A(SH[2]), .Y(n401) );
  INVX1 U406 ( .A(SH[1]), .Y(n398) );
  INVX1 U407 ( .A(SH[3]), .Y(n404) );
  INVX1 U408 ( .A(SH[4]), .Y(n405) );
  MUX2X1 U409 ( .B(n435), .A(n436), .S(n406), .Y(n434) );
  MUX2X1 U410 ( .B(n437), .A(n438), .S(n402), .Y(n436) );
  MUX2X1 U411 ( .B(n439), .A(n440), .S(SH[2]), .Y(n437) );
  MUX2X1 U412 ( .B(n441), .A(n442), .S(SH[1]), .Y(n439) );
  MUX2X1 U413 ( .B(A[31]), .A(A[30]), .S(SH[0]), .Y(n441) );
  MUX2X1 U414 ( .B(n444), .A(n445), .S(n405), .Y(n443) );
  MUX2X1 U415 ( .B(n446), .A(n447), .S(n403), .Y(n445) );
  MUX2X1 U416 ( .B(n448), .A(n449), .S(SH[2]), .Y(n446) );
  MUX2X1 U417 ( .B(n450), .A(n451), .S(SH[1]), .Y(n448) );
  MUX2X1 U418 ( .B(A[30]), .A(A[29]), .S(SH[0]), .Y(n450) );
  MUX2X1 U419 ( .B(n454), .A(n455), .S(n405), .Y(n453) );
  MUX2X1 U420 ( .B(n456), .A(n457), .S(n403), .Y(n455) );
  MUX2X1 U421 ( .B(n458), .A(n459), .S(SH[2]), .Y(n456) );
  MUX2X1 U422 ( .B(n442), .A(n460), .S(SH[1]), .Y(n458) );
  MUX2X1 U423 ( .B(A[29]), .A(A[28]), .S(SH[0]), .Y(n442) );
  MUX2X1 U424 ( .B(n462), .A(n463), .S(n405), .Y(n461) );
  MUX2X1 U425 ( .B(n464), .A(n465), .S(n403), .Y(n463) );
  MUX2X1 U426 ( .B(n466), .A(n467), .S(SH[2]), .Y(n464) );
  MUX2X1 U427 ( .B(n451), .A(n468), .S(n397), .Y(n466) );
  MUX2X1 U428 ( .B(A[28]), .A(A[27]), .S(SH[0]), .Y(n451) );
  MUX2X1 U429 ( .B(n469), .A(n426), .S(n405), .Y(B[27]) );
  MUX2X1 U430 ( .B(n471), .A(n472), .S(n403), .Y(n470) );
  MUX2X1 U431 ( .B(n440), .A(n473), .S(SH[2]), .Y(n471) );
  MUX2X1 U432 ( .B(n460), .A(n474), .S(n397), .Y(n440) );
  MUX2X1 U433 ( .B(A[27]), .A(A[26]), .S(SH[0]), .Y(n460) );
  MUX2X1 U434 ( .B(n475), .A(n425), .S(n406), .Y(B[26]) );
  MUX2X1 U435 ( .B(n477), .A(n478), .S(n403), .Y(n476) );
  MUX2X1 U436 ( .B(n449), .A(n479), .S(SH[2]), .Y(n477) );
  MUX2X1 U437 ( .B(n468), .A(n480), .S(n397), .Y(n449) );
  MUX2X1 U438 ( .B(A[26]), .A(A[25]), .S(SH[0]), .Y(n468) );
  MUX2X1 U439 ( .B(n427), .A(n424), .S(n406), .Y(B[25]) );
  MUX2X1 U440 ( .B(n482), .A(n483), .S(n403), .Y(n481) );
  MUX2X1 U441 ( .B(n459), .A(n484), .S(SH[2]), .Y(n482) );
  MUX2X1 U442 ( .B(n474), .A(n485), .S(n397), .Y(n459) );
  MUX2X1 U443 ( .B(A[25]), .A(A[24]), .S(SH[0]), .Y(n474) );
  MUX2X1 U444 ( .B(n414), .A(n486), .S(n403), .Y(n427) );
  MUX2X1 U445 ( .B(n428), .A(n423), .S(n406), .Y(B[24]) );
  MUX2X1 U446 ( .B(n489), .A(n490), .S(n403), .Y(n488) );
  MUX2X1 U447 ( .B(n467), .A(n491), .S(SH[2]), .Y(n489) );
  MUX2X1 U448 ( .B(n480), .A(n492), .S(n397), .Y(n467) );
  MUX2X1 U449 ( .B(A[24]), .A(A[23]), .S(SH[0]), .Y(n480) );
  MUX2X1 U450 ( .B(n412), .A(n493), .S(n403), .Y(n428) );
  MUX2X1 U451 ( .B(n429), .A(n422), .S(n406), .Y(B[23]) );
  MUX2X1 U452 ( .B(n438), .A(n496), .S(n403), .Y(n495) );
  MUX2X1 U453 ( .B(n473), .A(n497), .S(SH[2]), .Y(n438) );
  MUX2X1 U454 ( .B(n485), .A(n498), .S(n397), .Y(n473) );
  MUX2X1 U455 ( .B(A[23]), .A(A[22]), .S(SH[0]), .Y(n485) );
  OR2X1 U456 ( .A(n499), .B(SH[3]), .Y(n429) );
  MUX2X1 U457 ( .B(n430), .A(n421), .S(n406), .Y(B[22]) );
  MUX2X1 U458 ( .B(n447), .A(n501), .S(n402), .Y(n500) );
  MUX2X1 U459 ( .B(n502), .A(n479), .S(n401), .Y(n447) );
  MUX2X1 U460 ( .B(n492), .A(n503), .S(n397), .Y(n479) );
  MUX2X1 U461 ( .B(A[22]), .A(A[21]), .S(SH[0]), .Y(n492) );
  OR2X1 U462 ( .A(n504), .B(n403), .Y(n430) );
  MUX2X1 U463 ( .B(n431), .A(n420), .S(n406), .Y(B[21]) );
  MUX2X1 U464 ( .B(n457), .A(n506), .S(n402), .Y(n505) );
  MUX2X1 U465 ( .B(n484), .A(n507), .S(SH[2]), .Y(n457) );
  MUX2X1 U466 ( .B(n498), .A(n508), .S(n397), .Y(n484) );
  MUX2X1 U467 ( .B(A[21]), .A(A[20]), .S(SH[0]), .Y(n498) );
  OR2X1 U468 ( .A(n509), .B(n403), .Y(n431) );
  MUX2X1 U469 ( .B(n432), .A(n419), .S(n406), .Y(B[20]) );
  MUX2X1 U470 ( .B(n465), .A(n511), .S(n402), .Y(n510) );
  MUX2X1 U471 ( .B(n491), .A(n512), .S(SH[2]), .Y(n465) );
  MUX2X1 U472 ( .B(n503), .A(n513), .S(n397), .Y(n491) );
  MUX2X1 U473 ( .B(A[20]), .A(A[19]), .S(SH[0]), .Y(n503) );
  OR2X1 U474 ( .A(n514), .B(n402), .Y(n432) );
  MUX2X1 U475 ( .B(n392), .A(n418), .S(n406), .Y(B[19]) );
  MUX2X1 U476 ( .B(n472), .A(n517), .S(n402), .Y(n516) );
  MUX2X1 U477 ( .B(n497), .A(n518), .S(SH[2]), .Y(n472) );
  MUX2X1 U478 ( .B(n519), .A(n508), .S(n399), .Y(n497) );
  MUX2X1 U479 ( .B(A[19]), .A(A[18]), .S(SH[0]), .Y(n508) );
  MUX2X1 U480 ( .B(n385), .A(n416), .S(n406), .Y(B[18]) );
  MUX2X1 U481 ( .B(n478), .A(n522), .S(n402), .Y(n521) );
  MUX2X1 U482 ( .B(n502), .A(n523), .S(SH[2]), .Y(n478) );
  MUX2X1 U483 ( .B(n524), .A(n513), .S(n399), .Y(n502) );
  MUX2X1 U484 ( .B(A[18]), .A(A[17]), .S(SH[0]), .Y(n513) );
  MUX2X1 U485 ( .B(n389), .A(n413), .S(n406), .Y(B[17]) );
  MUX2X1 U486 ( .B(n483), .A(n487), .S(n402), .Y(n526) );
  MUX2X1 U487 ( .B(n527), .A(n528), .S(SH[2]), .Y(n487) );
  MUX2X1 U488 ( .B(n507), .A(n529), .S(SH[2]), .Y(n483) );
  MUX2X1 U489 ( .B(n530), .A(n519), .S(n399), .Y(n507) );
  MUX2X1 U490 ( .B(A[17]), .A(A[16]), .S(SH[0]), .Y(n519) );
  MUX2X1 U491 ( .B(n395), .A(n411), .S(n406), .Y(B[16]) );
  MUX2X1 U492 ( .B(n490), .A(n494), .S(n402), .Y(n533) );
  MUX2X1 U493 ( .B(n534), .A(n535), .S(SH[2]), .Y(n494) );
  MUX2X1 U494 ( .B(n512), .A(n536), .S(SH[2]), .Y(n490) );
  MUX2X1 U495 ( .B(n537), .A(n524), .S(n399), .Y(n512) );
  MUX2X1 U496 ( .B(A[16]), .A(A[15]), .S(SH[0]), .Y(n524) );
  AND2X1 U497 ( .A(n435), .B(n405), .Y(B[15]) );
  MUX2X1 U498 ( .B(n499), .A(n496), .S(n404), .Y(n435) );
  MUX2X1 U499 ( .B(n518), .A(n538), .S(SH[2]), .Y(n496) );
  MUX2X1 U500 ( .B(n539), .A(n530), .S(n399), .Y(n518) );
  MUX2X1 U501 ( .B(A[15]), .A(A[14]), .S(SH[0]), .Y(n530) );
  MUX2X1 U502 ( .B(n540), .A(n541), .S(SH[2]), .Y(n499) );
  AND2X1 U503 ( .A(n405), .B(n444), .Y(B[14]) );
  MUX2X1 U504 ( .B(n501), .A(n504), .S(n402), .Y(n444) );
  MUX2X1 U505 ( .B(n542), .A(n543), .S(SH[2]), .Y(n504) );
  MUX2X1 U506 ( .B(n523), .A(n544), .S(SH[2]), .Y(n501) );
  MUX2X1 U507 ( .B(n545), .A(n537), .S(n399), .Y(n523) );
  MUX2X1 U508 ( .B(A[14]), .A(A[13]), .S(SH[0]), .Y(n537) );
  AND2X1 U509 ( .A(n454), .B(n405), .Y(B[13]) );
  MUX2X1 U510 ( .B(n506), .A(n509), .S(n402), .Y(n454) );
  MUX2X1 U511 ( .B(n528), .A(n394), .S(SH[2]), .Y(n509) );
  MUX2X1 U512 ( .B(n547), .A(n548), .S(n399), .Y(n528) );
  MUX2X1 U513 ( .B(n529), .A(n527), .S(SH[2]), .Y(n506) );
  MUX2X1 U514 ( .B(n549), .A(n550), .S(n399), .Y(n527) );
  MUX2X1 U515 ( .B(n551), .A(n539), .S(n399), .Y(n529) );
  MUX2X1 U516 ( .B(A[13]), .A(A[12]), .S(SH[0]), .Y(n539) );
  AND2X1 U517 ( .A(n462), .B(n405), .Y(B[12]) );
  MUX2X1 U518 ( .B(n511), .A(n514), .S(n402), .Y(n462) );
  MUX2X1 U519 ( .B(n535), .A(n388), .S(SH[2]), .Y(n514) );
  MUX2X1 U520 ( .B(n553), .A(n554), .S(n399), .Y(n535) );
  MUX2X1 U521 ( .B(n536), .A(n534), .S(SH[2]), .Y(n511) );
  MUX2X1 U522 ( .B(n555), .A(n556), .S(n399), .Y(n534) );
  MUX2X1 U523 ( .B(n557), .A(n545), .S(n399), .Y(n536) );
  MUX2X1 U524 ( .B(A[12]), .A(A[11]), .S(SH[0]), .Y(n545) );
  MUX2X1 U525 ( .B(n417), .A(n520), .S(n402), .Y(n469) );
  AND2X1 U526 ( .A(n541), .B(n401), .Y(n520) );
  MUX2X1 U527 ( .B(n546), .A(n547), .S(n400), .Y(n541) );
  MUX2X1 U528 ( .B(A[3]), .A(A[2]), .S(SH[0]), .Y(n547) );
  MUX2X1 U529 ( .B(A[1]), .A(A[0]), .S(SH[0]), .Y(n546) );
  MUX2X1 U530 ( .B(n538), .A(n540), .S(SH[2]), .Y(n517) );
  MUX2X1 U531 ( .B(n548), .A(n549), .S(n400), .Y(n540) );
  MUX2X1 U532 ( .B(A[7]), .A(A[6]), .S(SH[0]), .Y(n549) );
  MUX2X1 U533 ( .B(A[5]), .A(A[4]), .S(SH[0]), .Y(n548) );
  MUX2X1 U534 ( .B(n550), .A(n551), .S(n400), .Y(n538) );
  MUX2X1 U535 ( .B(A[11]), .A(A[10]), .S(SH[0]), .Y(n551) );
  MUX2X1 U536 ( .B(A[9]), .A(A[8]), .S(SH[0]), .Y(n550) );
  MUX2X1 U537 ( .B(n415), .A(n525), .S(n403), .Y(n475) );
  AND2X1 U538 ( .A(n543), .B(n401), .Y(n525) );
  MUX2X1 U539 ( .B(n393), .A(n553), .S(n400), .Y(n543) );
  MUX2X1 U540 ( .B(A[2]), .A(A[1]), .S(SH[0]), .Y(n553) );
  MUX2X1 U541 ( .B(n544), .A(n542), .S(SH[2]), .Y(n522) );
  MUX2X1 U542 ( .B(n554), .A(n555), .S(n400), .Y(n542) );
  MUX2X1 U543 ( .B(A[6]), .A(A[5]), .S(SH[0]), .Y(n555) );
  MUX2X1 U544 ( .B(A[4]), .A(A[3]), .S(SH[0]), .Y(n554) );
  MUX2X1 U545 ( .B(n556), .A(n557), .S(n400), .Y(n544) );
  MUX2X1 U546 ( .B(A[10]), .A(A[9]), .S(SH[0]), .Y(n557) );
  MUX2X1 U547 ( .B(A[8]), .A(A[7]), .S(SH[0]), .Y(n556) );
endmodule


module alu_DW_leftsh_2 ( A, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  wire   n572, n571, n570, n569, n568, n567, n566, n565, n564, n563, n562,
         n561, n385, n388, n389, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560;

  AND2X1 U338 ( .A(n388), .B(n403), .Y(n495) );
  OR2X1 U339 ( .A(n432), .B(SH[4]), .Y(n566) );
  INVX1 U340 ( .A(n566), .Y(B[6]) );
  OR2X1 U341 ( .A(n385), .B(SH[4]), .Y(n570) );
  INVX1 U342 ( .A(n570), .Y(B[2]) );
  OR2X1 U343 ( .A(SH[4]), .B(n389), .Y(n571) );
  INVX1 U344 ( .A(n571), .Y(B[1]) );
  OR2X1 U345 ( .A(SH[4]), .B(n395), .Y(n572) );
  INVX1 U346 ( .A(n572), .Y(B[0]) );
  OR2X1 U347 ( .A(n392), .B(SH[4]), .Y(n569) );
  INVX1 U348 ( .A(n569), .Y(B[3]) );
  OR2X1 U349 ( .A(SH[4]), .B(n430), .Y(n564) );
  INVX1 U350 ( .A(n564), .Y(B[8]) );
  OR2X1 U351 ( .A(n434), .B(SH[4]), .Y(n568) );
  INVX1 U352 ( .A(n568), .Y(B[4]) );
  OR2X1 U353 ( .A(SH[4]), .B(n429), .Y(n563) );
  INVX1 U354 ( .A(n563), .Y(B[9]) );
  AND2X1 U355 ( .A(n527), .B(n406), .Y(n454) );
  INVX1 U356 ( .A(n454), .Y(n385) );
  OR2X1 U357 ( .A(n433), .B(SH[4]), .Y(n567) );
  INVX1 U358 ( .A(n567), .Y(B[5]) );
  OR2X1 U359 ( .A(SH[4]), .B(n477), .Y(n562) );
  INVX1 U360 ( .A(n562), .Y(B[10]) );
  OR2X1 U361 ( .A(n393), .B(n399), .Y(n554) );
  INVX1 U362 ( .A(n554), .Y(n388) );
  AND2X1 U363 ( .A(n488), .B(n406), .Y(n517) );
  INVX1 U364 ( .A(n517), .Y(n389) );
  AND2X1 U365 ( .A(n394), .B(n403), .Y(n488) );
  OR2X1 U366 ( .A(n431), .B(SH[4]), .Y(n565) );
  INVX1 U367 ( .A(n565), .Y(B[7]) );
  OR2X1 U368 ( .A(SH[4]), .B(n471), .Y(n561) );
  INVX1 U369 ( .A(n561), .Y(B[11]) );
  AND2X1 U370 ( .A(n522), .B(n406), .Y(n435) );
  INVX1 U371 ( .A(n435), .Y(n392) );
  AND2X1 U372 ( .A(A[0]), .B(n397), .Y(n560) );
  INVX1 U373 ( .A(n560), .Y(n393) );
  OR2X1 U374 ( .A(n548), .B(n399), .Y(n533) );
  INVX1 U375 ( .A(n533), .Y(n394) );
  AND2X1 U376 ( .A(n495), .B(n406), .Y(n534) );
  INVX1 U377 ( .A(n534), .Y(n395) );
  INVX1 U378 ( .A(n436), .Y(B[31]) );
  INVX1 U379 ( .A(n489), .Y(n416) );
  INVX1 U380 ( .A(n519), .Y(n419) );
  INVX1 U381 ( .A(n524), .Y(n417) );
  INVX1 U382 ( .A(n496), .Y(n414) );
  INVX1 U383 ( .A(n472), .Y(n428) );
  INVX1 U384 ( .A(n478), .Y(n427) );
  INVX1 U385 ( .A(n490), .Y(n425) );
  INVX1 U386 ( .A(n507), .Y(n422) );
  INVX1 U387 ( .A(n512), .Y(n421) );
  INVX1 U388 ( .A(n518), .Y(n420) );
  INVX1 U389 ( .A(n523), .Y(n418) );
  INVX1 U390 ( .A(n455), .Y(B[29]) );
  INVX1 U391 ( .A(n463), .Y(B[28]) );
  INVX1 U392 ( .A(n535), .Y(n413) );
  INVX1 U393 ( .A(n403), .Y(n402) );
  INVX1 U394 ( .A(n398), .Y(n401) );
  INVX1 U395 ( .A(n483), .Y(n426) );
  INVX1 U396 ( .A(n528), .Y(n415) );
  INVX1 U397 ( .A(n502), .Y(n423) );
  INVX1 U398 ( .A(n497), .Y(n424) );
  INVX1 U399 ( .A(n445), .Y(B[30]) );
  INVX1 U400 ( .A(n406), .Y(n405) );
  INVX1 U401 ( .A(n406), .Y(n404) );
  INVX1 U402 ( .A(n400), .Y(n399) );
  INVX1 U403 ( .A(n400), .Y(n398) );
  INVX1 U404 ( .A(SH[0]), .Y(n397) );
  INVX1 U405 ( .A(n397), .Y(n396) );
  INVX1 U406 ( .A(SH[4]), .Y(n408) );
  INVX1 U407 ( .A(SH[2]), .Y(n403) );
  INVX1 U408 ( .A(SH[1]), .Y(n400) );
  INVX1 U409 ( .A(SH[3]), .Y(n406) );
  INVX1 U410 ( .A(SH[4]), .Y(n407) );
  MUX2X1 U411 ( .B(n437), .A(n438), .S(n408), .Y(n436) );
  MUX2X1 U412 ( .B(n439), .A(n440), .S(n404), .Y(n438) );
  MUX2X1 U413 ( .B(n441), .A(n442), .S(n402), .Y(n439) );
  MUX2X1 U414 ( .B(n443), .A(n444), .S(n398), .Y(n441) );
  MUX2X1 U415 ( .B(A[31]), .A(A[30]), .S(n396), .Y(n443) );
  MUX2X1 U416 ( .B(n446), .A(n447), .S(n407), .Y(n445) );
  MUX2X1 U417 ( .B(n448), .A(n449), .S(n405), .Y(n447) );
  MUX2X1 U418 ( .B(n450), .A(n451), .S(n402), .Y(n448) );
  MUX2X1 U419 ( .B(n452), .A(n453), .S(n398), .Y(n450) );
  MUX2X1 U420 ( .B(A[30]), .A(A[29]), .S(n396), .Y(n452) );
  MUX2X1 U421 ( .B(n456), .A(n457), .S(n407), .Y(n455) );
  MUX2X1 U422 ( .B(n458), .A(n459), .S(n405), .Y(n457) );
  MUX2X1 U423 ( .B(n460), .A(n461), .S(n402), .Y(n458) );
  MUX2X1 U424 ( .B(n444), .A(n462), .S(n398), .Y(n460) );
  MUX2X1 U425 ( .B(A[29]), .A(A[28]), .S(n396), .Y(n444) );
  MUX2X1 U426 ( .B(n464), .A(n465), .S(n407), .Y(n463) );
  MUX2X1 U427 ( .B(n466), .A(n467), .S(n405), .Y(n465) );
  MUX2X1 U428 ( .B(n468), .A(n469), .S(n402), .Y(n466) );
  MUX2X1 U429 ( .B(n453), .A(n470), .S(n399), .Y(n468) );
  MUX2X1 U430 ( .B(A[28]), .A(A[27]), .S(n396), .Y(n453) );
  MUX2X1 U431 ( .B(n471), .A(n428), .S(n407), .Y(B[27]) );
  MUX2X1 U432 ( .B(n473), .A(n474), .S(n405), .Y(n472) );
  MUX2X1 U433 ( .B(n442), .A(n475), .S(n402), .Y(n473) );
  MUX2X1 U434 ( .B(n462), .A(n476), .S(n399), .Y(n442) );
  MUX2X1 U435 ( .B(A[27]), .A(A[26]), .S(n396), .Y(n462) );
  MUX2X1 U436 ( .B(n477), .A(n427), .S(n408), .Y(B[26]) );
  MUX2X1 U437 ( .B(n479), .A(n480), .S(n405), .Y(n478) );
  MUX2X1 U438 ( .B(n451), .A(n481), .S(n402), .Y(n479) );
  MUX2X1 U439 ( .B(n470), .A(n482), .S(n399), .Y(n451) );
  MUX2X1 U440 ( .B(A[26]), .A(A[25]), .S(n396), .Y(n470) );
  MUX2X1 U441 ( .B(n429), .A(n426), .S(n408), .Y(B[25]) );
  MUX2X1 U442 ( .B(n484), .A(n485), .S(n405), .Y(n483) );
  MUX2X1 U443 ( .B(n461), .A(n486), .S(n402), .Y(n484) );
  MUX2X1 U444 ( .B(n476), .A(n487), .S(n399), .Y(n461) );
  MUX2X1 U445 ( .B(A[25]), .A(A[24]), .S(n396), .Y(n476) );
  MUX2X1 U446 ( .B(n416), .A(n488), .S(n405), .Y(n429) );
  MUX2X1 U447 ( .B(n430), .A(n425), .S(n408), .Y(B[24]) );
  MUX2X1 U448 ( .B(n491), .A(n492), .S(n405), .Y(n490) );
  MUX2X1 U449 ( .B(n469), .A(n493), .S(n402), .Y(n491) );
  MUX2X1 U450 ( .B(n482), .A(n494), .S(n399), .Y(n469) );
  MUX2X1 U451 ( .B(A[24]), .A(A[23]), .S(n396), .Y(n482) );
  MUX2X1 U452 ( .B(n414), .A(n495), .S(n405), .Y(n430) );
  MUX2X1 U453 ( .B(n431), .A(n424), .S(n408), .Y(B[23]) );
  MUX2X1 U454 ( .B(n440), .A(n498), .S(n405), .Y(n497) );
  MUX2X1 U455 ( .B(n475), .A(n499), .S(n402), .Y(n440) );
  MUX2X1 U456 ( .B(n487), .A(n500), .S(n399), .Y(n475) );
  MUX2X1 U457 ( .B(A[23]), .A(A[22]), .S(n396), .Y(n487) );
  OR2X1 U458 ( .A(n501), .B(n405), .Y(n431) );
  MUX2X1 U459 ( .B(n432), .A(n423), .S(n408), .Y(B[22]) );
  MUX2X1 U460 ( .B(n449), .A(n503), .S(n404), .Y(n502) );
  MUX2X1 U461 ( .B(n504), .A(n481), .S(n403), .Y(n449) );
  MUX2X1 U462 ( .B(n494), .A(n505), .S(n399), .Y(n481) );
  MUX2X1 U463 ( .B(A[22]), .A(A[21]), .S(n396), .Y(n494) );
  OR2X1 U464 ( .A(n506), .B(n405), .Y(n432) );
  MUX2X1 U465 ( .B(n433), .A(n422), .S(n408), .Y(B[21]) );
  MUX2X1 U466 ( .B(n459), .A(n508), .S(n404), .Y(n507) );
  MUX2X1 U467 ( .B(n486), .A(n509), .S(n402), .Y(n459) );
  MUX2X1 U468 ( .B(n500), .A(n510), .S(n399), .Y(n486) );
  MUX2X1 U469 ( .B(A[21]), .A(A[20]), .S(n396), .Y(n500) );
  OR2X1 U470 ( .A(n511), .B(n405), .Y(n433) );
  MUX2X1 U471 ( .B(n434), .A(n421), .S(n408), .Y(B[20]) );
  MUX2X1 U472 ( .B(n467), .A(n513), .S(n404), .Y(n512) );
  MUX2X1 U473 ( .B(n493), .A(n514), .S(n402), .Y(n467) );
  MUX2X1 U474 ( .B(n505), .A(n515), .S(n399), .Y(n493) );
  MUX2X1 U475 ( .B(A[20]), .A(A[19]), .S(n396), .Y(n505) );
  OR2X1 U476 ( .A(n516), .B(n405), .Y(n434) );
  MUX2X1 U477 ( .B(n392), .A(n420), .S(n408), .Y(B[19]) );
  MUX2X1 U478 ( .B(n474), .A(n519), .S(n404), .Y(n518) );
  MUX2X1 U479 ( .B(n499), .A(n520), .S(n402), .Y(n474) );
  MUX2X1 U480 ( .B(n521), .A(n510), .S(n401), .Y(n499) );
  MUX2X1 U481 ( .B(A[19]), .A(A[18]), .S(SH[0]), .Y(n510) );
  MUX2X1 U482 ( .B(n385), .A(n418), .S(n408), .Y(B[18]) );
  MUX2X1 U483 ( .B(n480), .A(n524), .S(n404), .Y(n523) );
  MUX2X1 U484 ( .B(n504), .A(n525), .S(n402), .Y(n480) );
  MUX2X1 U485 ( .B(n526), .A(n515), .S(n401), .Y(n504) );
  MUX2X1 U486 ( .B(A[18]), .A(A[17]), .S(SH[0]), .Y(n515) );
  MUX2X1 U487 ( .B(n389), .A(n415), .S(n408), .Y(B[17]) );
  MUX2X1 U488 ( .B(n485), .A(n489), .S(n404), .Y(n528) );
  MUX2X1 U489 ( .B(n529), .A(n530), .S(SH[2]), .Y(n489) );
  MUX2X1 U490 ( .B(n509), .A(n531), .S(n402), .Y(n485) );
  MUX2X1 U491 ( .B(n532), .A(n521), .S(n401), .Y(n509) );
  MUX2X1 U492 ( .B(A[17]), .A(A[16]), .S(SH[0]), .Y(n521) );
  MUX2X1 U493 ( .B(n395), .A(n413), .S(n408), .Y(B[16]) );
  MUX2X1 U494 ( .B(n492), .A(n496), .S(n404), .Y(n535) );
  MUX2X1 U495 ( .B(n536), .A(n537), .S(SH[2]), .Y(n496) );
  MUX2X1 U496 ( .B(n514), .A(n538), .S(n402), .Y(n492) );
  MUX2X1 U497 ( .B(n539), .A(n526), .S(n401), .Y(n514) );
  MUX2X1 U498 ( .B(A[16]), .A(A[15]), .S(SH[0]), .Y(n526) );
  AND2X1 U499 ( .A(n437), .B(n407), .Y(B[15]) );
  MUX2X1 U500 ( .B(n501), .A(n498), .S(n406), .Y(n437) );
  MUX2X1 U501 ( .B(n520), .A(n540), .S(SH[2]), .Y(n498) );
  MUX2X1 U502 ( .B(n541), .A(n532), .S(n401), .Y(n520) );
  MUX2X1 U503 ( .B(A[15]), .A(A[14]), .S(SH[0]), .Y(n532) );
  MUX2X1 U504 ( .B(n542), .A(n543), .S(SH[2]), .Y(n501) );
  AND2X1 U505 ( .A(n407), .B(n446), .Y(B[14]) );
  MUX2X1 U506 ( .B(n503), .A(n506), .S(n404), .Y(n446) );
  MUX2X1 U507 ( .B(n544), .A(n545), .S(SH[2]), .Y(n506) );
  MUX2X1 U508 ( .B(n525), .A(n546), .S(SH[2]), .Y(n503) );
  MUX2X1 U509 ( .B(n547), .A(n539), .S(n401), .Y(n525) );
  MUX2X1 U510 ( .B(A[14]), .A(A[13]), .S(SH[0]), .Y(n539) );
  AND2X1 U511 ( .A(n456), .B(n407), .Y(B[13]) );
  MUX2X1 U512 ( .B(n508), .A(n511), .S(n404), .Y(n456) );
  MUX2X1 U513 ( .B(n530), .A(n394), .S(n402), .Y(n511) );
  MUX2X1 U514 ( .B(n549), .A(n550), .S(n401), .Y(n530) );
  MUX2X1 U515 ( .B(n531), .A(n529), .S(n402), .Y(n508) );
  MUX2X1 U516 ( .B(n551), .A(n552), .S(n401), .Y(n529) );
  MUX2X1 U517 ( .B(n553), .A(n541), .S(n401), .Y(n531) );
  MUX2X1 U518 ( .B(A[13]), .A(A[12]), .S(SH[0]), .Y(n541) );
  AND2X1 U519 ( .A(n464), .B(n407), .Y(B[12]) );
  MUX2X1 U520 ( .B(n513), .A(n516), .S(n404), .Y(n464) );
  MUX2X1 U521 ( .B(n537), .A(n388), .S(n402), .Y(n516) );
  MUX2X1 U522 ( .B(n555), .A(n556), .S(n401), .Y(n537) );
  MUX2X1 U523 ( .B(n538), .A(n536), .S(SH[2]), .Y(n513) );
  MUX2X1 U524 ( .B(n557), .A(n558), .S(n401), .Y(n536) );
  MUX2X1 U525 ( .B(n559), .A(n547), .S(n401), .Y(n538) );
  MUX2X1 U526 ( .B(A[12]), .A(A[11]), .S(SH[0]), .Y(n547) );
  MUX2X1 U527 ( .B(n419), .A(n522), .S(n404), .Y(n471) );
  AND2X1 U528 ( .A(n543), .B(n403), .Y(n522) );
  MUX2X1 U529 ( .B(n548), .A(n549), .S(n400), .Y(n543) );
  MUX2X1 U530 ( .B(A[3]), .A(A[2]), .S(SH[0]), .Y(n549) );
  MUX2X1 U531 ( .B(A[1]), .A(A[0]), .S(SH[0]), .Y(n548) );
  MUX2X1 U532 ( .B(n540), .A(n542), .S(n402), .Y(n519) );
  MUX2X1 U533 ( .B(n550), .A(n551), .S(n400), .Y(n542) );
  MUX2X1 U534 ( .B(A[7]), .A(A[6]), .S(SH[0]), .Y(n551) );
  MUX2X1 U535 ( .B(A[5]), .A(A[4]), .S(SH[0]), .Y(n550) );
  MUX2X1 U536 ( .B(n552), .A(n553), .S(n400), .Y(n540) );
  MUX2X1 U537 ( .B(A[11]), .A(A[10]), .S(n396), .Y(n553) );
  MUX2X1 U538 ( .B(A[9]), .A(A[8]), .S(SH[0]), .Y(n552) );
  MUX2X1 U539 ( .B(n417), .A(n527), .S(n405), .Y(n477) );
  AND2X1 U540 ( .A(n545), .B(n403), .Y(n527) );
  MUX2X1 U541 ( .B(n393), .A(n555), .S(n400), .Y(n545) );
  MUX2X1 U542 ( .B(A[2]), .A(A[1]), .S(SH[0]), .Y(n555) );
  MUX2X1 U543 ( .B(n546), .A(n544), .S(n402), .Y(n524) );
  MUX2X1 U544 ( .B(n556), .A(n557), .S(n400), .Y(n544) );
  MUX2X1 U545 ( .B(A[6]), .A(A[5]), .S(SH[0]), .Y(n557) );
  MUX2X1 U546 ( .B(A[4]), .A(A[3]), .S(SH[0]), .Y(n556) );
  MUX2X1 U547 ( .B(n558), .A(n559), .S(n400), .Y(n546) );
  MUX2X1 U548 ( .B(A[10]), .A(A[9]), .S(SH[0]), .Y(n559) );
  MUX2X1 U549 ( .B(A[8]), .A(A[7]), .S(SH[0]), .Y(n558) );
endmodule


module alu_DW_leftsh_15 ( A, SH, B );
  input [63:0] A;
  input [5:0] SH;
  output [63:0] B;
  wire   n1305, n1304, n1303, n1302, n1301, n1300, n1299, n1298, n1297, n1296,
         n1295, n1294, n1293, n1292, n1291, n1290, n1289, n1288, n1287, n1286,
         n1285, n1284, n1283, n1282, n1281, n1280, n1279, n1278, n1277, n1276,
         n1275, n1274, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n914, n915, n916, n918,
         n919, n920, n922, n923, n924, n925, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273;

  AND2X1 U801 ( .A(n905), .B(n949), .Y(n1071) );
  OR2X1 U802 ( .A(n903), .B(n951), .Y(n1296) );
  INVX1 U803 ( .A(n1296), .Y(B[9]) );
  OR2X1 U804 ( .A(n900), .B(n951), .Y(n1299) );
  INVX1 U805 ( .A(n1299), .Y(B[6]) );
  OR2X1 U806 ( .A(n952), .B(n1037), .Y(n1283) );
  INVX1 U807 ( .A(n1283), .Y(B[22]) );
  OR2X1 U808 ( .A(n952), .B(n935), .Y(n1301) );
  INVX1 U809 ( .A(n1301), .Y(B[4]) );
  OR2X1 U810 ( .A(n912), .B(n951), .Y(n1302) );
  INVX1 U811 ( .A(n1302), .Y(B[3]) );
  OR2X1 U812 ( .A(n952), .B(n1051), .Y(n1285) );
  INVX1 U813 ( .A(n1285), .Y(B[20]) );
  OR2X1 U814 ( .A(n916), .B(n952), .Y(n1294) );
  INVX1 U815 ( .A(n1294), .Y(B[11]) );
  OR2X1 U816 ( .A(n899), .B(n951), .Y(n1297) );
  INVX1 U817 ( .A(n1297), .Y(B[8]) );
  OR2X1 U818 ( .A(n901), .B(n951), .Y(n1300) );
  INVX1 U819 ( .A(n1300), .Y(B[5]) );
  OR2X1 U820 ( .A(n902), .B(n952), .Y(n1303) );
  INVX1 U821 ( .A(n1303), .Y(B[2]) );
  OR2X1 U822 ( .A(n952), .B(n988), .Y(n1277) );
  INVX1 U823 ( .A(n1277), .Y(B[28]) );
  OR2X1 U824 ( .A(n1014), .B(n952), .Y(n1280) );
  INVX1 U825 ( .A(n1280), .Y(B[25]) );
  OR2X1 U826 ( .A(n1022), .B(n952), .Y(n1281) );
  INVX1 U827 ( .A(n1281), .Y(B[24]) );
  OR2X1 U828 ( .A(n952), .B(n1044), .Y(n1284) );
  INVX1 U829 ( .A(n1284), .Y(B[21]) );
  OR2X1 U830 ( .A(n952), .B(n897), .Y(n1304) );
  INVX1 U831 ( .A(n1304), .Y(B[1]) );
  OR2X1 U832 ( .A(n952), .B(n1065), .Y(n1287) );
  INVX1 U833 ( .A(n1287), .Y(B[18]) );
  OR2X1 U834 ( .A(n951), .B(n1073), .Y(n1288) );
  INVX1 U835 ( .A(n1288), .Y(B[17]) );
  OR2X1 U836 ( .A(n952), .B(n1080), .Y(n1289) );
  INVX1 U837 ( .A(n1289), .Y(B[16]) );
  OR2X1 U838 ( .A(n908), .B(n952), .Y(n1290) );
  INVX1 U839 ( .A(n1290), .Y(B[15]) );
  OR2X1 U840 ( .A(n910), .B(n952), .Y(n1291) );
  INVX1 U841 ( .A(n1291), .Y(B[14]) );
  OR2X1 U842 ( .A(n906), .B(n952), .Y(n1292) );
  INVX1 U843 ( .A(n1292), .Y(B[13]) );
  OR2X1 U844 ( .A(n951), .B(n925), .Y(n1293) );
  INVX1 U845 ( .A(n1293), .Y(B[12]) );
  OR2X1 U846 ( .A(n904), .B(n952), .Y(n1295) );
  INVX1 U847 ( .A(n1295), .Y(B[10]) );
  OR2X1 U848 ( .A(n951), .B(n898), .Y(n1305) );
  INVX1 U849 ( .A(n1305), .Y(B[0]) );
  AND2X1 U850 ( .A(n911), .B(n949), .Y(n1172) );
  INVX1 U851 ( .A(n1172), .Y(n897) );
  AND2X1 U852 ( .A(n914), .B(n949), .Y(n1178) );
  INVX1 U853 ( .A(n1178), .Y(n898) );
  AND2X1 U854 ( .A(n1129), .B(n949), .Y(n955) );
  INVX1 U855 ( .A(n955), .Y(n899) );
  AND2X1 U856 ( .A(n918), .B(n949), .Y(n957) );
  INVX1 U857 ( .A(n957), .Y(n900) );
  AND2X1 U858 ( .A(n907), .B(n949), .Y(n996) );
  INVX1 U859 ( .A(n996), .Y(n901) );
  AND2X1 U860 ( .A(n909), .B(n949), .Y(n1166) );
  INVX1 U861 ( .A(n1166), .Y(n902) );
  AND2X1 U862 ( .A(n1123), .B(n949), .Y(n954) );
  INVX1 U863 ( .A(n954), .Y(n903) );
  AND2X1 U864 ( .A(n1204), .B(n949), .Y(n1117) );
  INVX1 U865 ( .A(n1117), .Y(n904) );
  OR2X1 U866 ( .A(n1233), .B(SH[3]), .Y(n1154) );
  INVX1 U867 ( .A(n1154), .Y(n905) );
  AND2X1 U868 ( .A(n1192), .B(n949), .Y(n1099) );
  INVX1 U869 ( .A(n1099), .Y(n906) );
  OR2X1 U870 ( .A(n1229), .B(SH[3]), .Y(n1148) );
  INVX1 U871 ( .A(n1148), .Y(n907) );
  AND2X1 U872 ( .A(n1183), .B(n949), .Y(n1087) );
  INVX1 U873 ( .A(n1087), .Y(n908) );
  OR2X1 U874 ( .A(n924), .B(n948), .Y(n1191) );
  INVX1 U875 ( .A(n1191), .Y(n909) );
  AND2X1 U876 ( .A(n1187), .B(n949), .Y(n1093) );
  INVX1 U877 ( .A(n1093), .Y(n910) );
  OR2X1 U878 ( .A(n915), .B(n947), .Y(n1234) );
  INVX1 U879 ( .A(n1234), .Y(n911) );
  AND2X1 U880 ( .A(n923), .B(n949), .Y(n1134) );
  INVX1 U881 ( .A(n1134), .Y(n912) );
  OR2X1 U882 ( .A(n920), .B(n951), .Y(n1298) );
  INVX1 U883 ( .A(n1298), .Y(B[7]) );
  OR2X1 U884 ( .A(n919), .B(SH[3]), .Y(n1248) );
  INVX1 U885 ( .A(n1248), .Y(n914) );
  AND2X1 U886 ( .A(n931), .B(n944), .Y(n1212) );
  INVX1 U887 ( .A(n1212), .Y(n915) );
  AND2X1 U888 ( .A(n1200), .B(n949), .Y(n1111) );
  INVX1 U889 ( .A(n1111), .Y(n916) );
  OR2X1 U890 ( .A(n952), .B(n1058), .Y(n1286) );
  INVX1 U891 ( .A(n1286), .Y(B[19]) );
  OR2X1 U892 ( .A(n1225), .B(SH[3]), .Y(n1142) );
  INVX1 U893 ( .A(n1142), .Y(n918) );
  AND2X1 U894 ( .A(n922), .B(n944), .Y(n1217) );
  INVX1 U895 ( .A(n1217), .Y(n919) );
  AND2X1 U896 ( .A(n932), .B(n949), .Y(n956) );
  INVX1 U897 ( .A(n956), .Y(n920) );
  OR2X1 U898 ( .A(n952), .B(n1030), .Y(n1282) );
  INVX1 U899 ( .A(n1282), .Y(B[23]) );
  OR2X1 U900 ( .A(n933), .B(n938), .Y(n1267) );
  INVX1 U901 ( .A(n1267), .Y(n922) );
  OR2X1 U902 ( .A(n934), .B(n947), .Y(n1160) );
  INVX1 U903 ( .A(n1160), .Y(n923) );
  AND2X1 U904 ( .A(n1257), .B(n944), .Y(n1242) );
  INVX1 U905 ( .A(n1242), .Y(n924) );
  AND2X1 U906 ( .A(n1196), .B(n949), .Y(n1105) );
  INVX1 U907 ( .A(n1105), .Y(n925) );
  OR2X1 U908 ( .A(n998), .B(n951), .Y(n1278) );
  INVX1 U909 ( .A(n1278), .Y(B[27]) );
  OR2X1 U910 ( .A(n952), .B(n959), .Y(n1274) );
  INVX1 U911 ( .A(n1274), .Y(B[31]) );
  OR2X1 U912 ( .A(n952), .B(n979), .Y(n1276) );
  INVX1 U913 ( .A(n1276), .Y(B[29]) );
  OR2X1 U914 ( .A(n1006), .B(n952), .Y(n1279) );
  INVX1 U915 ( .A(n1279), .Y(B[26]) );
  OR2X1 U916 ( .A(n969), .B(n952), .Y(n1275) );
  INVX1 U917 ( .A(n1275), .Y(B[30]) );
  OR2X1 U918 ( .A(n1263), .B(n938), .Y(n1247) );
  INVX1 U919 ( .A(n1247), .Y(n931) );
  OR2X1 U920 ( .A(n1221), .B(SH[3]), .Y(n1136) );
  INVX1 U921 ( .A(n1136), .Y(n932) );
  AND2X1 U922 ( .A(A[0]), .B(n936), .Y(n1273) );
  INVX1 U923 ( .A(n1273), .Y(n933) );
  AND2X1 U924 ( .A(n1253), .B(n944), .Y(n1238) );
  INVX1 U925 ( .A(n1238), .Y(n934) );
  INVX1 U926 ( .A(n1071), .Y(n935) );
  INVX1 U927 ( .A(n946), .Y(n947) );
  INVX1 U928 ( .A(n946), .Y(n948) );
  INVX1 U929 ( .A(n939), .Y(n940) );
  INVX1 U930 ( .A(n939), .Y(n941) );
  INVX1 U931 ( .A(n939), .Y(n943) );
  INVX1 U932 ( .A(n939), .Y(n942) );
  INVX1 U933 ( .A(SH[0]), .Y(n937) );
  INVX1 U934 ( .A(SH[2]), .Y(n945) );
  MUX2X1 U935 ( .B(n976), .A(n995), .S(n938), .Y(n994) );
  INVX1 U936 ( .A(SH[0]), .Y(n936) );
  INVX1 U937 ( .A(n939), .Y(n938) );
  INVX1 U938 ( .A(SH[1]), .Y(n939) );
  INVX1 U939 ( .A(SH[2]), .Y(n944) );
  INVX1 U940 ( .A(SH[3]), .Y(n946) );
  INVX1 U941 ( .A(SH[4]), .Y(n949) );
  INVX1 U942 ( .A(n953), .Y(n952) );
  INVX1 U943 ( .A(n953), .Y(n951) );
  INVX1 U944 ( .A(n953), .Y(n950) );
  INVX1 U945 ( .A(SH[5]), .Y(n953) );
  MUX2X1 U946 ( .B(n958), .A(n959), .S(n951), .Y(B[63]) );
  MUX2X1 U947 ( .B(n960), .A(n961), .S(n949), .Y(n958) );
  MUX2X1 U948 ( .B(n962), .A(n963), .S(n946), .Y(n961) );
  MUX2X1 U949 ( .B(n964), .A(n965), .S(n945), .Y(n963) );
  MUX2X1 U950 ( .B(n966), .A(n967), .S(n939), .Y(n965) );
  MUX2X1 U951 ( .B(A[62]), .A(A[63]), .S(n937), .Y(n967) );
  MUX2X1 U952 ( .B(n968), .A(n969), .S(n951), .Y(B[62]) );
  MUX2X1 U953 ( .B(n970), .A(n971), .S(n949), .Y(n968) );
  MUX2X1 U954 ( .B(n972), .A(n973), .S(n946), .Y(n971) );
  MUX2X1 U955 ( .B(n974), .A(n975), .S(n944), .Y(n973) );
  MUX2X1 U956 ( .B(n976), .A(n977), .S(n939), .Y(n975) );
  MUX2X1 U957 ( .B(A[61]), .A(A[62]), .S(n936), .Y(n977) );
  MUX2X1 U958 ( .B(n978), .A(n979), .S(n951), .Y(B[61]) );
  MUX2X1 U959 ( .B(n980), .A(n981), .S(n949), .Y(n978) );
  MUX2X1 U960 ( .B(n982), .A(n983), .S(n946), .Y(n981) );
  MUX2X1 U961 ( .B(n984), .A(n985), .S(n945), .Y(n983) );
  MUX2X1 U962 ( .B(n986), .A(n966), .S(n939), .Y(n985) );
  MUX2X1 U963 ( .B(A[60]), .A(A[61]), .S(n936), .Y(n966) );
  MUX2X1 U964 ( .B(n987), .A(n988), .S(n951), .Y(B[60]) );
  MUX2X1 U965 ( .B(n989), .A(n990), .S(n949), .Y(n987) );
  MUX2X1 U966 ( .B(n991), .A(n992), .S(n946), .Y(n990) );
  MUX2X1 U967 ( .B(n993), .A(n994), .S(n945), .Y(n992) );
  MUX2X1 U968 ( .B(A[59]), .A(A[60]), .S(n936), .Y(n976) );
  MUX2X1 U969 ( .B(n997), .A(n998), .S(n951), .Y(B[59]) );
  MUX2X1 U970 ( .B(n999), .A(n1000), .S(n949), .Y(n997) );
  MUX2X1 U971 ( .B(n1001), .A(n1002), .S(n946), .Y(n1000) );
  MUX2X1 U972 ( .B(n1003), .A(n964), .S(n945), .Y(n1002) );
  MUX2X1 U973 ( .B(n986), .A(n1004), .S(n940), .Y(n964) );
  MUX2X1 U974 ( .B(A[58]), .A(A[59]), .S(n936), .Y(n986) );
  MUX2X1 U975 ( .B(n1005), .A(n1006), .S(n951), .Y(B[58]) );
  MUX2X1 U976 ( .B(n1007), .A(n1008), .S(n949), .Y(n1005) );
  MUX2X1 U977 ( .B(n1009), .A(n1010), .S(n946), .Y(n1008) );
  MUX2X1 U978 ( .B(n1011), .A(n974), .S(n944), .Y(n1010) );
  MUX2X1 U979 ( .B(n995), .A(n1012), .S(n938), .Y(n974) );
  MUX2X1 U980 ( .B(A[57]), .A(A[58]), .S(n936), .Y(n995) );
  MUX2X1 U981 ( .B(n1013), .A(n1014), .S(n951), .Y(B[57]) );
  MUX2X1 U982 ( .B(n1015), .A(n1016), .S(n949), .Y(n1013) );
  MUX2X1 U983 ( .B(n1017), .A(n1018), .S(n946), .Y(n1016) );
  MUX2X1 U984 ( .B(n1019), .A(n984), .S(n945), .Y(n1018) );
  MUX2X1 U985 ( .B(n1004), .A(n1020), .S(n938), .Y(n984) );
  MUX2X1 U986 ( .B(A[56]), .A(A[57]), .S(n936), .Y(n1004) );
  MUX2X1 U987 ( .B(n1021), .A(n1022), .S(n951), .Y(B[56]) );
  MUX2X1 U988 ( .B(n1023), .A(n1024), .S(n949), .Y(n1021) );
  MUX2X1 U989 ( .B(n1025), .A(n1026), .S(n946), .Y(n1024) );
  MUX2X1 U990 ( .B(n1027), .A(n993), .S(n944), .Y(n1026) );
  MUX2X1 U991 ( .B(n1012), .A(n1028), .S(n938), .Y(n993) );
  MUX2X1 U992 ( .B(A[55]), .A(A[56]), .S(n936), .Y(n1012) );
  MUX2X1 U993 ( .B(n1029), .A(n1030), .S(n952), .Y(B[55]) );
  MUX2X1 U994 ( .B(n1031), .A(n1032), .S(n949), .Y(n1029) );
  MUX2X1 U995 ( .B(n1033), .A(n962), .S(n946), .Y(n1032) );
  MUX2X1 U996 ( .B(n1034), .A(n1003), .S(n944), .Y(n962) );
  MUX2X1 U997 ( .B(n1020), .A(n1035), .S(n938), .Y(n1003) );
  MUX2X1 U998 ( .B(A[54]), .A(A[55]), .S(n936), .Y(n1020) );
  MUX2X1 U999 ( .B(n1036), .A(n1037), .S(n951), .Y(B[54]) );
  MUX2X1 U1000 ( .B(n1038), .A(n1039), .S(n949), .Y(n1036) );
  MUX2X1 U1001 ( .B(n1040), .A(n972), .S(n946), .Y(n1039) );
  MUX2X1 U1002 ( .B(n1041), .A(n1011), .S(n944), .Y(n972) );
  MUX2X1 U1003 ( .B(n1028), .A(n1042), .S(n938), .Y(n1011) );
  MUX2X1 U1004 ( .B(A[53]), .A(A[54]), .S(n936), .Y(n1028) );
  MUX2X1 U1005 ( .B(n1043), .A(n1044), .S(n950), .Y(B[53]) );
  MUX2X1 U1006 ( .B(n1045), .A(n1046), .S(n949), .Y(n1043) );
  MUX2X1 U1007 ( .B(n1047), .A(n982), .S(n946), .Y(n1046) );
  MUX2X1 U1008 ( .B(n1048), .A(n1019), .S(n944), .Y(n982) );
  MUX2X1 U1009 ( .B(n1035), .A(n1049), .S(n938), .Y(n1019) );
  MUX2X1 U1010 ( .B(A[52]), .A(A[53]), .S(n936), .Y(n1035) );
  MUX2X1 U1011 ( .B(n1050), .A(n1051), .S(n951), .Y(B[52]) );
  MUX2X1 U1012 ( .B(n1052), .A(n1053), .S(n949), .Y(n1050) );
  MUX2X1 U1013 ( .B(n1054), .A(n991), .S(n946), .Y(n1053) );
  MUX2X1 U1014 ( .B(n1055), .A(n1027), .S(n944), .Y(n991) );
  MUX2X1 U1015 ( .B(n1042), .A(n1056), .S(n938), .Y(n1027) );
  MUX2X1 U1016 ( .B(A[51]), .A(A[52]), .S(n936), .Y(n1042) );
  MUX2X1 U1017 ( .B(n1057), .A(n1058), .S(n950), .Y(B[51]) );
  MUX2X1 U1018 ( .B(n1059), .A(n1060), .S(n949), .Y(n1057) );
  MUX2X1 U1019 ( .B(n1061), .A(n1001), .S(n946), .Y(n1060) );
  MUX2X1 U1020 ( .B(n1062), .A(n1034), .S(n945), .Y(n1001) );
  MUX2X1 U1021 ( .B(n1049), .A(n1063), .S(n938), .Y(n1034) );
  MUX2X1 U1022 ( .B(A[50]), .A(A[51]), .S(n937), .Y(n1049) );
  MUX2X1 U1023 ( .B(n1064), .A(n1065), .S(n951), .Y(B[50]) );
  MUX2X1 U1024 ( .B(n1066), .A(n1067), .S(n949), .Y(n1064) );
  MUX2X1 U1025 ( .B(n1068), .A(n1009), .S(n946), .Y(n1067) );
  MUX2X1 U1026 ( .B(n1069), .A(n1041), .S(n944), .Y(n1009) );
  MUX2X1 U1027 ( .B(n1056), .A(n1070), .S(n943), .Y(n1041) );
  MUX2X1 U1028 ( .B(A[49]), .A(A[50]), .S(n936), .Y(n1056) );
  MUX2X1 U1029 ( .B(n1072), .A(n1073), .S(n950), .Y(B[49]) );
  MUX2X1 U1030 ( .B(n1074), .A(n1075), .S(n949), .Y(n1072) );
  MUX2X1 U1031 ( .B(n1076), .A(n1017), .S(n946), .Y(n1075) );
  MUX2X1 U1032 ( .B(n1077), .A(n1048), .S(n944), .Y(n1017) );
  MUX2X1 U1033 ( .B(n1063), .A(n1078), .S(n938), .Y(n1048) );
  MUX2X1 U1034 ( .B(A[48]), .A(A[49]), .S(n937), .Y(n1063) );
  MUX2X1 U1035 ( .B(n1079), .A(n1080), .S(n950), .Y(B[48]) );
  MUX2X1 U1036 ( .B(n1081), .A(n1082), .S(n949), .Y(n1079) );
  MUX2X1 U1037 ( .B(n1083), .A(n1025), .S(n946), .Y(n1082) );
  MUX2X1 U1038 ( .B(n1084), .A(n1055), .S(n944), .Y(n1025) );
  MUX2X1 U1039 ( .B(n1070), .A(n1085), .S(n943), .Y(n1055) );
  MUX2X1 U1040 ( .B(A[47]), .A(A[48]), .S(n937), .Y(n1070) );
  MUX2X1 U1041 ( .B(n1086), .A(n908), .S(n950), .Y(B[47]) );
  MUX2X1 U1042 ( .B(n1088), .A(n960), .S(n949), .Y(n1086) );
  MUX2X1 U1043 ( .B(n1033), .A(n1089), .S(n948), .Y(n960) );
  MUX2X1 U1044 ( .B(n1090), .A(n1062), .S(n944), .Y(n1033) );
  MUX2X1 U1045 ( .B(n1078), .A(n1091), .S(n938), .Y(n1062) );
  MUX2X1 U1046 ( .B(A[46]), .A(A[47]), .S(n936), .Y(n1078) );
  MUX2X1 U1047 ( .B(n1092), .A(n910), .S(n950), .Y(B[46]) );
  MUX2X1 U1048 ( .B(n1094), .A(n970), .S(n949), .Y(n1092) );
  MUX2X1 U1049 ( .B(n1040), .A(n1095), .S(SH[3]), .Y(n970) );
  MUX2X1 U1050 ( .B(n1096), .A(n1069), .S(n944), .Y(n1040) );
  MUX2X1 U1051 ( .B(n1085), .A(n1097), .S(n943), .Y(n1069) );
  MUX2X1 U1052 ( .B(A[45]), .A(A[46]), .S(n936), .Y(n1085) );
  MUX2X1 U1053 ( .B(n1098), .A(n906), .S(n950), .Y(B[45]) );
  MUX2X1 U1054 ( .B(n1100), .A(n980), .S(n949), .Y(n1098) );
  MUX2X1 U1055 ( .B(n1047), .A(n1101), .S(SH[3]), .Y(n980) );
  MUX2X1 U1056 ( .B(n1102), .A(n1077), .S(n944), .Y(n1047) );
  MUX2X1 U1057 ( .B(n1091), .A(n1103), .S(n943), .Y(n1077) );
  MUX2X1 U1058 ( .B(A[44]), .A(A[45]), .S(n936), .Y(n1091) );
  MUX2X1 U1059 ( .B(n1104), .A(n925), .S(n950), .Y(B[44]) );
  MUX2X1 U1060 ( .B(n1106), .A(n989), .S(n949), .Y(n1104) );
  MUX2X1 U1061 ( .B(n1054), .A(n1107), .S(SH[3]), .Y(n989) );
  MUX2X1 U1062 ( .B(n1108), .A(n1084), .S(n944), .Y(n1054) );
  MUX2X1 U1063 ( .B(n1097), .A(n1109), .S(n943), .Y(n1084) );
  MUX2X1 U1064 ( .B(A[43]), .A(A[44]), .S(n936), .Y(n1097) );
  MUX2X1 U1065 ( .B(n1110), .A(n916), .S(n950), .Y(B[43]) );
  MUX2X1 U1066 ( .B(n1112), .A(n999), .S(n949), .Y(n1110) );
  MUX2X1 U1067 ( .B(n1061), .A(n1113), .S(SH[3]), .Y(n999) );
  MUX2X1 U1068 ( .B(n1114), .A(n1090), .S(n944), .Y(n1061) );
  MUX2X1 U1069 ( .B(n1103), .A(n1115), .S(n943), .Y(n1090) );
  MUX2X1 U1070 ( .B(A[42]), .A(A[43]), .S(n937), .Y(n1103) );
  MUX2X1 U1071 ( .B(n1116), .A(n904), .S(n951), .Y(B[42]) );
  MUX2X1 U1072 ( .B(n1118), .A(n1007), .S(n949), .Y(n1116) );
  MUX2X1 U1073 ( .B(n1068), .A(n1119), .S(SH[3]), .Y(n1007) );
  MUX2X1 U1074 ( .B(n1120), .A(n1096), .S(n944), .Y(n1068) );
  MUX2X1 U1075 ( .B(n1109), .A(n1121), .S(n943), .Y(n1096) );
  MUX2X1 U1076 ( .B(A[41]), .A(A[42]), .S(n936), .Y(n1109) );
  MUX2X1 U1077 ( .B(n1122), .A(n903), .S(n951), .Y(B[41]) );
  MUX2X1 U1078 ( .B(n1124), .A(n1015), .S(n949), .Y(n1122) );
  MUX2X1 U1079 ( .B(n1076), .A(n1125), .S(SH[3]), .Y(n1015) );
  MUX2X1 U1080 ( .B(n1126), .A(n1102), .S(n944), .Y(n1076) );
  MUX2X1 U1081 ( .B(n1115), .A(n1127), .S(n943), .Y(n1102) );
  MUX2X1 U1082 ( .B(A[40]), .A(A[41]), .S(n936), .Y(n1115) );
  MUX2X1 U1083 ( .B(n1128), .A(n899), .S(n951), .Y(B[40]) );
  MUX2X1 U1084 ( .B(n1130), .A(n1023), .S(n949), .Y(n1128) );
  MUX2X1 U1085 ( .B(n1083), .A(n1131), .S(SH[3]), .Y(n1023) );
  MUX2X1 U1086 ( .B(n1132), .A(n1108), .S(n944), .Y(n1083) );
  MUX2X1 U1087 ( .B(n1121), .A(n1133), .S(n943), .Y(n1108) );
  MUX2X1 U1088 ( .B(A[39]), .A(A[40]), .S(n937), .Y(n1121) );
  MUX2X1 U1089 ( .B(n1135), .A(n920), .S(n951), .Y(B[39]) );
  MUX2X1 U1090 ( .B(n1137), .A(n1031), .S(n949), .Y(n1135) );
  MUX2X1 U1091 ( .B(n1089), .A(n1138), .S(SH[3]), .Y(n1031) );
  MUX2X1 U1092 ( .B(n1139), .A(n1114), .S(n944), .Y(n1089) );
  MUX2X1 U1093 ( .B(n1127), .A(n1140), .S(n943), .Y(n1114) );
  MUX2X1 U1094 ( .B(A[38]), .A(A[39]), .S(n936), .Y(n1127) );
  MUX2X1 U1095 ( .B(n1141), .A(n900), .S(n951), .Y(B[38]) );
  MUX2X1 U1096 ( .B(n1143), .A(n1038), .S(n949), .Y(n1141) );
  MUX2X1 U1097 ( .B(n1095), .A(n1144), .S(SH[3]), .Y(n1038) );
  MUX2X1 U1098 ( .B(n1145), .A(n1120), .S(n945), .Y(n1095) );
  MUX2X1 U1099 ( .B(n1133), .A(n1146), .S(n943), .Y(n1120) );
  MUX2X1 U1100 ( .B(A[37]), .A(A[38]), .S(n937), .Y(n1133) );
  MUX2X1 U1101 ( .B(n1147), .A(n901), .S(n951), .Y(B[37]) );
  MUX2X1 U1102 ( .B(n1149), .A(n1045), .S(n949), .Y(n1147) );
  MUX2X1 U1103 ( .B(n1101), .A(n1150), .S(SH[3]), .Y(n1045) );
  MUX2X1 U1104 ( .B(n1151), .A(n1126), .S(n945), .Y(n1101) );
  MUX2X1 U1105 ( .B(n1140), .A(n1152), .S(n943), .Y(n1126) );
  MUX2X1 U1106 ( .B(A[36]), .A(A[37]), .S(n937), .Y(n1140) );
  MUX2X1 U1107 ( .B(n1153), .A(n935), .S(n950), .Y(B[36]) );
  MUX2X1 U1108 ( .B(n1155), .A(n1052), .S(n949), .Y(n1153) );
  MUX2X1 U1109 ( .B(n1107), .A(n1156), .S(SH[3]), .Y(n1052) );
  MUX2X1 U1110 ( .B(n1157), .A(n1132), .S(n945), .Y(n1107) );
  MUX2X1 U1111 ( .B(n1146), .A(n1158), .S(n942), .Y(n1132) );
  MUX2X1 U1112 ( .B(A[35]), .A(A[36]), .S(n937), .Y(n1146) );
  MUX2X1 U1113 ( .B(n1159), .A(n912), .S(n951), .Y(B[35]) );
  MUX2X1 U1114 ( .B(n1161), .A(n1059), .S(n949), .Y(n1159) );
  MUX2X1 U1115 ( .B(n1113), .A(n1162), .S(SH[3]), .Y(n1059) );
  MUX2X1 U1116 ( .B(n1163), .A(n1139), .S(n945), .Y(n1113) );
  MUX2X1 U1117 ( .B(n1152), .A(n1164), .S(n942), .Y(n1139) );
  MUX2X1 U1118 ( .B(A[34]), .A(A[35]), .S(n936), .Y(n1152) );
  MUX2X1 U1119 ( .B(n1165), .A(n902), .S(n950), .Y(B[34]) );
  MUX2X1 U1120 ( .B(n1167), .A(n1066), .S(n949), .Y(n1165) );
  MUX2X1 U1121 ( .B(n1119), .A(n1168), .S(SH[3]), .Y(n1066) );
  MUX2X1 U1122 ( .B(n1169), .A(n1145), .S(n945), .Y(n1119) );
  MUX2X1 U1123 ( .B(n1158), .A(n1170), .S(n942), .Y(n1145) );
  MUX2X1 U1124 ( .B(A[33]), .A(A[34]), .S(n936), .Y(n1158) );
  MUX2X1 U1125 ( .B(n1171), .A(n897), .S(n951), .Y(B[33]) );
  MUX2X1 U1126 ( .B(n1173), .A(n1074), .S(n949), .Y(n1171) );
  MUX2X1 U1127 ( .B(n1125), .A(n1174), .S(SH[3]), .Y(n1074) );
  MUX2X1 U1128 ( .B(n1175), .A(n1151), .S(n945), .Y(n1125) );
  MUX2X1 U1129 ( .B(n1164), .A(n1176), .S(n942), .Y(n1151) );
  MUX2X1 U1130 ( .B(A[32]), .A(A[33]), .S(n937), .Y(n1164) );
  MUX2X1 U1131 ( .B(n1177), .A(n898), .S(n950), .Y(B[32]) );
  MUX2X1 U1132 ( .B(n1179), .A(n1081), .S(n949), .Y(n1177) );
  MUX2X1 U1133 ( .B(n1131), .A(n1180), .S(SH[3]), .Y(n1081) );
  MUX2X1 U1134 ( .B(n1181), .A(n1157), .S(n945), .Y(n1131) );
  MUX2X1 U1135 ( .B(n1170), .A(n1182), .S(n942), .Y(n1157) );
  MUX2X1 U1136 ( .B(A[31]), .A(A[32]), .S(n937), .Y(n1170) );
  MUX2X1 U1137 ( .B(n1183), .A(n1088), .S(n949), .Y(n959) );
  MUX2X1 U1138 ( .B(n1138), .A(n1184), .S(SH[3]), .Y(n1088) );
  MUX2X1 U1139 ( .B(n1185), .A(n1163), .S(n945), .Y(n1138) );
  MUX2X1 U1140 ( .B(n1176), .A(n1186), .S(n942), .Y(n1163) );
  MUX2X1 U1141 ( .B(A[30]), .A(A[31]), .S(n937), .Y(n1176) );
  MUX2X1 U1142 ( .B(n1187), .A(n1094), .S(n949), .Y(n969) );
  MUX2X1 U1143 ( .B(n1144), .A(n1188), .S(n948), .Y(n1094) );
  MUX2X1 U1144 ( .B(n1189), .A(n1169), .S(n945), .Y(n1144) );
  MUX2X1 U1145 ( .B(n1182), .A(n1190), .S(n942), .Y(n1169) );
  MUX2X1 U1146 ( .B(A[29]), .A(A[30]), .S(n936), .Y(n1182) );
  MUX2X1 U1147 ( .B(n1192), .A(n1100), .S(n949), .Y(n979) );
  MUX2X1 U1148 ( .B(n1150), .A(n1193), .S(n948), .Y(n1100) );
  MUX2X1 U1149 ( .B(n1194), .A(n1175), .S(n945), .Y(n1150) );
  MUX2X1 U1150 ( .B(n1186), .A(n1195), .S(n942), .Y(n1175) );
  MUX2X1 U1151 ( .B(A[28]), .A(A[29]), .S(n936), .Y(n1186) );
  MUX2X1 U1152 ( .B(n1196), .A(n1106), .S(n949), .Y(n988) );
  MUX2X1 U1153 ( .B(n1156), .A(n1197), .S(n948), .Y(n1106) );
  MUX2X1 U1154 ( .B(n1198), .A(n1181), .S(n945), .Y(n1156) );
  MUX2X1 U1155 ( .B(n1190), .A(n1199), .S(n942), .Y(n1181) );
  MUX2X1 U1156 ( .B(A[27]), .A(A[28]), .S(n937), .Y(n1190) );
  MUX2X1 U1157 ( .B(n1200), .A(n1112), .S(n949), .Y(n998) );
  MUX2X1 U1158 ( .B(n1162), .A(n1201), .S(n948), .Y(n1112) );
  MUX2X1 U1159 ( .B(n1202), .A(n1185), .S(n944), .Y(n1162) );
  MUX2X1 U1160 ( .B(n1195), .A(n1203), .S(n942), .Y(n1185) );
  MUX2X1 U1161 ( .B(A[26]), .A(A[27]), .S(n937), .Y(n1195) );
  MUX2X1 U1162 ( .B(n1204), .A(n1118), .S(n949), .Y(n1006) );
  MUX2X1 U1163 ( .B(n1168), .A(n1205), .S(n948), .Y(n1118) );
  MUX2X1 U1164 ( .B(n1206), .A(n1189), .S(n944), .Y(n1168) );
  MUX2X1 U1165 ( .B(n1199), .A(n1207), .S(n942), .Y(n1189) );
  MUX2X1 U1166 ( .B(A[25]), .A(A[26]), .S(n936), .Y(n1199) );
  MUX2X1 U1167 ( .B(n1123), .A(n1124), .S(n949), .Y(n1014) );
  MUX2X1 U1168 ( .B(n1174), .A(n1208), .S(n948), .Y(n1124) );
  MUX2X1 U1169 ( .B(n1209), .A(n1194), .S(n944), .Y(n1174) );
  MUX2X1 U1170 ( .B(n1203), .A(n1210), .S(n941), .Y(n1194) );
  MUX2X1 U1171 ( .B(A[24]), .A(A[25]), .S(n936), .Y(n1203) );
  MUX2X1 U1172 ( .B(n1211), .A(n915), .S(n948), .Y(n1123) );
  MUX2X1 U1173 ( .B(n1129), .A(n1130), .S(n949), .Y(n1022) );
  MUX2X1 U1174 ( .B(n1180), .A(n1213), .S(n948), .Y(n1130) );
  MUX2X1 U1175 ( .B(n1214), .A(n1198), .S(n944), .Y(n1180) );
  MUX2X1 U1176 ( .B(n1207), .A(n1215), .S(n941), .Y(n1198) );
  MUX2X1 U1177 ( .B(A[23]), .A(A[24]), .S(n937), .Y(n1207) );
  MUX2X1 U1178 ( .B(n1216), .A(n919), .S(n948), .Y(n1129) );
  MUX2X1 U1179 ( .B(n932), .A(n1137), .S(n949), .Y(n1030) );
  MUX2X1 U1180 ( .B(n1184), .A(n1218), .S(n948), .Y(n1137) );
  MUX2X1 U1181 ( .B(n1219), .A(n1202), .S(n945), .Y(n1184) );
  MUX2X1 U1182 ( .B(n1210), .A(n1220), .S(n941), .Y(n1202) );
  MUX2X1 U1183 ( .B(A[22]), .A(A[23]), .S(n937), .Y(n1210) );
  MUX2X1 U1184 ( .B(n918), .A(n1143), .S(n949), .Y(n1037) );
  MUX2X1 U1185 ( .B(n1188), .A(n1222), .S(n948), .Y(n1143) );
  MUX2X1 U1186 ( .B(n1223), .A(n1206), .S(n945), .Y(n1188) );
  MUX2X1 U1187 ( .B(n1215), .A(n1224), .S(n941), .Y(n1206) );
  MUX2X1 U1188 ( .B(A[21]), .A(A[22]), .S(n936), .Y(n1215) );
  MUX2X1 U1189 ( .B(n907), .A(n1149), .S(n949), .Y(n1044) );
  MUX2X1 U1190 ( .B(n1193), .A(n1226), .S(n947), .Y(n1149) );
  MUX2X1 U1191 ( .B(n1227), .A(n1209), .S(n945), .Y(n1193) );
  MUX2X1 U1192 ( .B(n1220), .A(n1228), .S(n941), .Y(n1209) );
  MUX2X1 U1193 ( .B(A[20]), .A(A[21]), .S(n936), .Y(n1220) );
  MUX2X1 U1194 ( .B(n905), .A(n1155), .S(n949), .Y(n1051) );
  MUX2X1 U1195 ( .B(n1197), .A(n1230), .S(n947), .Y(n1155) );
  MUX2X1 U1196 ( .B(n1231), .A(n1214), .S(n945), .Y(n1197) );
  MUX2X1 U1197 ( .B(n1224), .A(n1232), .S(n941), .Y(n1214) );
  MUX2X1 U1198 ( .B(A[19]), .A(A[20]), .S(n937), .Y(n1224) );
  MUX2X1 U1199 ( .B(n923), .A(n1161), .S(n949), .Y(n1058) );
  MUX2X1 U1200 ( .B(n1201), .A(n1235), .S(n947), .Y(n1161) );
  MUX2X1 U1201 ( .B(n1236), .A(n1219), .S(n945), .Y(n1201) );
  MUX2X1 U1202 ( .B(n1228), .A(n1237), .S(n941), .Y(n1219) );
  MUX2X1 U1203 ( .B(A[18]), .A(A[19]), .S(n937), .Y(n1228) );
  MUX2X1 U1204 ( .B(n909), .A(n1167), .S(n949), .Y(n1065) );
  MUX2X1 U1205 ( .B(n1205), .A(n1239), .S(n947), .Y(n1167) );
  MUX2X1 U1206 ( .B(n1240), .A(n1223), .S(n945), .Y(n1205) );
  MUX2X1 U1207 ( .B(n1232), .A(n1241), .S(n941), .Y(n1223) );
  MUX2X1 U1208 ( .B(A[17]), .A(A[18]), .S(n936), .Y(n1232) );
  MUX2X1 U1209 ( .B(n911), .A(n1173), .S(n949), .Y(n1073) );
  MUX2X1 U1210 ( .B(n1208), .A(n1211), .S(n947), .Y(n1173) );
  MUX2X1 U1211 ( .B(n1243), .A(n1244), .S(n945), .Y(n1211) );
  MUX2X1 U1212 ( .B(n1245), .A(n1227), .S(n945), .Y(n1208) );
  MUX2X1 U1213 ( .B(n1237), .A(n1246), .S(n941), .Y(n1227) );
  MUX2X1 U1214 ( .B(A[16]), .A(A[17]), .S(n937), .Y(n1237) );
  MUX2X1 U1215 ( .B(n914), .A(n1179), .S(n949), .Y(n1080) );
  MUX2X1 U1216 ( .B(n1213), .A(n1216), .S(n947), .Y(n1179) );
  MUX2X1 U1217 ( .B(n1249), .A(n1250), .S(n945), .Y(n1216) );
  MUX2X1 U1218 ( .B(n1251), .A(n1231), .S(n945), .Y(n1213) );
  MUX2X1 U1219 ( .B(n1241), .A(n1252), .S(n941), .Y(n1231) );
  MUX2X1 U1220 ( .B(A[15]), .A(A[16]), .S(n937), .Y(n1241) );
  MUX2X1 U1221 ( .B(n1218), .A(n1221), .S(n947), .Y(n1183) );
  MUX2X1 U1222 ( .B(n1253), .A(n1254), .S(n944), .Y(n1221) );
  MUX2X1 U1223 ( .B(n1255), .A(n1236), .S(n944), .Y(n1218) );
  MUX2X1 U1224 ( .B(n1246), .A(n1256), .S(n941), .Y(n1236) );
  MUX2X1 U1225 ( .B(A[14]), .A(A[15]), .S(n937), .Y(n1246) );
  MUX2X1 U1226 ( .B(n1222), .A(n1225), .S(n947), .Y(n1187) );
  MUX2X1 U1227 ( .B(n1257), .A(n1258), .S(n944), .Y(n1225) );
  MUX2X1 U1228 ( .B(n1259), .A(n1240), .S(n944), .Y(n1222) );
  MUX2X1 U1229 ( .B(n1252), .A(n1260), .S(n942), .Y(n1240) );
  MUX2X1 U1230 ( .B(A[13]), .A(A[14]), .S(n937), .Y(n1252) );
  MUX2X1 U1231 ( .B(n1226), .A(n1229), .S(n947), .Y(n1192) );
  MUX2X1 U1232 ( .B(n931), .A(n1243), .S(n944), .Y(n1229) );
  MUX2X1 U1233 ( .B(n1261), .A(n1262), .S(n941), .Y(n1243) );
  MUX2X1 U1234 ( .B(n1244), .A(n1245), .S(n944), .Y(n1226) );
  MUX2X1 U1235 ( .B(n1256), .A(n1264), .S(n940), .Y(n1245) );
  MUX2X1 U1236 ( .B(A[12]), .A(A[13]), .S(n937), .Y(n1256) );
  MUX2X1 U1237 ( .B(n1265), .A(n1266), .S(n940), .Y(n1244) );
  MUX2X1 U1238 ( .B(n1230), .A(n1233), .S(n947), .Y(n1196) );
  MUX2X1 U1239 ( .B(n922), .A(n1249), .S(n945), .Y(n1233) );
  MUX2X1 U1240 ( .B(n1268), .A(n1269), .S(n940), .Y(n1249) );
  MUX2X1 U1241 ( .B(n1250), .A(n1251), .S(n944), .Y(n1230) );
  MUX2X1 U1242 ( .B(n1260), .A(n1270), .S(n940), .Y(n1251) );
  MUX2X1 U1243 ( .B(A[11]), .A(A[12]), .S(n937), .Y(n1260) );
  MUX2X1 U1244 ( .B(n1271), .A(n1272), .S(n940), .Y(n1250) );
  MUX2X1 U1245 ( .B(n1235), .A(n934), .S(n947), .Y(n1200) );
  MUX2X1 U1246 ( .B(n1262), .A(n1263), .S(n940), .Y(n1253) );
  MUX2X1 U1247 ( .B(A[0]), .A(A[1]), .S(n937), .Y(n1263) );
  MUX2X1 U1248 ( .B(A[2]), .A(A[3]), .S(n937), .Y(n1262) );
  MUX2X1 U1249 ( .B(n1254), .A(n1255), .S(n945), .Y(n1235) );
  MUX2X1 U1250 ( .B(n1264), .A(n1265), .S(n940), .Y(n1255) );
  MUX2X1 U1251 ( .B(A[8]), .A(A[9]), .S(n937), .Y(n1265) );
  MUX2X1 U1252 ( .B(A[10]), .A(A[11]), .S(n937), .Y(n1264) );
  MUX2X1 U1253 ( .B(n1266), .A(n1261), .S(n940), .Y(n1254) );
  MUX2X1 U1254 ( .B(A[4]), .A(A[5]), .S(n937), .Y(n1261) );
  MUX2X1 U1255 ( .B(A[6]), .A(A[7]), .S(n937), .Y(n1266) );
  MUX2X1 U1256 ( .B(n1239), .A(n924), .S(n947), .Y(n1204) );
  MUX2X1 U1257 ( .B(n1269), .A(n933), .S(n940), .Y(n1257) );
  MUX2X1 U1258 ( .B(A[1]), .A(A[2]), .S(n937), .Y(n1269) );
  MUX2X1 U1259 ( .B(n1258), .A(n1259), .S(n945), .Y(n1239) );
  MUX2X1 U1260 ( .B(n1270), .A(n1271), .S(n940), .Y(n1259) );
  MUX2X1 U1261 ( .B(A[7]), .A(A[8]), .S(n937), .Y(n1271) );
  MUX2X1 U1262 ( .B(A[9]), .A(A[10]), .S(n936), .Y(n1270) );
  MUX2X1 U1263 ( .B(n1272), .A(n1268), .S(n940), .Y(n1258) );
  MUX2X1 U1264 ( .B(A[3]), .A(A[4]), .S(n936), .Y(n1268) );
  MUX2X1 U1265 ( .B(A[5]), .A(A[6]), .S(n936), .Y(n1272) );
endmodule


module alu_DW_leftsh_16 ( A, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  wire   n574, n573, n572, n571, n570, n569, n568, n567, n566, n565, n564,
         n563, n388, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562;

  AND2X1 U338 ( .A(n394), .B(n405), .Y(n490) );
  AND2X1 U339 ( .A(n390), .B(n405), .Y(n497) );
  OR2X1 U340 ( .A(n409), .B(n431), .Y(n565) );
  INVX1 U341 ( .A(n565), .Y(B[9]) );
  OR2X1 U342 ( .A(n409), .B(n432), .Y(n566) );
  INVX1 U343 ( .A(n566), .Y(B[8]) );
  OR2X1 U344 ( .A(n433), .B(SH[4]), .Y(n567) );
  INVX1 U345 ( .A(n567), .Y(B[7]) );
  OR2X1 U346 ( .A(n435), .B(n409), .Y(n569) );
  INVX1 U347 ( .A(n569), .Y(B[5]) );
  OR2X1 U348 ( .A(n436), .B(SH[4]), .Y(n570) );
  INVX1 U349 ( .A(n570), .Y(B[4]) );
  OR2X1 U350 ( .A(n392), .B(n409), .Y(n571) );
  INVX1 U351 ( .A(n571), .Y(B[3]) );
  OR2X1 U352 ( .A(n388), .B(n409), .Y(n572) );
  INVX1 U353 ( .A(n572), .Y(B[2]) );
  OR2X1 U354 ( .A(n409), .B(n473), .Y(n563) );
  INVX1 U355 ( .A(n563), .Y(B[11]) );
  OR2X1 U356 ( .A(n409), .B(n479), .Y(n564) );
  INVX1 U357 ( .A(n564), .Y(B[10]) );
  OR2X1 U358 ( .A(n409), .B(n391), .Y(n574) );
  INVX1 U359 ( .A(n574), .Y(B[0]) );
  OR2X1 U360 ( .A(n409), .B(n395), .Y(n573) );
  INVX1 U361 ( .A(n573), .Y(B[1]) );
  AND2X1 U362 ( .A(n529), .B(n408), .Y(n456) );
  INVX1 U363 ( .A(n456), .Y(n388) );
  OR2X1 U364 ( .A(n434), .B(n409), .Y(n568) );
  INVX1 U365 ( .A(n568), .Y(B[6]) );
  OR2X1 U366 ( .A(n393), .B(n401), .Y(n556) );
  INVX1 U367 ( .A(n556), .Y(n390) );
  AND2X1 U368 ( .A(n497), .B(n408), .Y(n536) );
  INVX1 U369 ( .A(n536), .Y(n391) );
  AND2X1 U370 ( .A(n524), .B(n408), .Y(n437) );
  INVX1 U371 ( .A(n437), .Y(n392) );
  AND2X1 U372 ( .A(A[0]), .B(n399), .Y(n562) );
  INVX1 U373 ( .A(n562), .Y(n393) );
  OR2X1 U374 ( .A(n550), .B(n401), .Y(n535) );
  INVX1 U375 ( .A(n535), .Y(n394) );
  AND2X1 U376 ( .A(n490), .B(n408), .Y(n519) );
  INVX1 U377 ( .A(n519), .Y(n395) );
  INVX1 U378 ( .A(n491), .Y(n427) );
  INVX1 U379 ( .A(n521), .Y(n428) );
  INVX1 U380 ( .A(n498), .Y(n429) );
  INVX1 U381 ( .A(n457), .Y(B[29]) );
  INVX1 U382 ( .A(n465), .Y(B[28]) );
  INVX1 U383 ( .A(n525), .Y(n424) );
  INVX1 U384 ( .A(n530), .Y(n425) );
  INVX1 U385 ( .A(n499), .Y(n419) );
  INVX1 U386 ( .A(n526), .Y(n430) );
  INVX1 U387 ( .A(n474), .Y(n415) );
  INVX1 U388 ( .A(n480), .Y(n416) );
  INVX1 U389 ( .A(n485), .Y(n417) );
  INVX1 U390 ( .A(n492), .Y(n418) );
  INVX1 U391 ( .A(n520), .Y(n423) );
  INVX1 U392 ( .A(n537), .Y(n426) );
  INVX1 U393 ( .A(n504), .Y(n420) );
  INVX1 U394 ( .A(n509), .Y(n421) );
  INVX1 U395 ( .A(n514), .Y(n422) );
  INVX1 U396 ( .A(n447), .Y(B[30]) );
  INVX1 U397 ( .A(n408), .Y(n407) );
  INVX1 U398 ( .A(n405), .Y(n403) );
  INVX1 U399 ( .A(n405), .Y(n404) );
  INVX1 U400 ( .A(n408), .Y(n406) );
  INVX1 U401 ( .A(n438), .Y(B[31]) );
  INVX1 U402 ( .A(n402), .Y(n401) );
  INVX1 U403 ( .A(n402), .Y(n400) );
  INVX1 U404 ( .A(n399), .Y(n398) );
  INVX1 U405 ( .A(n410), .Y(n409) );
  INVX1 U406 ( .A(n399), .Y(n396) );
  INVX1 U407 ( .A(n399), .Y(n397) );
  INVX1 U408 ( .A(SH[0]), .Y(n399) );
  INVX1 U409 ( .A(SH[2]), .Y(n405) );
  INVX1 U410 ( .A(SH[1]), .Y(n402) );
  INVX1 U411 ( .A(SH[3]), .Y(n408) );
  INVX1 U412 ( .A(SH[4]), .Y(n410) );
  MUX2X1 U413 ( .B(n439), .A(n440), .S(n410), .Y(n438) );
  MUX2X1 U414 ( .B(n441), .A(n442), .S(n406), .Y(n440) );
  MUX2X1 U415 ( .B(n443), .A(n444), .S(n403), .Y(n441) );
  MUX2X1 U416 ( .B(n445), .A(n446), .S(n400), .Y(n443) );
  MUX2X1 U417 ( .B(A[31]), .A(A[30]), .S(n396), .Y(n445) );
  MUX2X1 U418 ( .B(n448), .A(n449), .S(n410), .Y(n447) );
  MUX2X1 U419 ( .B(n450), .A(n451), .S(n407), .Y(n449) );
  MUX2X1 U420 ( .B(n452), .A(n453), .S(n403), .Y(n450) );
  MUX2X1 U421 ( .B(n454), .A(n455), .S(n400), .Y(n452) );
  MUX2X1 U422 ( .B(A[30]), .A(A[29]), .S(n396), .Y(n454) );
  MUX2X1 U423 ( .B(n458), .A(n459), .S(n410), .Y(n457) );
  MUX2X1 U424 ( .B(n460), .A(n461), .S(n407), .Y(n459) );
  MUX2X1 U425 ( .B(n462), .A(n463), .S(n403), .Y(n460) );
  MUX2X1 U426 ( .B(n446), .A(n464), .S(n400), .Y(n462) );
  MUX2X1 U427 ( .B(A[29]), .A(A[28]), .S(n396), .Y(n446) );
  MUX2X1 U428 ( .B(n466), .A(n467), .S(n410), .Y(n465) );
  MUX2X1 U429 ( .B(n468), .A(n469), .S(n407), .Y(n467) );
  MUX2X1 U430 ( .B(n470), .A(n471), .S(n403), .Y(n468) );
  MUX2X1 U431 ( .B(n455), .A(n472), .S(n401), .Y(n470) );
  MUX2X1 U432 ( .B(A[28]), .A(A[27]), .S(n396), .Y(n455) );
  MUX2X1 U433 ( .B(n473), .A(n415), .S(n410), .Y(B[27]) );
  MUX2X1 U434 ( .B(n475), .A(n476), .S(n407), .Y(n474) );
  MUX2X1 U435 ( .B(n444), .A(n477), .S(n403), .Y(n475) );
  MUX2X1 U436 ( .B(n464), .A(n478), .S(n401), .Y(n444) );
  MUX2X1 U437 ( .B(A[27]), .A(A[26]), .S(n396), .Y(n464) );
  MUX2X1 U438 ( .B(n479), .A(n416), .S(n410), .Y(B[26]) );
  MUX2X1 U439 ( .B(n481), .A(n482), .S(n407), .Y(n480) );
  MUX2X1 U440 ( .B(n453), .A(n483), .S(n403), .Y(n481) );
  MUX2X1 U441 ( .B(n472), .A(n484), .S(n401), .Y(n453) );
  MUX2X1 U442 ( .B(A[26]), .A(A[25]), .S(n396), .Y(n472) );
  MUX2X1 U443 ( .B(n431), .A(n417), .S(n410), .Y(B[25]) );
  MUX2X1 U444 ( .B(n486), .A(n487), .S(n407), .Y(n485) );
  MUX2X1 U445 ( .B(n463), .A(n488), .S(n403), .Y(n486) );
  MUX2X1 U446 ( .B(n478), .A(n489), .S(n401), .Y(n463) );
  MUX2X1 U447 ( .B(A[25]), .A(A[24]), .S(n396), .Y(n478) );
  MUX2X1 U448 ( .B(n427), .A(n490), .S(n407), .Y(n431) );
  MUX2X1 U449 ( .B(n432), .A(n418), .S(n410), .Y(B[24]) );
  MUX2X1 U450 ( .B(n493), .A(n494), .S(n407), .Y(n492) );
  MUX2X1 U451 ( .B(n471), .A(n495), .S(n403), .Y(n493) );
  MUX2X1 U452 ( .B(n484), .A(n496), .S(n401), .Y(n471) );
  MUX2X1 U453 ( .B(A[24]), .A(A[23]), .S(n396), .Y(n484) );
  MUX2X1 U454 ( .B(n429), .A(n497), .S(n407), .Y(n432) );
  MUX2X1 U455 ( .B(n433), .A(n419), .S(n410), .Y(B[23]) );
  MUX2X1 U456 ( .B(n442), .A(n500), .S(n407), .Y(n499) );
  MUX2X1 U457 ( .B(n477), .A(n501), .S(n403), .Y(n442) );
  MUX2X1 U458 ( .B(n489), .A(n502), .S(n401), .Y(n477) );
  MUX2X1 U459 ( .B(A[23]), .A(A[22]), .S(n396), .Y(n489) );
  OR2X1 U460 ( .A(n503), .B(n406), .Y(n433) );
  MUX2X1 U461 ( .B(n434), .A(n420), .S(n410), .Y(B[22]) );
  MUX2X1 U462 ( .B(n451), .A(n505), .S(n406), .Y(n504) );
  MUX2X1 U463 ( .B(n506), .A(n483), .S(n405), .Y(n451) );
  MUX2X1 U464 ( .B(n496), .A(n507), .S(n401), .Y(n483) );
  MUX2X1 U465 ( .B(A[22]), .A(A[21]), .S(n396), .Y(n496) );
  OR2X1 U466 ( .A(n508), .B(n407), .Y(n434) );
  MUX2X1 U467 ( .B(n435), .A(n421), .S(n410), .Y(B[21]) );
  MUX2X1 U468 ( .B(n461), .A(n510), .S(n406), .Y(n509) );
  MUX2X1 U469 ( .B(n488), .A(n511), .S(n403), .Y(n461) );
  MUX2X1 U470 ( .B(n502), .A(n512), .S(n401), .Y(n488) );
  MUX2X1 U471 ( .B(A[21]), .A(A[20]), .S(n396), .Y(n502) );
  OR2X1 U472 ( .A(n513), .B(n407), .Y(n435) );
  MUX2X1 U473 ( .B(n436), .A(n422), .S(n410), .Y(B[20]) );
  MUX2X1 U474 ( .B(n469), .A(n515), .S(n406), .Y(n514) );
  MUX2X1 U475 ( .B(n495), .A(n516), .S(n403), .Y(n469) );
  MUX2X1 U476 ( .B(n507), .A(n517), .S(n401), .Y(n495) );
  MUX2X1 U477 ( .B(A[20]), .A(A[19]), .S(n396), .Y(n507) );
  OR2X1 U478 ( .A(n518), .B(n406), .Y(n436) );
  MUX2X1 U479 ( .B(n392), .A(n423), .S(n410), .Y(B[19]) );
  MUX2X1 U480 ( .B(n476), .A(n521), .S(n406), .Y(n520) );
  MUX2X1 U481 ( .B(n501), .A(n522), .S(n403), .Y(n476) );
  MUX2X1 U482 ( .B(n523), .A(n512), .S(n402), .Y(n501) );
  MUX2X1 U483 ( .B(A[19]), .A(A[18]), .S(n397), .Y(n512) );
  MUX2X1 U484 ( .B(n388), .A(n424), .S(n410), .Y(B[18]) );
  MUX2X1 U485 ( .B(n482), .A(n526), .S(n406), .Y(n525) );
  MUX2X1 U486 ( .B(n506), .A(n527), .S(n404), .Y(n482) );
  MUX2X1 U487 ( .B(n528), .A(n517), .S(n402), .Y(n506) );
  MUX2X1 U488 ( .B(A[18]), .A(A[17]), .S(n397), .Y(n517) );
  MUX2X1 U489 ( .B(n395), .A(n425), .S(n410), .Y(B[17]) );
  MUX2X1 U490 ( .B(n487), .A(n491), .S(n406), .Y(n530) );
  MUX2X1 U491 ( .B(n531), .A(n532), .S(n404), .Y(n491) );
  MUX2X1 U492 ( .B(n511), .A(n533), .S(n404), .Y(n487) );
  MUX2X1 U493 ( .B(n534), .A(n523), .S(n402), .Y(n511) );
  MUX2X1 U494 ( .B(A[17]), .A(A[16]), .S(n397), .Y(n523) );
  MUX2X1 U495 ( .B(n391), .A(n426), .S(n410), .Y(B[16]) );
  MUX2X1 U496 ( .B(n494), .A(n498), .S(n406), .Y(n537) );
  MUX2X1 U497 ( .B(n538), .A(n539), .S(n404), .Y(n498) );
  MUX2X1 U498 ( .B(n516), .A(n540), .S(n404), .Y(n494) );
  MUX2X1 U499 ( .B(n541), .A(n528), .S(n402), .Y(n516) );
  MUX2X1 U500 ( .B(A[16]), .A(A[15]), .S(n397), .Y(n528) );
  AND2X1 U501 ( .A(n439), .B(n410), .Y(B[15]) );
  MUX2X1 U502 ( .B(n503), .A(n500), .S(n408), .Y(n439) );
  MUX2X1 U503 ( .B(n522), .A(n542), .S(n404), .Y(n500) );
  MUX2X1 U504 ( .B(n543), .A(n534), .S(n402), .Y(n522) );
  MUX2X1 U505 ( .B(A[15]), .A(A[14]), .S(n397), .Y(n534) );
  MUX2X1 U506 ( .B(n544), .A(n545), .S(n404), .Y(n503) );
  AND2X1 U507 ( .A(n410), .B(n448), .Y(B[14]) );
  MUX2X1 U508 ( .B(n505), .A(n508), .S(n406), .Y(n448) );
  MUX2X1 U509 ( .B(n546), .A(n547), .S(n404), .Y(n508) );
  MUX2X1 U510 ( .B(n527), .A(n548), .S(n404), .Y(n505) );
  MUX2X1 U511 ( .B(n549), .A(n541), .S(n402), .Y(n527) );
  MUX2X1 U512 ( .B(A[14]), .A(A[13]), .S(n397), .Y(n541) );
  AND2X1 U513 ( .A(n458), .B(n410), .Y(B[13]) );
  MUX2X1 U514 ( .B(n510), .A(n513), .S(n406), .Y(n458) );
  MUX2X1 U515 ( .B(n532), .A(n394), .S(n404), .Y(n513) );
  MUX2X1 U516 ( .B(n551), .A(n552), .S(n402), .Y(n532) );
  MUX2X1 U517 ( .B(n533), .A(n531), .S(n404), .Y(n510) );
  MUX2X1 U518 ( .B(n553), .A(n554), .S(n402), .Y(n531) );
  MUX2X1 U519 ( .B(n555), .A(n543), .S(n402), .Y(n533) );
  MUX2X1 U520 ( .B(A[13]), .A(A[12]), .S(n397), .Y(n543) );
  AND2X1 U521 ( .A(n466), .B(n410), .Y(B[12]) );
  MUX2X1 U522 ( .B(n515), .A(n518), .S(n406), .Y(n466) );
  MUX2X1 U523 ( .B(n539), .A(n390), .S(n404), .Y(n518) );
  MUX2X1 U524 ( .B(n557), .A(n558), .S(n402), .Y(n539) );
  MUX2X1 U525 ( .B(n540), .A(n538), .S(n403), .Y(n515) );
  MUX2X1 U526 ( .B(n559), .A(n560), .S(n402), .Y(n538) );
  MUX2X1 U527 ( .B(n561), .A(n549), .S(n402), .Y(n540) );
  MUX2X1 U528 ( .B(A[12]), .A(A[11]), .S(n397), .Y(n549) );
  MUX2X1 U529 ( .B(n428), .A(n524), .S(n406), .Y(n473) );
  AND2X1 U530 ( .A(n545), .B(n405), .Y(n524) );
  MUX2X1 U531 ( .B(n550), .A(n551), .S(n402), .Y(n545) );
  MUX2X1 U532 ( .B(A[3]), .A(A[2]), .S(n397), .Y(n551) );
  MUX2X1 U533 ( .B(A[1]), .A(A[0]), .S(n397), .Y(n550) );
  MUX2X1 U534 ( .B(n542), .A(n544), .S(n403), .Y(n521) );
  MUX2X1 U535 ( .B(n552), .A(n553), .S(n402), .Y(n544) );
  MUX2X1 U536 ( .B(A[7]), .A(A[6]), .S(n397), .Y(n553) );
  MUX2X1 U537 ( .B(A[5]), .A(A[4]), .S(n397), .Y(n552) );
  MUX2X1 U538 ( .B(n554), .A(n555), .S(n402), .Y(n542) );
  MUX2X1 U539 ( .B(A[11]), .A(A[10]), .S(n398), .Y(n555) );
  MUX2X1 U540 ( .B(A[9]), .A(A[8]), .S(n398), .Y(n554) );
  MUX2X1 U541 ( .B(n430), .A(n529), .S(n407), .Y(n479) );
  AND2X1 U542 ( .A(n547), .B(n405), .Y(n529) );
  MUX2X1 U543 ( .B(n393), .A(n557), .S(n402), .Y(n547) );
  MUX2X1 U544 ( .B(A[2]), .A(A[1]), .S(n398), .Y(n557) );
  MUX2X1 U545 ( .B(n548), .A(n546), .S(n403), .Y(n526) );
  MUX2X1 U546 ( .B(n558), .A(n559), .S(n402), .Y(n546) );
  MUX2X1 U547 ( .B(A[6]), .A(A[5]), .S(n398), .Y(n559) );
  MUX2X1 U548 ( .B(A[4]), .A(A[3]), .S(n398), .Y(n558) );
  MUX2X1 U549 ( .B(n560), .A(n561), .S(n402), .Y(n548) );
  MUX2X1 U550 ( .B(A[10]), .A(A[9]), .S(n398), .Y(n561) );
  MUX2X1 U551 ( .B(A[8]), .A(A[7]), .S(n398), .Y(n560) );
endmodule


module alu_DW_leftsh_17 ( A, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  wire   n573, n572, n571, n570, n569, n568, n567, n566, n565, n564, n563,
         n562, n388, n389, n390, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561;

  AND2X1 U338 ( .A(n394), .B(n404), .Y(n489) );
  AND2X1 U339 ( .A(n389), .B(n404), .Y(n496) );
  OR2X1 U340 ( .A(n408), .B(n430), .Y(n564) );
  INVX1 U341 ( .A(n564), .Y(B[9]) );
  OR2X1 U342 ( .A(n408), .B(n431), .Y(n565) );
  INVX1 U343 ( .A(n565), .Y(B[8]) );
  OR2X1 U344 ( .A(n432), .B(n408), .Y(n566) );
  INVX1 U345 ( .A(n566), .Y(B[7]) );
  OR2X1 U346 ( .A(n434), .B(n408), .Y(n568) );
  INVX1 U347 ( .A(n568), .Y(B[5]) );
  OR2X1 U348 ( .A(n435), .B(n408), .Y(n569) );
  INVX1 U349 ( .A(n569), .Y(B[4]) );
  OR2X1 U350 ( .A(n392), .B(n408), .Y(n570) );
  INVX1 U351 ( .A(n570), .Y(B[3]) );
  OR2X1 U352 ( .A(n408), .B(n472), .Y(n562) );
  INVX1 U353 ( .A(n562), .Y(B[11]) );
  OR2X1 U354 ( .A(n408), .B(n478), .Y(n563) );
  INVX1 U355 ( .A(n563), .Y(B[10]) );
  OR2X1 U356 ( .A(n408), .B(n390), .Y(n573) );
  INVX1 U357 ( .A(n573), .Y(B[0]) );
  OR2X1 U358 ( .A(n408), .B(n395), .Y(n572) );
  INVX1 U359 ( .A(n572), .Y(B[1]) );
  OR2X1 U360 ( .A(n388), .B(n408), .Y(n571) );
  INVX1 U361 ( .A(n571), .Y(B[2]) );
  AND2X1 U362 ( .A(n528), .B(n407), .Y(n455) );
  INVX1 U363 ( .A(n455), .Y(n388) );
  OR2X1 U364 ( .A(n393), .B(n401), .Y(n555) );
  INVX1 U365 ( .A(n555), .Y(n389) );
  AND2X1 U366 ( .A(n496), .B(n407), .Y(n535) );
  INVX1 U367 ( .A(n535), .Y(n390) );
  OR2X1 U368 ( .A(n433), .B(n408), .Y(n567) );
  INVX1 U369 ( .A(n567), .Y(B[6]) );
  AND2X1 U370 ( .A(n523), .B(n407), .Y(n436) );
  INVX1 U371 ( .A(n436), .Y(n392) );
  AND2X1 U372 ( .A(A[0]), .B(n399), .Y(n561) );
  INVX1 U373 ( .A(n561), .Y(n393) );
  OR2X1 U374 ( .A(n549), .B(n401), .Y(n534) );
  INVX1 U375 ( .A(n534), .Y(n394) );
  AND2X1 U376 ( .A(n489), .B(n407), .Y(n518) );
  INVX1 U377 ( .A(n518), .Y(n395) );
  INVX1 U378 ( .A(n490), .Y(n426) );
  INVX1 U379 ( .A(n520), .Y(n427) );
  INVX1 U380 ( .A(n525), .Y(n429) );
  INVX1 U381 ( .A(n497), .Y(n428) );
  INVX1 U382 ( .A(n536), .Y(n425) );
  INVX1 U383 ( .A(n407), .Y(n406) );
  INVX1 U384 ( .A(n407), .Y(n405) );
  INVX1 U385 ( .A(n404), .Y(n403) );
  INVX1 U386 ( .A(n519), .Y(n422) );
  INVX1 U387 ( .A(n524), .Y(n423) );
  INVX1 U388 ( .A(n529), .Y(n424) );
  INVX1 U389 ( .A(n503), .Y(n419) );
  INVX1 U390 ( .A(n508), .Y(n420) );
  INVX1 U391 ( .A(n513), .Y(n421) );
  INVX1 U392 ( .A(n498), .Y(n418) );
  INVX1 U393 ( .A(n464), .Y(B[28]) );
  INVX1 U394 ( .A(n402), .Y(n400) );
  INVX1 U395 ( .A(n437), .Y(B[31]) );
  INVX1 U396 ( .A(SH[3]), .Y(n407) );
  INVX1 U397 ( .A(n402), .Y(n401) );
  INVX1 U398 ( .A(SH[2]), .Y(n404) );
  INVX1 U399 ( .A(n473), .Y(n414) );
  INVX1 U400 ( .A(n479), .Y(n415) );
  INVX1 U401 ( .A(n484), .Y(n416) );
  INVX1 U402 ( .A(n491), .Y(n417) );
  INVX1 U403 ( .A(n456), .Y(B[29]) );
  INVX1 U404 ( .A(n409), .Y(n408) );
  INVX1 U405 ( .A(SH[1]), .Y(n402) );
  INVX1 U406 ( .A(n399), .Y(n398) );
  INVX1 U407 ( .A(SH[4]), .Y(n409) );
  INVX1 U408 ( .A(n446), .Y(B[30]) );
  INVX1 U409 ( .A(n399), .Y(n396) );
  INVX1 U410 ( .A(n399), .Y(n397) );
  INVX1 U411 ( .A(SH[0]), .Y(n399) );
  MUX2X1 U412 ( .B(n438), .A(n439), .S(n409), .Y(n437) );
  MUX2X1 U413 ( .B(n440), .A(n441), .S(n405), .Y(n439) );
  MUX2X1 U414 ( .B(n442), .A(n443), .S(n403), .Y(n440) );
  MUX2X1 U415 ( .B(n444), .A(n445), .S(n400), .Y(n442) );
  MUX2X1 U416 ( .B(A[31]), .A(A[30]), .S(n396), .Y(n444) );
  MUX2X1 U417 ( .B(n447), .A(n448), .S(n409), .Y(n446) );
  MUX2X1 U418 ( .B(n449), .A(n450), .S(n406), .Y(n448) );
  MUX2X1 U419 ( .B(n451), .A(n452), .S(n403), .Y(n449) );
  MUX2X1 U420 ( .B(n453), .A(n454), .S(n400), .Y(n451) );
  MUX2X1 U421 ( .B(A[30]), .A(A[29]), .S(n396), .Y(n453) );
  MUX2X1 U422 ( .B(n457), .A(n458), .S(n409), .Y(n456) );
  MUX2X1 U423 ( .B(n459), .A(n460), .S(n406), .Y(n458) );
  MUX2X1 U424 ( .B(n461), .A(n462), .S(n403), .Y(n459) );
  MUX2X1 U425 ( .B(n445), .A(n463), .S(n400), .Y(n461) );
  MUX2X1 U426 ( .B(A[29]), .A(A[28]), .S(n396), .Y(n445) );
  MUX2X1 U427 ( .B(n465), .A(n466), .S(n409), .Y(n464) );
  MUX2X1 U428 ( .B(n467), .A(n468), .S(n406), .Y(n466) );
  MUX2X1 U429 ( .B(n469), .A(n470), .S(n403), .Y(n467) );
  MUX2X1 U430 ( .B(n454), .A(n471), .S(n401), .Y(n469) );
  MUX2X1 U431 ( .B(A[28]), .A(A[27]), .S(n396), .Y(n454) );
  MUX2X1 U432 ( .B(n472), .A(n414), .S(n409), .Y(B[27]) );
  MUX2X1 U433 ( .B(n474), .A(n475), .S(n406), .Y(n473) );
  MUX2X1 U434 ( .B(n443), .A(n476), .S(n403), .Y(n474) );
  MUX2X1 U435 ( .B(n463), .A(n477), .S(n401), .Y(n443) );
  MUX2X1 U436 ( .B(A[27]), .A(A[26]), .S(n396), .Y(n463) );
  MUX2X1 U437 ( .B(n478), .A(n415), .S(n409), .Y(B[26]) );
  MUX2X1 U438 ( .B(n480), .A(n481), .S(n406), .Y(n479) );
  MUX2X1 U439 ( .B(n452), .A(n482), .S(n403), .Y(n480) );
  MUX2X1 U440 ( .B(n471), .A(n483), .S(n401), .Y(n452) );
  MUX2X1 U441 ( .B(A[26]), .A(A[25]), .S(n396), .Y(n471) );
  MUX2X1 U442 ( .B(n430), .A(n416), .S(n409), .Y(B[25]) );
  MUX2X1 U443 ( .B(n485), .A(n486), .S(n406), .Y(n484) );
  MUX2X1 U444 ( .B(n462), .A(n487), .S(n403), .Y(n485) );
  MUX2X1 U445 ( .B(n477), .A(n488), .S(n401), .Y(n462) );
  MUX2X1 U446 ( .B(A[25]), .A(A[24]), .S(n396), .Y(n477) );
  MUX2X1 U447 ( .B(n426), .A(n489), .S(n406), .Y(n430) );
  MUX2X1 U448 ( .B(n431), .A(n417), .S(n409), .Y(B[24]) );
  MUX2X1 U449 ( .B(n492), .A(n493), .S(n406), .Y(n491) );
  MUX2X1 U450 ( .B(n470), .A(n494), .S(n403), .Y(n492) );
  MUX2X1 U451 ( .B(n483), .A(n495), .S(n401), .Y(n470) );
  MUX2X1 U452 ( .B(A[24]), .A(A[23]), .S(n396), .Y(n483) );
  MUX2X1 U453 ( .B(n428), .A(n496), .S(n406), .Y(n431) );
  MUX2X1 U454 ( .B(n432), .A(n418), .S(n409), .Y(B[23]) );
  MUX2X1 U455 ( .B(n441), .A(n499), .S(n406), .Y(n498) );
  MUX2X1 U456 ( .B(n476), .A(n500), .S(n403), .Y(n441) );
  MUX2X1 U457 ( .B(n488), .A(n501), .S(n401), .Y(n476) );
  MUX2X1 U458 ( .B(A[23]), .A(A[22]), .S(n396), .Y(n488) );
  OR2X1 U459 ( .A(n502), .B(n406), .Y(n432) );
  MUX2X1 U460 ( .B(n433), .A(n419), .S(n409), .Y(B[22]) );
  MUX2X1 U461 ( .B(n450), .A(n504), .S(n405), .Y(n503) );
  MUX2X1 U462 ( .B(n505), .A(n482), .S(n404), .Y(n450) );
  MUX2X1 U463 ( .B(n495), .A(n506), .S(n401), .Y(n482) );
  MUX2X1 U464 ( .B(A[22]), .A(A[21]), .S(n396), .Y(n495) );
  OR2X1 U465 ( .A(n507), .B(n406), .Y(n433) );
  MUX2X1 U466 ( .B(n434), .A(n420), .S(n409), .Y(B[21]) );
  MUX2X1 U467 ( .B(n460), .A(n509), .S(n405), .Y(n508) );
  MUX2X1 U468 ( .B(n487), .A(n510), .S(n403), .Y(n460) );
  MUX2X1 U469 ( .B(n501), .A(n511), .S(n401), .Y(n487) );
  MUX2X1 U470 ( .B(A[21]), .A(A[20]), .S(n396), .Y(n501) );
  OR2X1 U471 ( .A(n512), .B(n406), .Y(n434) );
  MUX2X1 U472 ( .B(n435), .A(n421), .S(n409), .Y(B[20]) );
  MUX2X1 U473 ( .B(n468), .A(n514), .S(n405), .Y(n513) );
  MUX2X1 U474 ( .B(n494), .A(n515), .S(n403), .Y(n468) );
  MUX2X1 U475 ( .B(n506), .A(n516), .S(n401), .Y(n494) );
  MUX2X1 U476 ( .B(A[20]), .A(A[19]), .S(n396), .Y(n506) );
  OR2X1 U477 ( .A(n517), .B(n406), .Y(n435) );
  MUX2X1 U478 ( .B(n392), .A(n422), .S(n409), .Y(B[19]) );
  MUX2X1 U479 ( .B(n475), .A(n520), .S(n405), .Y(n519) );
  MUX2X1 U480 ( .B(n500), .A(n521), .S(n403), .Y(n475) );
  MUX2X1 U481 ( .B(n522), .A(n511), .S(n402), .Y(n500) );
  MUX2X1 U482 ( .B(A[19]), .A(A[18]), .S(n397), .Y(n511) );
  MUX2X1 U483 ( .B(n388), .A(n423), .S(n409), .Y(B[18]) );
  MUX2X1 U484 ( .B(n481), .A(n525), .S(n405), .Y(n524) );
  MUX2X1 U485 ( .B(n505), .A(n526), .S(SH[2]), .Y(n481) );
  MUX2X1 U486 ( .B(n527), .A(n516), .S(n402), .Y(n505) );
  MUX2X1 U487 ( .B(A[18]), .A(A[17]), .S(n397), .Y(n516) );
  MUX2X1 U488 ( .B(n395), .A(n424), .S(n409), .Y(B[17]) );
  MUX2X1 U489 ( .B(n486), .A(n490), .S(n405), .Y(n529) );
  MUX2X1 U490 ( .B(n530), .A(n531), .S(SH[2]), .Y(n490) );
  MUX2X1 U491 ( .B(n510), .A(n532), .S(SH[2]), .Y(n486) );
  MUX2X1 U492 ( .B(n533), .A(n522), .S(n402), .Y(n510) );
  MUX2X1 U493 ( .B(A[17]), .A(A[16]), .S(n397), .Y(n522) );
  MUX2X1 U494 ( .B(n390), .A(n425), .S(n409), .Y(B[16]) );
  MUX2X1 U495 ( .B(n493), .A(n497), .S(n405), .Y(n536) );
  MUX2X1 U496 ( .B(n537), .A(n538), .S(SH[2]), .Y(n497) );
  MUX2X1 U497 ( .B(n515), .A(n539), .S(SH[2]), .Y(n493) );
  MUX2X1 U498 ( .B(n540), .A(n527), .S(n402), .Y(n515) );
  MUX2X1 U499 ( .B(A[16]), .A(A[15]), .S(n397), .Y(n527) );
  AND2X1 U500 ( .A(n438), .B(n409), .Y(B[15]) );
  MUX2X1 U501 ( .B(n502), .A(n499), .S(n407), .Y(n438) );
  MUX2X1 U502 ( .B(n521), .A(n541), .S(SH[2]), .Y(n499) );
  MUX2X1 U503 ( .B(n542), .A(n533), .S(n402), .Y(n521) );
  MUX2X1 U504 ( .B(A[15]), .A(A[14]), .S(n397), .Y(n533) );
  MUX2X1 U505 ( .B(n543), .A(n544), .S(SH[2]), .Y(n502) );
  AND2X1 U506 ( .A(n409), .B(n447), .Y(B[14]) );
  MUX2X1 U507 ( .B(n504), .A(n507), .S(n405), .Y(n447) );
  MUX2X1 U508 ( .B(n545), .A(n546), .S(SH[2]), .Y(n507) );
  MUX2X1 U509 ( .B(n526), .A(n547), .S(SH[2]), .Y(n504) );
  MUX2X1 U510 ( .B(n548), .A(n540), .S(n402), .Y(n526) );
  MUX2X1 U511 ( .B(A[14]), .A(A[13]), .S(n397), .Y(n540) );
  AND2X1 U512 ( .A(n457), .B(n409), .Y(B[13]) );
  MUX2X1 U513 ( .B(n509), .A(n512), .S(n405), .Y(n457) );
  MUX2X1 U514 ( .B(n531), .A(n394), .S(SH[2]), .Y(n512) );
  MUX2X1 U515 ( .B(n550), .A(n551), .S(n402), .Y(n531) );
  MUX2X1 U516 ( .B(n532), .A(n530), .S(SH[2]), .Y(n509) );
  MUX2X1 U517 ( .B(n552), .A(n553), .S(n402), .Y(n530) );
  MUX2X1 U518 ( .B(n554), .A(n542), .S(n402), .Y(n532) );
  MUX2X1 U519 ( .B(A[13]), .A(A[12]), .S(n397), .Y(n542) );
  AND2X1 U520 ( .A(n465), .B(n409), .Y(B[12]) );
  MUX2X1 U521 ( .B(n514), .A(n517), .S(n405), .Y(n465) );
  MUX2X1 U522 ( .B(n538), .A(n389), .S(SH[2]), .Y(n517) );
  MUX2X1 U523 ( .B(n556), .A(n557), .S(n402), .Y(n538) );
  MUX2X1 U524 ( .B(n539), .A(n537), .S(SH[2]), .Y(n514) );
  MUX2X1 U525 ( .B(n558), .A(n559), .S(n402), .Y(n537) );
  MUX2X1 U526 ( .B(n560), .A(n548), .S(n402), .Y(n539) );
  MUX2X1 U527 ( .B(A[12]), .A(A[11]), .S(n397), .Y(n548) );
  MUX2X1 U528 ( .B(n427), .A(n523), .S(n405), .Y(n472) );
  AND2X1 U529 ( .A(n544), .B(n404), .Y(n523) );
  MUX2X1 U530 ( .B(n549), .A(n550), .S(n402), .Y(n544) );
  MUX2X1 U531 ( .B(A[3]), .A(A[2]), .S(n397), .Y(n550) );
  MUX2X1 U532 ( .B(A[1]), .A(A[0]), .S(n397), .Y(n549) );
  MUX2X1 U533 ( .B(n541), .A(n543), .S(SH[2]), .Y(n520) );
  MUX2X1 U534 ( .B(n551), .A(n552), .S(n402), .Y(n543) );
  MUX2X1 U535 ( .B(A[7]), .A(A[6]), .S(n397), .Y(n552) );
  MUX2X1 U536 ( .B(A[5]), .A(A[4]), .S(n397), .Y(n551) );
  MUX2X1 U537 ( .B(n553), .A(n554), .S(n402), .Y(n541) );
  MUX2X1 U538 ( .B(A[11]), .A(A[10]), .S(n398), .Y(n554) );
  MUX2X1 U539 ( .B(A[9]), .A(A[8]), .S(n398), .Y(n553) );
  MUX2X1 U540 ( .B(n429), .A(n528), .S(n406), .Y(n478) );
  AND2X1 U541 ( .A(n546), .B(n404), .Y(n528) );
  MUX2X1 U542 ( .B(n393), .A(n556), .S(n402), .Y(n546) );
  MUX2X1 U543 ( .B(A[2]), .A(A[1]), .S(n398), .Y(n556) );
  MUX2X1 U544 ( .B(n547), .A(n545), .S(n403), .Y(n525) );
  MUX2X1 U545 ( .B(n557), .A(n558), .S(n402), .Y(n545) );
  MUX2X1 U546 ( .B(A[6]), .A(A[5]), .S(n398), .Y(n558) );
  MUX2X1 U547 ( .B(A[4]), .A(A[3]), .S(n398), .Y(n557) );
  MUX2X1 U548 ( .B(n559), .A(n560), .S(n402), .Y(n547) );
  MUX2X1 U549 ( .B(A[10]), .A(A[9]), .S(n398), .Y(n560) );
  MUX2X1 U550 ( .B(A[8]), .A(A[7]), .S(n398), .Y(n559) );
endmodule


module alu_DW01_sub_7 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [7:2] carry;

  FAX1 U2_7 ( .A(A[7]), .B(n8), .C(carry[7]), .YC(), .YS(DIFF[7]) );
  FAX1 U2_6 ( .A(A[6]), .B(n7), .C(carry[6]), .YC(carry[7]), .YS(DIFF[6]) );
  FAX1 U2_5 ( .A(A[5]), .B(n6), .C(carry[5]), .YC(carry[6]), .YS(DIFF[5]) );
  FAX1 U2_4 ( .A(A[4]), .B(n5), .C(carry[4]), .YC(carry[5]), .YS(DIFF[4]) );
  FAX1 U2_3 ( .A(A[3]), .B(n4), .C(carry[3]), .YC(carry[4]), .YS(DIFF[3]) );
  FAX1 U2_2 ( .A(A[2]), .B(n3), .C(carry[2]), .YC(carry[3]), .YS(DIFF[2]) );
  FAX1 U2_1 ( .A(A[1]), .B(n2), .C(n9), .YC(carry[2]), .YS(DIFF[1]) );
  OR2X1 U1 ( .A(A[0]), .B(n1), .Y(n9) );
  INVX1 U2 ( .A(B[1]), .Y(n2) );
  INVX1 U3 ( .A(B[4]), .Y(n5) );
  INVX1 U4 ( .A(B[3]), .Y(n4) );
  INVX1 U5 ( .A(B[0]), .Y(n1) );
  INVX1 U6 ( .A(B[6]), .Y(n7) );
  INVX1 U7 ( .A(B[2]), .Y(n3) );
  INVX1 U8 ( .A(B[7]), .Y(n8) );
  INVX1 U9 ( .A(B[5]), .Y(n6) );
  XNOR2X1 U10 ( .A(n1), .B(A[0]), .Y(DIFF[0]) );
endmodule


module alu_DW01_sub_8 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [7:2] carry;

  FAX1 U2_7 ( .A(A[7]), .B(n8), .C(carry[7]), .YC(), .YS(DIFF[7]) );
  FAX1 U2_6 ( .A(A[6]), .B(n7), .C(carry[6]), .YC(carry[7]), .YS(DIFF[6]) );
  FAX1 U2_5 ( .A(A[5]), .B(n6), .C(carry[5]), .YC(carry[6]), .YS(DIFF[5]) );
  FAX1 U2_4 ( .A(A[4]), .B(n5), .C(carry[4]), .YC(carry[5]), .YS(DIFF[4]) );
  FAX1 U2_3 ( .A(A[3]), .B(n4), .C(carry[3]), .YC(carry[4]), .YS(DIFF[3]) );
  FAX1 U2_2 ( .A(A[2]), .B(n3), .C(carry[2]), .YC(carry[3]), .YS(DIFF[2]) );
  FAX1 U2_1 ( .A(A[1]), .B(n2), .C(n9), .YC(carry[2]), .YS(DIFF[1]) );
  OR2X1 U1 ( .A(A[0]), .B(n1), .Y(n9) );
  INVX1 U2 ( .A(B[1]), .Y(n2) );
  INVX1 U3 ( .A(B[6]), .Y(n7) );
  INVX1 U4 ( .A(B[3]), .Y(n4) );
  INVX1 U5 ( .A(B[5]), .Y(n6) );
  INVX1 U6 ( .A(B[4]), .Y(n5) );
  INVX1 U7 ( .A(B[7]), .Y(n8) );
  INVX1 U8 ( .A(B[2]), .Y(n3) );
  INVX1 U9 ( .A(B[0]), .Y(n1) );
  XNOR2X1 U10 ( .A(n1), .B(A[0]), .Y(DIFF[0]) );
endmodule


module alu_DW01_sub_9 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [7:2] carry;

  FAX1 U2_7 ( .A(A[7]), .B(n9), .C(carry[7]), .YC(), .YS(DIFF[7]) );
  FAX1 U2_6 ( .A(A[6]), .B(n8), .C(carry[6]), .YC(carry[7]), .YS(DIFF[6]) );
  FAX1 U2_5 ( .A(A[5]), .B(n7), .C(carry[5]), .YC(carry[6]), .YS(DIFF[5]) );
  FAX1 U2_4 ( .A(A[4]), .B(n6), .C(carry[4]), .YC(carry[5]), .YS(DIFF[4]) );
  FAX1 U2_3 ( .A(A[3]), .B(n5), .C(carry[3]), .YC(carry[4]), .YS(DIFF[3]) );
  FAX1 U2_2 ( .A(A[2]), .B(n4), .C(carry[2]), .YC(carry[3]), .YS(DIFF[2]) );
  FAX1 U2_1 ( .A(A[1]), .B(n3), .C(n1), .YC(carry[2]), .YS(DIFF[1]) );
  INVX1 U1 ( .A(B[3]), .Y(n5) );
  INVX1 U2 ( .A(B[2]), .Y(n4) );
  OR2X1 U3 ( .A(A[0]), .B(n2), .Y(n1) );
  INVX1 U4 ( .A(B[0]), .Y(n2) );
  INVX1 U5 ( .A(B[5]), .Y(n7) );
  INVX1 U6 ( .A(B[6]), .Y(n8) );
  INVX1 U7 ( .A(B[7]), .Y(n9) );
  INVX1 U8 ( .A(B[1]), .Y(n3) );
  INVX1 U9 ( .A(B[4]), .Y(n6) );
  XNOR2X1 U10 ( .A(n2), .B(A[0]), .Y(DIFF[0]) );
endmodule


module alu_DW01_sub_10 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [7:2] carry;

  FAX1 U2_7 ( .A(A[7]), .B(n8), .C(carry[7]), .YC(), .YS(DIFF[7]) );
  FAX1 U2_6 ( .A(A[6]), .B(n7), .C(carry[6]), .YC(carry[7]), .YS(DIFF[6]) );
  FAX1 U2_5 ( .A(A[5]), .B(n6), .C(carry[5]), .YC(carry[6]), .YS(DIFF[5]) );
  FAX1 U2_4 ( .A(A[4]), .B(n5), .C(carry[4]), .YC(carry[5]), .YS(DIFF[4]) );
  FAX1 U2_3 ( .A(A[3]), .B(n4), .C(carry[3]), .YC(carry[4]), .YS(DIFF[3]) );
  FAX1 U2_2 ( .A(A[2]), .B(n3), .C(carry[2]), .YC(carry[3]), .YS(DIFF[2]) );
  FAX1 U2_1 ( .A(A[1]), .B(n2), .C(n9), .YC(carry[2]), .YS(DIFF[1]) );
  OR2X1 U1 ( .A(A[0]), .B(n1), .Y(n9) );
  INVX1 U2 ( .A(B[1]), .Y(n2) );
  INVX1 U3 ( .A(B[2]), .Y(n3) );
  INVX1 U4 ( .A(B[0]), .Y(n1) );
  INVX1 U5 ( .A(B[5]), .Y(n6) );
  INVX1 U6 ( .A(B[6]), .Y(n7) );
  INVX1 U7 ( .A(B[3]), .Y(n4) );
  INVX1 U8 ( .A(B[4]), .Y(n5) );
  INVX1 U9 ( .A(B[7]), .Y(n8) );
  XNOR2X1 U10 ( .A(n1), .B(A[0]), .Y(DIFF[0]) );
endmodule


module alu_DW01_sub_11 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [7:2] carry;

  FAX1 U2_7 ( .A(A[7]), .B(n8), .C(carry[7]), .YC(), .YS(DIFF[7]) );
  FAX1 U2_6 ( .A(A[6]), .B(n7), .C(carry[6]), .YC(carry[7]), .YS(DIFF[6]) );
  FAX1 U2_5 ( .A(A[5]), .B(n6), .C(carry[5]), .YC(carry[6]), .YS(DIFF[5]) );
  FAX1 U2_4 ( .A(A[4]), .B(n5), .C(carry[4]), .YC(carry[5]), .YS(DIFF[4]) );
  FAX1 U2_3 ( .A(A[3]), .B(n4), .C(carry[3]), .YC(carry[4]), .YS(DIFF[3]) );
  FAX1 U2_2 ( .A(A[2]), .B(n3), .C(carry[2]), .YC(carry[3]), .YS(DIFF[2]) );
  FAX1 U2_1 ( .A(A[1]), .B(n2), .C(n9), .YC(carry[2]), .YS(DIFF[1]) );
  OR2X1 U1 ( .A(A[0]), .B(n1), .Y(n9) );
  INVX1 U2 ( .A(B[2]), .Y(n3) );
  INVX1 U3 ( .A(B[1]), .Y(n2) );
  INVX1 U4 ( .A(B[4]), .Y(n5) );
  INVX1 U5 ( .A(B[3]), .Y(n4) );
  INVX1 U6 ( .A(B[6]), .Y(n7) );
  INVX1 U7 ( .A(B[5]), .Y(n6) );
  INVX1 U8 ( .A(B[0]), .Y(n1) );
  INVX1 U9 ( .A(B[7]), .Y(n8) );
  XNOR2X1 U10 ( .A(n1), .B(A[0]), .Y(DIFF[0]) );
endmodule


module alu_DW01_sub_12 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [7:2] carry;

  FAX1 U2_7 ( .A(A[7]), .B(n8), .C(carry[7]), .YC(), .YS(DIFF[7]) );
  FAX1 U2_6 ( .A(A[6]), .B(n7), .C(carry[6]), .YC(carry[7]), .YS(DIFF[6]) );
  FAX1 U2_5 ( .A(A[5]), .B(n6), .C(carry[5]), .YC(carry[6]), .YS(DIFF[5]) );
  FAX1 U2_4 ( .A(A[4]), .B(n5), .C(carry[4]), .YC(carry[5]), .YS(DIFF[4]) );
  FAX1 U2_3 ( .A(A[3]), .B(n4), .C(carry[3]), .YC(carry[4]), .YS(DIFF[3]) );
  FAX1 U2_2 ( .A(A[2]), .B(n3), .C(carry[2]), .YC(carry[3]), .YS(DIFF[2]) );
  FAX1 U2_1 ( .A(A[1]), .B(n2), .C(n9), .YC(carry[2]), .YS(DIFF[1]) );
  OR2X1 U1 ( .A(A[0]), .B(n1), .Y(n9) );
  INVX1 U2 ( .A(B[2]), .Y(n3) );
  INVX1 U3 ( .A(B[1]), .Y(n2) );
  INVX1 U4 ( .A(B[6]), .Y(n7) );
  INVX1 U5 ( .A(B[0]), .Y(n1) );
  INVX1 U6 ( .A(B[4]), .Y(n5) );
  INVX1 U7 ( .A(B[3]), .Y(n4) );
  INVX1 U8 ( .A(B[5]), .Y(n6) );
  INVX1 U9 ( .A(B[7]), .Y(n8) );
  XNOR2X1 U10 ( .A(n1), .B(A[0]), .Y(DIFF[0]) );
endmodule


module alu_DW01_sub_13 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [7:2] carry;

  FAX1 U2_7 ( .A(A[7]), .B(n8), .C(carry[7]), .YC(), .YS(DIFF[7]) );
  FAX1 U2_6 ( .A(A[6]), .B(n7), .C(carry[6]), .YC(carry[7]), .YS(DIFF[6]) );
  FAX1 U2_5 ( .A(A[5]), .B(n6), .C(carry[5]), .YC(carry[6]), .YS(DIFF[5]) );
  FAX1 U2_4 ( .A(A[4]), .B(n5), .C(carry[4]), .YC(carry[5]), .YS(DIFF[4]) );
  FAX1 U2_3 ( .A(A[3]), .B(n4), .C(carry[3]), .YC(carry[4]), .YS(DIFF[3]) );
  FAX1 U2_2 ( .A(A[2]), .B(n3), .C(carry[2]), .YC(carry[3]), .YS(DIFF[2]) );
  FAX1 U2_1 ( .A(A[1]), .B(n2), .C(n9), .YC(carry[2]), .YS(DIFF[1]) );
  OR2X1 U1 ( .A(A[0]), .B(n1), .Y(n9) );
  INVX1 U2 ( .A(B[2]), .Y(n3) );
  INVX1 U3 ( .A(B[3]), .Y(n4) );
  INVX1 U4 ( .A(B[0]), .Y(n1) );
  INVX1 U5 ( .A(B[4]), .Y(n5) );
  INVX1 U6 ( .A(B[5]), .Y(n6) );
  INVX1 U7 ( .A(B[1]), .Y(n2) );
  INVX1 U8 ( .A(B[6]), .Y(n7) );
  INVX1 U9 ( .A(B[7]), .Y(n8) );
  XNOR2X1 U10 ( .A(n1), .B(A[0]), .Y(DIFF[0]) );
endmodule


module alu_DW01_sub_14 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [7:2] carry;

  FAX1 U2_7 ( .A(A[7]), .B(n8), .C(carry[7]), .YC(), .YS(DIFF[7]) );
  FAX1 U2_6 ( .A(A[6]), .B(n7), .C(carry[6]), .YC(carry[7]), .YS(DIFF[6]) );
  FAX1 U2_5 ( .A(A[5]), .B(n6), .C(carry[5]), .YC(carry[6]), .YS(DIFF[5]) );
  FAX1 U2_4 ( .A(A[4]), .B(n5), .C(carry[4]), .YC(carry[5]), .YS(DIFF[4]) );
  FAX1 U2_3 ( .A(A[3]), .B(n4), .C(carry[3]), .YC(carry[4]), .YS(DIFF[3]) );
  FAX1 U2_2 ( .A(A[2]), .B(n3), .C(carry[2]), .YC(carry[3]), .YS(DIFF[2]) );
  FAX1 U2_1 ( .A(A[1]), .B(n2), .C(n9), .YC(carry[2]), .YS(DIFF[1]) );
  OR2X1 U1 ( .A(A[0]), .B(n1), .Y(n9) );
  INVX1 U2 ( .A(B[1]), .Y(n2) );
  INVX1 U3 ( .A(B[2]), .Y(n3) );
  INVX1 U4 ( .A(B[0]), .Y(n1) );
  INVX1 U5 ( .A(B[3]), .Y(n4) );
  INVX1 U6 ( .A(B[5]), .Y(n6) );
  INVX1 U7 ( .A(B[6]), .Y(n7) );
  INVX1 U8 ( .A(B[4]), .Y(n5) );
  INVX1 U9 ( .A(B[7]), .Y(n8) );
  XNOR2X1 U10 ( .A(n1), .B(A[0]), .Y(DIFF[0]) );
endmodule


module alu_DW01_add_7 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:2] carry;

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X1 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module alu_DW01_add_8 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:2] carry;

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X1 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module alu_DW01_add_9 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:2] carry;

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module alu_DW01_add_10 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:2] carry;

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X1 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module alu_DW01_add_11 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:2] carry;

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X1 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module alu_DW01_add_12 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:2] carry;

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X1 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module alu_DW01_add_13 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:2] carry;

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X1 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module alu_DW01_add_14 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:2] carry;

  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X1 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module alu_DW_mult_uns_23 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71;
  assign product[0] = b[0];

  FAX1 U2 ( .A(a[7]), .B(n44), .C(n2), .YC(product[15]), .YS(product[14]) );
  FAX1 U3 ( .A(n45), .B(n14), .C(n3), .YC(n2), .YS(product[13]) );
  FAX1 U4 ( .A(n15), .B(n16), .C(n4), .YC(n3), .YS(product[12]) );
  FAX1 U5 ( .A(n17), .B(n18), .C(n5), .YC(n4), .YS(product[11]) );
  FAX1 U6 ( .A(n22), .B(n19), .C(n6), .YC(n5), .YS(product[10]) );
  FAX1 U7 ( .A(n26), .B(n23), .C(n7), .YC(n6), .YS(product[9]) );
  FAX1 U8 ( .A(n32), .B(n27), .C(n8), .YC(n7), .YS(product[8]) );
  FAX1 U9 ( .A(n36), .B(n33), .C(n9), .YC(n8), .YS(product[7]) );
  FAX1 U10 ( .A(n39), .B(n37), .C(n10), .YC(n9), .YS(product[6]) );
  FAX1 U11 ( .A(n42), .B(n41), .C(n11), .YC(n10), .YS(product[5]) );
  FAX1 U12 ( .A(n68), .B(n43), .C(n12), .YC(n11), .YS(product[4]) );
  HAX1 U13 ( .A(n70), .B(n13), .YC(n12), .YS(product[3]) );
  HAX1 U14 ( .A(a[1]), .B(n71), .YC(n13), .YS(product[2]) );
  FAX1 U15 ( .A(a[6]), .B(n51), .C(n46), .YC(n14), .YS(n15) );
  FAX1 U16 ( .A(n52), .B(n47), .C(n20), .YC(n16), .YS(n17) );
  FAX1 U17 ( .A(n53), .B(n24), .C(n21), .YC(n18), .YS(n19) );
  FAX1 U18 ( .A(a[5]), .B(n57), .C(n48), .YC(n20), .YS(n21) );
  FAX1 U19 ( .A(n30), .B(n28), .C(n25), .YC(n22), .YS(n23) );
  FAX1 U20 ( .A(n58), .B(n49), .C(n54), .YC(n24), .YS(n25) );
  FAX1 U21 ( .A(n34), .B(n31), .C(n29), .YC(n26), .YS(n27) );
  FAX1 U22 ( .A(n62), .B(n50), .C(n59), .YC(n28), .YS(n29) );
  HAX1 U23 ( .A(a[4]), .B(n55), .YC(n30), .YS(n31) );
  FAX1 U24 ( .A(n60), .B(n38), .C(n35), .YC(n32), .YS(n33) );
  HAX1 U25 ( .A(n63), .B(n56), .YC(n34), .YS(n35) );
  FAX1 U26 ( .A(n64), .B(n61), .C(n40), .YC(n36), .YS(n37) );
  HAX1 U27 ( .A(a[3]), .B(n66), .YC(n38), .YS(n39) );
  HAX1 U28 ( .A(n67), .B(n65), .YC(n40), .YS(n41) );
  HAX1 U29 ( .A(a[2]), .B(n69), .YC(n42), .YS(n43) );
  AND2X1 U75 ( .A(b[3]), .B(b[1]), .Y(n67) );
  AND2X1 U76 ( .A(b[5]), .B(b[2]), .Y(n59) );
  AND2X1 U77 ( .A(b[4]), .B(b[3]), .Y(n62) );
  AND2X1 U78 ( .A(b[6]), .B(b[3]), .Y(n53) );
  AND2X1 U79 ( .A(b[7]), .B(b[5]), .Y(n45) );
  AND2X1 U80 ( .A(b[3]), .B(b[0]), .Y(n68) );
  AND2X1 U81 ( .A(b[1]), .B(b[0]), .Y(n71) );
  AND2X1 U82 ( .A(b[3]), .B(b[2]), .Y(n66) );
  AND2X1 U83 ( .A(b[5]), .B(b[0]), .Y(n61) );
  AND2X2 U84 ( .A(b[6]), .B(b[5]), .Y(n51) );
  AND2X2 U85 ( .A(b[5]), .B(b[4]), .Y(n57) );
  AND2X2 U86 ( .A(b[5]), .B(b[1]), .Y(n60) );
  AND2X2 U87 ( .A(b[2]), .B(b[1]), .Y(n69) );
  AND2X2 U88 ( .A(b[7]), .B(b[3]), .Y(n47) );
  AND2X2 U89 ( .A(b[5]), .B(b[3]), .Y(n58) );
  AND2X1 U90 ( .A(b[4]), .B(b[0]), .Y(n65) );
  AND2X1 U91 ( .A(b[2]), .B(b[0]), .Y(n70) );
  AND2X1 U92 ( .A(b[7]), .B(b[0]), .Y(n50) );
  AND2X1 U93 ( .A(b[6]), .B(b[2]), .Y(n54) );
  AND2X1 U94 ( .A(b[7]), .B(b[2]), .Y(n48) );
  AND2X1 U95 ( .A(b[4]), .B(b[2]), .Y(n63) );
  AND2X1 U96 ( .A(b[6]), .B(b[0]), .Y(n56) );
  AND2X1 U97 ( .A(b[4]), .B(b[1]), .Y(n64) );
  AND2X1 U98 ( .A(b[6]), .B(b[1]), .Y(n55) );
  AND2X1 U99 ( .A(b[6]), .B(b[4]), .Y(n52) );
  AND2X1 U100 ( .A(b[7]), .B(b[1]), .Y(n49) );
  AND2X1 U101 ( .A(b[7]), .B(b[4]), .Y(n46) );
  AND2X1 U102 ( .A(b[7]), .B(b[6]), .Y(n44) );
endmodule


module alu_DW_mult_uns_22 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161;

  FAX1 U2 ( .A(n99), .B(n15), .C(n2), .YC(product[15]), .YS(product[14]) );
  FAX1 U3 ( .A(n16), .B(n17), .C(n3), .YC(n2), .YS(product[13]) );
  FAX1 U4 ( .A(n18), .B(n21), .C(n4), .YC(n3), .YS(product[12]) );
  FAX1 U5 ( .A(n22), .B(n27), .C(n5), .YC(n4), .YS(product[11]) );
  FAX1 U6 ( .A(n35), .B(n28), .C(n6), .YC(n5), .YS(product[10]) );
  FAX1 U7 ( .A(n45), .B(n36), .C(n7), .YC(n6), .YS(product[9]) );
  FAX1 U8 ( .A(n57), .B(n46), .C(n8), .YC(n7), .YS(product[8]) );
  FAX1 U9 ( .A(n69), .B(n58), .C(n9), .YC(n8), .YS(product[7]) );
  FAX1 U10 ( .A(n79), .B(n70), .C(n10), .YC(n9), .YS(product[6]) );
  FAX1 U11 ( .A(n87), .B(n80), .C(n11), .YC(n10), .YS(product[5]) );
  FAX1 U12 ( .A(n93), .B(n88), .C(n12), .YC(n11), .YS(product[4]) );
  FAX1 U13 ( .A(n96), .B(n94), .C(n13), .YC(n12), .YS(product[3]) );
  FAX1 U14 ( .A(n146), .B(n14), .C(n98), .YC(n13), .YS(product[2]) );
  HAX1 U15 ( .A(n154), .B(n161), .YC(n14), .YS(product[1]) );
  FAX1 U16 ( .A(n107), .B(n100), .C(n19), .YC(n15), .YS(n16) );
  FAX1 U17 ( .A(n25), .B(n20), .C(n23), .YC(n17), .YS(n18) );
  FAX1 U18 ( .A(n115), .B(n101), .C(n108), .YC(n19), .YS(n20) );
  FAX1 U19 ( .A(n31), .B(n24), .C(n29), .YC(n21), .YS(n22) );
  FAX1 U20 ( .A(n116), .B(n33), .C(n26), .YC(n23), .YS(n24) );
  FAX1 U21 ( .A(n123), .B(n102), .C(n109), .YC(n25), .YS(n26) );
  FAX1 U22 ( .A(n39), .B(n37), .C(n30), .YC(n27), .YS(n28) );
  FAX1 U23 ( .A(n41), .B(n34), .C(n32), .YC(n29), .YS(n30) );
  FAX1 U24 ( .A(n124), .B(n117), .C(n43), .YC(n31), .YS(n32) );
  FAX1 U25 ( .A(n131), .B(n103), .C(n110), .YC(n33), .YS(n34) );
  FAX1 U26 ( .A(n40), .B(n47), .C(n38), .YC(n35), .YS(n36) );
  FAX1 U27 ( .A(n44), .B(n51), .C(n49), .YC(n37), .YS(n38) );
  FAX1 U28 ( .A(n55), .B(n53), .C(n42), .YC(n39), .YS(n40) );
  FAX1 U29 ( .A(n118), .B(n125), .C(n132), .YC(n41), .YS(n42) );
  FAX1 U30 ( .A(n139), .B(n104), .C(n111), .YC(n43), .YS(n44) );
  FAX1 U31 ( .A(n50), .B(n59), .C(n48), .YC(n45), .YS(n46) );
  FAX1 U32 ( .A(n54), .B(n52), .C(n61), .YC(n47), .YS(n48) );
  FAX1 U33 ( .A(n56), .B(n65), .C(n63), .YC(n49), .YS(n50) );
  FAX1 U34 ( .A(n140), .B(n133), .C(n67), .YC(n51), .YS(n52) );
  FAX1 U35 ( .A(n126), .B(n119), .C(n147), .YC(n53), .YS(n54) );
  HAX1 U36 ( .A(n112), .B(n105), .YC(n55), .YS(n56) );
  FAX1 U37 ( .A(n62), .B(n71), .C(n60), .YC(n57), .YS(n58) );
  FAX1 U38 ( .A(n64), .B(n66), .C(n73), .YC(n59), .YS(n60) );
  FAX1 U39 ( .A(n77), .B(n68), .C(n75), .YC(n61), .YS(n62) );
  FAX1 U40 ( .A(n141), .B(n127), .C(n134), .YC(n63), .YS(n64) );
  FAX1 U41 ( .A(n155), .B(n120), .C(n148), .YC(n65), .YS(n66) );
  HAX1 U42 ( .A(n113), .B(n106), .YC(n67), .YS(n68) );
  FAX1 U43 ( .A(n74), .B(n81), .C(n72), .YC(n69), .YS(n70) );
  FAX1 U44 ( .A(n78), .B(n83), .C(n76), .YC(n71), .YS(n72) );
  FAX1 U45 ( .A(n142), .B(n135), .C(n85), .YC(n73), .YS(n74) );
  FAX1 U46 ( .A(n156), .B(n128), .C(n149), .YC(n75), .YS(n76) );
  HAX1 U47 ( .A(n121), .B(n114), .YC(n77), .YS(n78) );
  FAX1 U48 ( .A(n89), .B(n84), .C(n82), .YC(n79), .YS(n80) );
  FAX1 U49 ( .A(n150), .B(n91), .C(n86), .YC(n81), .YS(n82) );
  FAX1 U50 ( .A(n157), .B(n136), .C(n143), .YC(n83), .YS(n84) );
  HAX1 U51 ( .A(n129), .B(n122), .YC(n85), .YS(n86) );
  FAX1 U52 ( .A(n95), .B(n92), .C(n90), .YC(n87), .YS(n88) );
  FAX1 U53 ( .A(n158), .B(n144), .C(n151), .YC(n89), .YS(n90) );
  HAX1 U54 ( .A(n137), .B(n130), .YC(n91), .YS(n92) );
  FAX1 U55 ( .A(n159), .B(n152), .C(n97), .YC(n93), .YS(n94) );
  HAX1 U56 ( .A(n145), .B(n138), .YC(n95), .YS(n96) );
  HAX1 U57 ( .A(n160), .B(n153), .YC(n97), .YS(n98) );
  AND2X1 U140 ( .A(a[3]), .B(b[5]), .Y(n133) );
  AND2X1 U141 ( .A(a[4]), .B(b[1]), .Y(n129) );
  AND2X1 U142 ( .A(a[5]), .B(b[4]), .Y(n118) );
  AND2X1 U143 ( .A(a[3]), .B(b[6]), .Y(n132) );
  AND2X1 U144 ( .A(a[5]), .B(b[5]), .Y(n117) );
  AND2X1 U145 ( .A(a[5]), .B(b[6]), .Y(n116) );
  AND2X1 U146 ( .A(a[5]), .B(b[3]), .Y(n119) );
  AND2X1 U147 ( .A(b[1]), .B(a[7]), .Y(n105) );
  AND2X1 U148 ( .A(a[3]), .B(b[4]), .Y(n134) );
  AND2X1 U149 ( .A(a[5]), .B(b[2]), .Y(n120) );
  AND2X1 U150 ( .A(a[6]), .B(b[1]), .Y(n113) );
  AND2X1 U151 ( .A(a[5]), .B(b[7]), .Y(n115) );
  AND2X1 U152 ( .A(a[3]), .B(b[1]), .Y(n137) );
  AND2X1 U153 ( .A(a[5]), .B(b[1]), .Y(n121) );
  AND2X1 U154 ( .A(b[6]), .B(a[0]), .Y(n156) );
  AND2X1 U155 ( .A(a[2]), .B(b[1]), .Y(n145) );
  AND2X1 U156 ( .A(a[3]), .B(b[0]), .Y(n138) );
  AND2X1 U157 ( .A(a[3]), .B(b[2]), .Y(n136) );
  AND2X1 U158 ( .A(a[3]), .B(b[3]), .Y(n135) );
  AND2X1 U159 ( .A(a[1]), .B(b[1]), .Y(n153) );
  AND2X1 U160 ( .A(b[1]), .B(a[0]), .Y(n161) );
  AND2X2 U161 ( .A(a[5]), .B(b[0]), .Y(n122) );
  AND2X2 U162 ( .A(a[3]), .B(b[7]), .Y(n131) );
  AND2X1 U163 ( .A(a[6]), .B(b[2]), .Y(n112) );
  AND2X1 U164 ( .A(a[1]), .B(b[0]), .Y(n154) );
  AND2X1 U165 ( .A(a[4]), .B(b[0]), .Y(n130) );
  AND2X1 U166 ( .A(a[7]), .B(b[0]), .Y(n106) );
  AND2X1 U167 ( .A(b[2]), .B(a[0]), .Y(n160) );
  AND2X1 U168 ( .A(a[2]), .B(b[0]), .Y(n146) );
  AND2X1 U169 ( .A(a[6]), .B(b[0]), .Y(n114) );
  AND2X1 U170 ( .A(b[0]), .B(a[0]), .Y(product[0]) );
  AND2X1 U171 ( .A(b[2]), .B(a[7]), .Y(n104) );
  AND2X1 U172 ( .A(a[1]), .B(b[2]), .Y(n152) );
  AND2X1 U173 ( .A(a[2]), .B(b[2]), .Y(n144) );
  AND2X1 U174 ( .A(a[4]), .B(b[2]), .Y(n128) );
  AND2X1 U175 ( .A(b[7]), .B(a[7]), .Y(n99) );
  AND2X1 U176 ( .A(b[3]), .B(a[0]), .Y(n159) );
  AND2X1 U177 ( .A(b[4]), .B(a[0]), .Y(n158) );
  AND2X1 U178 ( .A(b[5]), .B(a[0]), .Y(n157) );
  AND2X1 U179 ( .A(b[7]), .B(a[0]), .Y(n155) );
  AND2X1 U180 ( .A(a[1]), .B(b[3]), .Y(n151) );
  AND2X1 U181 ( .A(a[1]), .B(b[4]), .Y(n150) );
  AND2X1 U182 ( .A(a[1]), .B(b[5]), .Y(n149) );
  AND2X1 U183 ( .A(a[1]), .B(b[6]), .Y(n148) );
  AND2X1 U184 ( .A(a[1]), .B(b[7]), .Y(n147) );
  AND2X1 U185 ( .A(a[2]), .B(b[3]), .Y(n143) );
  AND2X1 U186 ( .A(a[2]), .B(b[4]), .Y(n142) );
  AND2X1 U187 ( .A(a[2]), .B(b[5]), .Y(n141) );
  AND2X1 U188 ( .A(a[2]), .B(b[6]), .Y(n140) );
  AND2X1 U189 ( .A(a[2]), .B(b[7]), .Y(n139) );
  AND2X1 U190 ( .A(a[4]), .B(b[3]), .Y(n127) );
  AND2X1 U191 ( .A(a[4]), .B(b[4]), .Y(n126) );
  AND2X1 U192 ( .A(a[4]), .B(b[5]), .Y(n125) );
  AND2X1 U193 ( .A(a[4]), .B(b[6]), .Y(n124) );
  AND2X1 U194 ( .A(a[4]), .B(b[7]), .Y(n123) );
  AND2X1 U195 ( .A(a[6]), .B(b[3]), .Y(n111) );
  AND2X1 U196 ( .A(a[6]), .B(b[4]), .Y(n110) );
  AND2X1 U197 ( .A(a[6]), .B(b[5]), .Y(n109) );
  AND2X1 U198 ( .A(a[6]), .B(b[6]), .Y(n108) );
  AND2X1 U199 ( .A(a[6]), .B(b[7]), .Y(n107) );
  AND2X1 U200 ( .A(b[3]), .B(a[7]), .Y(n103) );
  AND2X1 U201 ( .A(b[4]), .B(a[7]), .Y(n102) );
  AND2X1 U202 ( .A(b[5]), .B(a[7]), .Y(n101) );
  AND2X1 U203 ( .A(b[6]), .B(a[7]), .Y(n100) );
endmodule


module alu_DW_mult_uns_19 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71;
  assign product[0] = b[0];

  FAX1 U2 ( .A(a[7]), .B(n44), .C(n2), .YC(product[15]), .YS(product[14]) );
  FAX1 U3 ( .A(n45), .B(n14), .C(n3), .YC(n2), .YS(product[13]) );
  FAX1 U4 ( .A(n15), .B(n16), .C(n4), .YC(n3), .YS(product[12]) );
  FAX1 U5 ( .A(n17), .B(n18), .C(n5), .YC(n4), .YS(product[11]) );
  FAX1 U6 ( .A(n22), .B(n19), .C(n6), .YC(n5), .YS(product[10]) );
  FAX1 U7 ( .A(n26), .B(n23), .C(n7), .YC(n6), .YS(product[9]) );
  FAX1 U8 ( .A(n32), .B(n27), .C(n8), .YC(n7), .YS(product[8]) );
  FAX1 U9 ( .A(n36), .B(n33), .C(n9), .YC(n8), .YS(product[7]) );
  FAX1 U10 ( .A(n39), .B(n37), .C(n10), .YC(n9), .YS(product[6]) );
  FAX1 U11 ( .A(n42), .B(n41), .C(n11), .YC(n10), .YS(product[5]) );
  FAX1 U12 ( .A(n68), .B(n43), .C(n12), .YC(n11), .YS(product[4]) );
  HAX1 U13 ( .A(n70), .B(n13), .YC(n12), .YS(product[3]) );
  HAX1 U14 ( .A(b[1]), .B(n71), .YC(n13), .YS(product[2]) );
  FAX1 U15 ( .A(a[6]), .B(n51), .C(n46), .YC(n14), .YS(n15) );
  FAX1 U16 ( .A(n52), .B(n47), .C(n20), .YC(n16), .YS(n17) );
  FAX1 U17 ( .A(n53), .B(n24), .C(n21), .YC(n18), .YS(n19) );
  FAX1 U18 ( .A(a[5]), .B(n57), .C(n48), .YC(n20), .YS(n21) );
  FAX1 U19 ( .A(n30), .B(n28), .C(n25), .YC(n22), .YS(n23) );
  FAX1 U20 ( .A(n58), .B(n49), .C(n54), .YC(n24), .YS(n25) );
  FAX1 U21 ( .A(n34), .B(n31), .C(n29), .YC(n26), .YS(n27) );
  FAX1 U22 ( .A(n62), .B(n50), .C(n59), .YC(n28), .YS(n29) );
  HAX1 U23 ( .A(a[4]), .B(n55), .YC(n30), .YS(n31) );
  FAX1 U24 ( .A(n60), .B(n38), .C(n35), .YC(n32), .YS(n33) );
  HAX1 U25 ( .A(n63), .B(n56), .YC(n34), .YS(n35) );
  FAX1 U26 ( .A(n64), .B(n61), .C(n40), .YC(n36), .YS(n37) );
  HAX1 U27 ( .A(a[3]), .B(n66), .YC(n38), .YS(n39) );
  HAX1 U28 ( .A(n67), .B(n65), .YC(n40), .YS(n41) );
  HAX1 U29 ( .A(a[2]), .B(n69), .YC(n42), .YS(n43) );
  AND2X2 U75 ( .A(b[5]), .B(b[1]), .Y(n60) );
  AND2X2 U76 ( .A(b[5]), .B(b[2]), .Y(n59) );
  AND2X1 U77 ( .A(b[3]), .B(b[1]), .Y(n67) );
  AND2X1 U78 ( .A(b[4]), .B(b[3]), .Y(n62) );
  AND2X1 U79 ( .A(b[6]), .B(b[3]), .Y(n53) );
  AND2X1 U80 ( .A(b[5]), .B(b[0]), .Y(n61) );
  AND2X1 U81 ( .A(b[7]), .B(b[5]), .Y(n45) );
  AND2X1 U82 ( .A(b[3]), .B(b[0]), .Y(n68) );
  AND2X2 U83 ( .A(b[7]), .B(b[6]), .Y(n44) );
  AND2X2 U84 ( .A(b[6]), .B(b[5]), .Y(n51) );
  AND2X2 U85 ( .A(b[5]), .B(b[4]), .Y(n57) );
  AND2X2 U86 ( .A(b[7]), .B(b[3]), .Y(n47) );
  AND2X2 U87 ( .A(b[5]), .B(b[3]), .Y(n58) );
  AND2X2 U88 ( .A(b[3]), .B(b[2]), .Y(n66) );
  AND2X1 U89 ( .A(b[4]), .B(b[1]), .Y(n64) );
  AND2X1 U90 ( .A(b[6]), .B(b[1]), .Y(n55) );
  AND2X1 U91 ( .A(b[2]), .B(b[1]), .Y(n69) );
  AND2X1 U92 ( .A(b[7]), .B(b[1]), .Y(n49) );
  AND2X1 U93 ( .A(b[1]), .B(b[0]), .Y(n71) );
  AND2X1 U94 ( .A(b[2]), .B(b[0]), .Y(n70) );
  AND2X1 U95 ( .A(b[4]), .B(b[0]), .Y(n65) );
  AND2X1 U96 ( .A(b[4]), .B(b[2]), .Y(n63) );
  AND2X1 U97 ( .A(b[6]), .B(b[0]), .Y(n56) );
  AND2X1 U98 ( .A(b[6]), .B(b[2]), .Y(n54) );
  AND2X1 U99 ( .A(b[6]), .B(b[4]), .Y(n52) );
  AND2X1 U100 ( .A(b[7]), .B(b[0]), .Y(n50) );
  AND2X1 U101 ( .A(b[7]), .B(b[2]), .Y(n48) );
  AND2X1 U102 ( .A(b[7]), .B(b[4]), .Y(n46) );
endmodule


module alu_DW_mult_uns_18 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n214;

  FAX1 U2 ( .A(n99), .B(n15), .C(n2), .YC(product[15]), .YS(product[14]) );
  FAX1 U3 ( .A(n16), .B(n17), .C(n3), .YC(n2), .YS(product[13]) );
  FAX1 U4 ( .A(n18), .B(n21), .C(n4), .YC(n3), .YS(product[12]) );
  FAX1 U5 ( .A(n22), .B(n27), .C(n5), .YC(n4), .YS(product[11]) );
  FAX1 U6 ( .A(n35), .B(n28), .C(n6), .YC(n5), .YS(product[10]) );
  FAX1 U7 ( .A(n45), .B(n36), .C(n7), .YC(n6), .YS(product[9]) );
  FAX1 U8 ( .A(n57), .B(n46), .C(n8), .YC(n7), .YS(product[8]) );
  FAX1 U9 ( .A(n69), .B(n58), .C(n9), .YC(n8), .YS(product[7]) );
  FAX1 U10 ( .A(n79), .B(n70), .C(n10), .YC(n9), .YS(product[6]) );
  FAX1 U11 ( .A(n87), .B(n80), .C(n11), .YC(n10), .YS(product[5]) );
  FAX1 U12 ( .A(n93), .B(n88), .C(n12), .YC(n11), .YS(product[4]) );
  FAX1 U13 ( .A(n96), .B(n94), .C(n13), .YC(n12), .YS(product[3]) );
  FAX1 U14 ( .A(n146), .B(n14), .C(n98), .YC(n13), .YS(product[2]) );
  HAX1 U15 ( .A(n154), .B(n161), .YC(n14), .YS(product[1]) );
  FAX1 U16 ( .A(n107), .B(n100), .C(n19), .YC(n15), .YS(n16) );
  FAX1 U17 ( .A(n25), .B(n20), .C(n23), .YC(n17), .YS(n18) );
  FAX1 U18 ( .A(n115), .B(n101), .C(n108), .YC(n19), .YS(n20) );
  FAX1 U19 ( .A(n31), .B(n24), .C(n29), .YC(n21), .YS(n22) );
  FAX1 U20 ( .A(n116), .B(n33), .C(n26), .YC(n23), .YS(n24) );
  FAX1 U21 ( .A(n123), .B(n102), .C(n109), .YC(n25), .YS(n26) );
  FAX1 U22 ( .A(n39), .B(n37), .C(n30), .YC(n27), .YS(n28) );
  FAX1 U23 ( .A(n41), .B(n34), .C(n32), .YC(n29), .YS(n30) );
  FAX1 U24 ( .A(n124), .B(n117), .C(n43), .YC(n31), .YS(n32) );
  FAX1 U25 ( .A(n131), .B(n103), .C(n110), .YC(n33), .YS(n34) );
  FAX1 U26 ( .A(n40), .B(n47), .C(n38), .YC(n35), .YS(n36) );
  FAX1 U27 ( .A(n44), .B(n51), .C(n49), .YC(n37), .YS(n38) );
  FAX1 U28 ( .A(n55), .B(n53), .C(n42), .YC(n39), .YS(n40) );
  FAX1 U29 ( .A(n118), .B(n125), .C(n132), .YC(n41), .YS(n42) );
  FAX1 U30 ( .A(n139), .B(n104), .C(n111), .YC(n43), .YS(n44) );
  FAX1 U31 ( .A(n50), .B(n59), .C(n48), .YC(n45), .YS(n46) );
  FAX1 U32 ( .A(n54), .B(n52), .C(n61), .YC(n47), .YS(n48) );
  FAX1 U33 ( .A(n56), .B(n65), .C(n63), .YC(n49), .YS(n50) );
  FAX1 U34 ( .A(n140), .B(n133), .C(n67), .YC(n51), .YS(n52) );
  FAX1 U35 ( .A(n126), .B(n119), .C(n147), .YC(n53), .YS(n54) );
  HAX1 U36 ( .A(n112), .B(n105), .YC(n55), .YS(n56) );
  FAX1 U37 ( .A(n62), .B(n71), .C(n60), .YC(n57), .YS(n58) );
  FAX1 U38 ( .A(n64), .B(n66), .C(n73), .YC(n59), .YS(n60) );
  FAX1 U39 ( .A(n77), .B(n68), .C(n75), .YC(n61), .YS(n62) );
  FAX1 U40 ( .A(n141), .B(n127), .C(n134), .YC(n63), .YS(n64) );
  FAX1 U41 ( .A(n155), .B(n120), .C(n148), .YC(n65), .YS(n66) );
  HAX1 U42 ( .A(n113), .B(n106), .YC(n67), .YS(n68) );
  FAX1 U43 ( .A(n74), .B(n81), .C(n72), .YC(n69), .YS(n70) );
  FAX1 U44 ( .A(n78), .B(n83), .C(n76), .YC(n71), .YS(n72) );
  FAX1 U45 ( .A(n142), .B(n135), .C(n85), .YC(n73), .YS(n74) );
  FAX1 U46 ( .A(n156), .B(n128), .C(n149), .YC(n75), .YS(n76) );
  HAX1 U47 ( .A(n121), .B(n114), .YC(n77), .YS(n78) );
  FAX1 U48 ( .A(n89), .B(n84), .C(n82), .YC(n79), .YS(n80) );
  FAX1 U49 ( .A(n150), .B(n91), .C(n86), .YC(n81), .YS(n82) );
  FAX1 U50 ( .A(n157), .B(n136), .C(n143), .YC(n83), .YS(n84) );
  HAX1 U51 ( .A(n129), .B(n122), .YC(n85), .YS(n86) );
  FAX1 U52 ( .A(n95), .B(n92), .C(n90), .YC(n87), .YS(n88) );
  FAX1 U53 ( .A(n158), .B(n144), .C(n151), .YC(n89), .YS(n90) );
  HAX1 U54 ( .A(n137), .B(n130), .YC(n91), .YS(n92) );
  FAX1 U55 ( .A(n159), .B(n152), .C(n97), .YC(n93), .YS(n94) );
  HAX1 U56 ( .A(n145), .B(n138), .YC(n95), .YS(n96) );
  HAX1 U57 ( .A(n160), .B(n153), .YC(n97), .YS(n98) );
  AND2X2 U140 ( .A(b[7]), .B(a[7]), .Y(n99) );
  AND2X2 U141 ( .A(a[4]), .B(b[7]), .Y(n123) );
  AND2X2 U142 ( .A(b[7]), .B(a[0]), .Y(n155) );
  AND2X2 U143 ( .A(a[1]), .B(b[7]), .Y(n147) );
  AND2X2 U144 ( .A(a[3]), .B(b[7]), .Y(n131) );
  AND2X2 U145 ( .A(a[6]), .B(b[6]), .Y(n108) );
  AND2X2 U146 ( .A(n214), .B(b[6]), .Y(n116) );
  AND2X2 U147 ( .A(a[4]), .B(b[6]), .Y(n124) );
  AND2X2 U148 ( .A(a[3]), .B(b[6]), .Y(n132) );
  AND2X2 U149 ( .A(a[2]), .B(b[6]), .Y(n140) );
  AND2X2 U150 ( .A(a[1]), .B(b[6]), .Y(n148) );
  AND2X2 U151 ( .A(b[6]), .B(a[0]), .Y(n156) );
  AND2X1 U152 ( .A(n214), .B(b[4]), .Y(n118) );
  AND2X1 U153 ( .A(b[3]), .B(a[7]), .Y(n103) );
  AND2X1 U154 ( .A(n214), .B(b[3]), .Y(n119) );
  AND2X1 U155 ( .A(a[3]), .B(b[5]), .Y(n133) );
  AND2X1 U156 ( .A(b[1]), .B(a[7]), .Y(n105) );
  AND2X1 U157 ( .A(a[3]), .B(b[2]), .Y(n136) );
  AND2X1 U158 ( .A(a[2]), .B(b[3]), .Y(n143) );
  AND2X1 U159 ( .A(a[3]), .B(b[4]), .Y(n134) );
  AND2X1 U160 ( .A(a[4]), .B(b[3]), .Y(n127) );
  AND2X1 U161 ( .A(n214), .B(b[2]), .Y(n120) );
  AND2X1 U162 ( .A(a[1]), .B(b[5]), .Y(n149) );
  AND2X1 U163 ( .A(a[4]), .B(b[2]), .Y(n128) );
  AND2X1 U164 ( .A(a[5]), .B(b[1]), .Y(n121) );
  AND2X1 U165 ( .A(n214), .B(b[5]), .Y(n117) );
  AND2X1 U166 ( .A(a[3]), .B(b[3]), .Y(n135) );
  AND2X1 U167 ( .A(a[2]), .B(b[2]), .Y(n144) );
  AND2X1 U168 ( .A(a[1]), .B(b[3]), .Y(n151) );
  AND2X1 U169 ( .A(a[3]), .B(b[1]), .Y(n137) );
  AND2X1 U170 ( .A(a[3]), .B(b[0]), .Y(n138) );
  AND2X1 U171 ( .A(a[1]), .B(b[1]), .Y(n153) );
  AND2X1 U172 ( .A(a[1]), .B(b[0]), .Y(n154) );
  AND2X2 U173 ( .A(b[6]), .B(a[7]), .Y(n100) );
  AND2X2 U174 ( .A(a[4]), .B(b[1]), .Y(n129) );
  BUFX2 U175 ( .A(a[5]), .Y(n214) );
  AND2X2 U176 ( .A(a[1]), .B(b[4]), .Y(n150) );
  AND2X2 U177 ( .A(a[1]), .B(b[2]), .Y(n152) );
  AND2X2 U178 ( .A(a[6]), .B(b[3]), .Y(n111) );
  AND2X2 U179 ( .A(b[3]), .B(a[0]), .Y(n159) );
  AND2X2 U180 ( .A(a[6]), .B(b[7]), .Y(n107) );
  AND2X2 U181 ( .A(n214), .B(b[7]), .Y(n115) );
  AND2X2 U182 ( .A(a[2]), .B(b[7]), .Y(n139) );
  AND2X1 U183 ( .A(a[5]), .B(b[0]), .Y(n122) );
  AND2X1 U184 ( .A(b[0]), .B(a[0]), .Y(product[0]) );
  AND2X1 U185 ( .A(b[1]), .B(a[0]), .Y(n161) );
  AND2X1 U186 ( .A(b[2]), .B(a[0]), .Y(n160) );
  AND2X1 U187 ( .A(b[4]), .B(a[0]), .Y(n158) );
  AND2X1 U188 ( .A(b[5]), .B(a[0]), .Y(n157) );
  AND2X1 U189 ( .A(a[2]), .B(b[0]), .Y(n146) );
  AND2X1 U190 ( .A(a[2]), .B(b[1]), .Y(n145) );
  AND2X1 U191 ( .A(a[2]), .B(b[4]), .Y(n142) );
  AND2X1 U192 ( .A(a[2]), .B(b[5]), .Y(n141) );
  AND2X1 U193 ( .A(a[4]), .B(b[0]), .Y(n130) );
  AND2X1 U194 ( .A(a[4]), .B(b[4]), .Y(n126) );
  AND2X1 U195 ( .A(a[4]), .B(b[5]), .Y(n125) );
  AND2X1 U196 ( .A(a[6]), .B(b[0]), .Y(n114) );
  AND2X1 U197 ( .A(a[6]), .B(b[1]), .Y(n113) );
  AND2X1 U198 ( .A(a[6]), .B(b[2]), .Y(n112) );
  AND2X1 U199 ( .A(a[6]), .B(b[4]), .Y(n110) );
  AND2X1 U200 ( .A(a[6]), .B(b[5]), .Y(n109) );
  AND2X1 U201 ( .A(a[7]), .B(b[0]), .Y(n106) );
  AND2X1 U202 ( .A(b[2]), .B(a[7]), .Y(n104) );
  AND2X1 U203 ( .A(b[4]), .B(a[7]), .Y(n102) );
  AND2X1 U204 ( .A(b[5]), .B(a[7]), .Y(n101) );
endmodule


module alu_DW_mult_uns_11 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71;
  assign product[0] = b[0];

  FAX1 U2 ( .A(a[7]), .B(n44), .C(n2), .YC(product[15]), .YS(product[14]) );
  FAX1 U3 ( .A(n45), .B(n14), .C(n3), .YC(n2), .YS(product[13]) );
  FAX1 U4 ( .A(n15), .B(n16), .C(n4), .YC(n3), .YS(product[12]) );
  FAX1 U5 ( .A(n17), .B(n18), .C(n5), .YC(n4), .YS(product[11]) );
  FAX1 U6 ( .A(n22), .B(n19), .C(n6), .YC(n5), .YS(product[10]) );
  FAX1 U7 ( .A(n26), .B(n23), .C(n7), .YC(n6), .YS(product[9]) );
  FAX1 U8 ( .A(n32), .B(n27), .C(n8), .YC(n7), .YS(product[8]) );
  FAX1 U9 ( .A(n36), .B(n33), .C(n9), .YC(n8), .YS(product[7]) );
  FAX1 U10 ( .A(n39), .B(n37), .C(n10), .YC(n9), .YS(product[6]) );
  FAX1 U11 ( .A(n42), .B(n41), .C(n11), .YC(n10), .YS(product[5]) );
  FAX1 U12 ( .A(n68), .B(n43), .C(n12), .YC(n11), .YS(product[4]) );
  HAX1 U13 ( .A(n70), .B(n13), .YC(n12), .YS(product[3]) );
  HAX1 U14 ( .A(a[1]), .B(n71), .YC(n13), .YS(product[2]) );
  FAX1 U15 ( .A(a[6]), .B(n51), .C(n46), .YC(n14), .YS(n15) );
  FAX1 U16 ( .A(n52), .B(n47), .C(n20), .YC(n16), .YS(n17) );
  FAX1 U17 ( .A(n53), .B(n24), .C(n21), .YC(n18), .YS(n19) );
  FAX1 U18 ( .A(a[5]), .B(n57), .C(n48), .YC(n20), .YS(n21) );
  FAX1 U19 ( .A(n30), .B(n28), .C(n25), .YC(n22), .YS(n23) );
  FAX1 U20 ( .A(n58), .B(n49), .C(n54), .YC(n24), .YS(n25) );
  FAX1 U21 ( .A(n34), .B(n31), .C(n29), .YC(n26), .YS(n27) );
  FAX1 U22 ( .A(n62), .B(n50), .C(n59), .YC(n28), .YS(n29) );
  HAX1 U23 ( .A(a[4]), .B(n55), .YC(n30), .YS(n31) );
  FAX1 U24 ( .A(n60), .B(n38), .C(n35), .YC(n32), .YS(n33) );
  HAX1 U25 ( .A(n63), .B(n56), .YC(n34), .YS(n35) );
  FAX1 U26 ( .A(n64), .B(n61), .C(n40), .YC(n36), .YS(n37) );
  HAX1 U27 ( .A(a[3]), .B(n66), .YC(n38), .YS(n39) );
  HAX1 U28 ( .A(n67), .B(n65), .YC(n40), .YS(n41) );
  HAX1 U29 ( .A(a[2]), .B(n69), .YC(n42), .YS(n43) );
  AND2X1 U75 ( .A(b[5]), .B(b[3]), .Y(n58) );
  AND2X1 U76 ( .A(b[5]), .B(b[4]), .Y(n57) );
  AND2X1 U77 ( .A(b[2]), .B(b[0]), .Y(n70) );
  AND2X1 U78 ( .A(b[5]), .B(b[2]), .Y(n59) );
  AND2X1 U79 ( .A(b[6]), .B(b[1]), .Y(n55) );
  AND2X1 U80 ( .A(b[6]), .B(b[4]), .Y(n52) );
  AND2X1 U81 ( .A(b[7]), .B(b[3]), .Y(n47) );
  AND2X1 U82 ( .A(b[6]), .B(b[3]), .Y(n53) );
  AND2X1 U83 ( .A(b[6]), .B(b[0]), .Y(n56) );
  AND2X1 U84 ( .A(b[3]), .B(b[0]), .Y(n68) );
  AND2X1 U85 ( .A(b[3]), .B(b[2]), .Y(n66) );
  AND2X1 U86 ( .A(b[5]), .B(b[0]), .Y(n61) );
  AND2X1 U87 ( .A(b[7]), .B(b[6]), .Y(n44) );
  AND2X1 U88 ( .A(b[1]), .B(b[0]), .Y(n71) );
  AND2X1 U89 ( .A(b[4]), .B(b[0]), .Y(n65) );
  AND2X1 U90 ( .A(b[4]), .B(b[1]), .Y(n64) );
  AND2X1 U91 ( .A(b[4]), .B(b[2]), .Y(n63) );
  AND2X1 U92 ( .A(b[4]), .B(b[3]), .Y(n62) );
  AND2X2 U93 ( .A(b[7]), .B(b[1]), .Y(n49) );
  AND2X2 U94 ( .A(b[7]), .B(b[2]), .Y(n48) );
  AND2X2 U95 ( .A(b[2]), .B(b[1]), .Y(n69) );
  AND2X2 U96 ( .A(b[6]), .B(b[2]), .Y(n54) );
  AND2X2 U97 ( .A(b[3]), .B(b[1]), .Y(n67) );
  AND2X2 U98 ( .A(b[7]), .B(b[5]), .Y(n45) );
  AND2X2 U99 ( .A(b[6]), .B(b[5]), .Y(n51) );
  AND2X2 U100 ( .A(b[5]), .B(b[1]), .Y(n60) );
  AND2X2 U101 ( .A(b[7]), .B(b[4]), .Y(n46) );
  AND2X1 U102 ( .A(b[7]), .B(b[0]), .Y(n50) );
endmodule


module alu_DW_mult_uns_10 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n214;

  FAX1 U2 ( .A(n99), .B(n15), .C(n2), .YC(product[15]), .YS(product[14]) );
  FAX1 U3 ( .A(n16), .B(n17), .C(n3), .YC(n2), .YS(product[13]) );
  FAX1 U4 ( .A(n18), .B(n21), .C(n4), .YC(n3), .YS(product[12]) );
  FAX1 U5 ( .A(n22), .B(n27), .C(n5), .YC(n4), .YS(product[11]) );
  FAX1 U6 ( .A(n35), .B(n28), .C(n6), .YC(n5), .YS(product[10]) );
  FAX1 U7 ( .A(n45), .B(n36), .C(n7), .YC(n6), .YS(product[9]) );
  FAX1 U8 ( .A(n57), .B(n46), .C(n8), .YC(n7), .YS(product[8]) );
  FAX1 U9 ( .A(n69), .B(n58), .C(n9), .YC(n8), .YS(product[7]) );
  FAX1 U10 ( .A(n79), .B(n70), .C(n10), .YC(n9), .YS(product[6]) );
  FAX1 U11 ( .A(n87), .B(n80), .C(n11), .YC(n10), .YS(product[5]) );
  FAX1 U12 ( .A(n93), .B(n88), .C(n12), .YC(n11), .YS(product[4]) );
  FAX1 U13 ( .A(n96), .B(n94), .C(n13), .YC(n12), .YS(product[3]) );
  FAX1 U14 ( .A(n146), .B(n14), .C(n98), .YC(n13), .YS(product[2]) );
  HAX1 U15 ( .A(n154), .B(n161), .YC(n14), .YS(product[1]) );
  FAX1 U16 ( .A(n107), .B(n100), .C(n19), .YC(n15), .YS(n16) );
  FAX1 U17 ( .A(n25), .B(n20), .C(n23), .YC(n17), .YS(n18) );
  FAX1 U18 ( .A(n115), .B(n101), .C(n108), .YC(n19), .YS(n20) );
  FAX1 U19 ( .A(n31), .B(n24), .C(n29), .YC(n21), .YS(n22) );
  FAX1 U20 ( .A(n116), .B(n33), .C(n26), .YC(n23), .YS(n24) );
  FAX1 U21 ( .A(n123), .B(n102), .C(n109), .YC(n25), .YS(n26) );
  FAX1 U22 ( .A(n39), .B(n37), .C(n30), .YC(n27), .YS(n28) );
  FAX1 U23 ( .A(n41), .B(n34), .C(n32), .YC(n29), .YS(n30) );
  FAX1 U24 ( .A(n124), .B(n117), .C(n43), .YC(n31), .YS(n32) );
  FAX1 U25 ( .A(n131), .B(n103), .C(n110), .YC(n33), .YS(n34) );
  FAX1 U26 ( .A(n40), .B(n47), .C(n38), .YC(n35), .YS(n36) );
  FAX1 U27 ( .A(n44), .B(n51), .C(n49), .YC(n37), .YS(n38) );
  FAX1 U28 ( .A(n55), .B(n53), .C(n42), .YC(n39), .YS(n40) );
  FAX1 U29 ( .A(n118), .B(n125), .C(n132), .YC(n41), .YS(n42) );
  FAX1 U30 ( .A(n139), .B(n104), .C(n111), .YC(n43), .YS(n44) );
  FAX1 U31 ( .A(n50), .B(n59), .C(n48), .YC(n45), .YS(n46) );
  FAX1 U32 ( .A(n54), .B(n52), .C(n61), .YC(n47), .YS(n48) );
  FAX1 U33 ( .A(n56), .B(n65), .C(n63), .YC(n49), .YS(n50) );
  FAX1 U34 ( .A(n140), .B(n133), .C(n67), .YC(n51), .YS(n52) );
  FAX1 U35 ( .A(n126), .B(n119), .C(n147), .YC(n53), .YS(n54) );
  HAX1 U36 ( .A(n112), .B(n105), .YC(n55), .YS(n56) );
  FAX1 U37 ( .A(n62), .B(n71), .C(n60), .YC(n57), .YS(n58) );
  FAX1 U38 ( .A(n64), .B(n66), .C(n73), .YC(n59), .YS(n60) );
  FAX1 U39 ( .A(n77), .B(n68), .C(n75), .YC(n61), .YS(n62) );
  FAX1 U40 ( .A(n141), .B(n127), .C(n134), .YC(n63), .YS(n64) );
  FAX1 U41 ( .A(n155), .B(n120), .C(n148), .YC(n65), .YS(n66) );
  HAX1 U42 ( .A(n113), .B(n106), .YC(n67), .YS(n68) );
  FAX1 U43 ( .A(n74), .B(n81), .C(n72), .YC(n69), .YS(n70) );
  FAX1 U44 ( .A(n78), .B(n83), .C(n76), .YC(n71), .YS(n72) );
  FAX1 U45 ( .A(n142), .B(n135), .C(n85), .YC(n73), .YS(n74) );
  FAX1 U46 ( .A(n156), .B(n128), .C(n149), .YC(n75), .YS(n76) );
  HAX1 U47 ( .A(n121), .B(n114), .YC(n77), .YS(n78) );
  FAX1 U48 ( .A(n89), .B(n84), .C(n82), .YC(n79), .YS(n80) );
  FAX1 U49 ( .A(n150), .B(n91), .C(n86), .YC(n81), .YS(n82) );
  FAX1 U50 ( .A(n157), .B(n136), .C(n143), .YC(n83), .YS(n84) );
  HAX1 U51 ( .A(n129), .B(n122), .YC(n85), .YS(n86) );
  FAX1 U52 ( .A(n95), .B(n92), .C(n90), .YC(n87), .YS(n88) );
  FAX1 U53 ( .A(n151), .B(n144), .C(n158), .YC(n89), .YS(n90) );
  HAX1 U54 ( .A(n137), .B(n130), .YC(n91), .YS(n92) );
  FAX1 U55 ( .A(n159), .B(n152), .C(n97), .YC(n93), .YS(n94) );
  HAX1 U56 ( .A(n145), .B(n138), .YC(n95), .YS(n96) );
  HAX1 U57 ( .A(n160), .B(n153), .YC(n97), .YS(n98) );
  BUFX2 U140 ( .A(b[1]), .Y(n214) );
  AND2X2 U141 ( .A(a[6]), .B(n214), .Y(n113) );
  AND2X2 U142 ( .A(a[6]), .B(b[2]), .Y(n112) );
  AND2X1 U143 ( .A(a[2]), .B(b[7]), .Y(n139) );
  AND2X1 U144 ( .A(a[3]), .B(b[5]), .Y(n133) );
  AND2X1 U145 ( .A(a[2]), .B(b[6]), .Y(n140) );
  AND2X1 U146 ( .A(a[3]), .B(b[7]), .Y(n131) );
  AND2X1 U147 ( .A(a[4]), .B(b[7]), .Y(n123) );
  AND2X1 U148 ( .A(a[5]), .B(b[0]), .Y(n122) );
  AND2X1 U149 ( .A(a[5]), .B(b[7]), .Y(n115) );
  AND2X1 U150 ( .A(b[0]), .B(a[0]), .Y(product[0]) );
  AND2X1 U151 ( .A(a[2]), .B(b[0]), .Y(n146) );
  AND2X1 U152 ( .A(a[4]), .B(b[5]), .Y(n125) );
  AND2X1 U153 ( .A(a[3]), .B(b[6]), .Y(n132) );
  AND2X1 U154 ( .A(a[1]), .B(b[7]), .Y(n147) );
  AND2X1 U155 ( .A(a[5]), .B(b[3]), .Y(n119) );
  AND2X1 U156 ( .A(n214), .B(a[7]), .Y(n105) );
  AND2X1 U157 ( .A(a[5]), .B(b[5]), .Y(n117) );
  AND2X1 U158 ( .A(a[4]), .B(b[6]), .Y(n124) );
  AND2X1 U159 ( .A(a[2]), .B(b[5]), .Y(n141) );
  AND2X1 U160 ( .A(a[1]), .B(b[6]), .Y(n148) );
  AND2X1 U161 ( .A(a[5]), .B(b[2]), .Y(n120) );
  AND2X1 U162 ( .A(a[7]), .B(b[0]), .Y(n106) );
  AND2X1 U163 ( .A(a[5]), .B(b[6]), .Y(n116) );
  AND2X1 U164 ( .A(a[3]), .B(b[1]), .Y(n137) );
  AND2X1 U165 ( .A(a[1]), .B(b[5]), .Y(n149) );
  AND2X1 U166 ( .A(a[6]), .B(b[0]), .Y(n114) );
  AND2X1 U167 ( .A(a[5]), .B(n214), .Y(n121) );
  AND2X1 U168 ( .A(a[1]), .B(b[3]), .Y(n151) );
  AND2X1 U169 ( .A(a[2]), .B(b[2]), .Y(n144) );
  AND2X1 U170 ( .A(a[2]), .B(b[3]), .Y(n143) );
  AND2X1 U171 ( .A(a[3]), .B(b[2]), .Y(n136) );
  AND2X1 U172 ( .A(a[3]), .B(b[3]), .Y(n135) );
  AND2X1 U173 ( .A(a[2]), .B(n214), .Y(n145) );
  AND2X1 U174 ( .A(a[3]), .B(b[0]), .Y(n138) );
  AND2X1 U175 ( .A(a[6]), .B(b[7]), .Y(n107) );
  AND2X1 U176 ( .A(b[2]), .B(a[0]), .Y(n160) );
  AND2X1 U177 ( .A(a[1]), .B(b[1]), .Y(n153) );
  AND2X1 U178 ( .A(a[4]), .B(b[0]), .Y(n130) );
  AND2X1 U179 ( .A(a[4]), .B(n214), .Y(n129) );
  AND2X1 U180 ( .A(a[4]), .B(b[2]), .Y(n128) );
  AND2X1 U181 ( .A(a[4]), .B(b[3]), .Y(n127) );
  AND2X2 U182 ( .A(b[4]), .B(a[7]), .Y(n102) );
  AND2X2 U183 ( .A(a[2]), .B(b[4]), .Y(n142) );
  AND2X2 U184 ( .A(b[4]), .B(a[0]), .Y(n158) );
  AND2X2 U185 ( .A(a[1]), .B(b[4]), .Y(n150) );
  AND2X2 U186 ( .A(a[6]), .B(b[6]), .Y(n108) );
  AND2X2 U187 ( .A(a[6]), .B(b[5]), .Y(n109) );
  AND2X2 U188 ( .A(a[6]), .B(b[4]), .Y(n110) );
  AND2X2 U189 ( .A(a[3]), .B(b[4]), .Y(n134) );
  AND2X2 U190 ( .A(a[1]), .B(b[0]), .Y(n154) );
  AND2X2 U191 ( .A(b[2]), .B(a[7]), .Y(n104) );
  AND2X2 U192 ( .A(a[5]), .B(b[4]), .Y(n118) );
  AND2X2 U193 ( .A(a[6]), .B(b[3]), .Y(n111) );
  AND2X2 U194 ( .A(b[1]), .B(a[0]), .Y(n161) );
  AND2X2 U195 ( .A(a[1]), .B(b[2]), .Y(n152) );
  AND2X2 U196 ( .A(a[4]), .B(b[4]), .Y(n126) );
  AND2X1 U197 ( .A(b[5]), .B(a[0]), .Y(n157) );
  AND2X1 U198 ( .A(b[7]), .B(a[0]), .Y(n155) );
  AND2X1 U199 ( .A(b[3]), .B(a[0]), .Y(n159) );
  AND2X1 U200 ( .A(b[6]), .B(a[0]), .Y(n156) );
  AND2X1 U201 ( .A(b[7]), .B(a[7]), .Y(n99) );
  AND2X1 U202 ( .A(b[3]), .B(a[7]), .Y(n103) );
  AND2X1 U203 ( .A(b[5]), .B(a[7]), .Y(n101) );
  AND2X1 U204 ( .A(b[6]), .B(a[7]), .Y(n100) );
endmodule


module alu_DW_mult_uns_15 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71;
  assign product[0] = b[0];

  FAX1 U2 ( .A(a[7]), .B(n44), .C(n2), .YC(product[15]), .YS(product[14]) );
  FAX1 U3 ( .A(n45), .B(n14), .C(n3), .YC(n2), .YS(product[13]) );
  FAX1 U4 ( .A(n15), .B(n16), .C(n4), .YC(n3), .YS(product[12]) );
  FAX1 U5 ( .A(n17), .B(n18), .C(n5), .YC(n4), .YS(product[11]) );
  FAX1 U6 ( .A(n22), .B(n19), .C(n6), .YC(n5), .YS(product[10]) );
  FAX1 U7 ( .A(n26), .B(n23), .C(n7), .YC(n6), .YS(product[9]) );
  FAX1 U8 ( .A(n32), .B(n27), .C(n8), .YC(n7), .YS(product[8]) );
  FAX1 U9 ( .A(n36), .B(n33), .C(n9), .YC(n8), .YS(product[7]) );
  FAX1 U10 ( .A(n39), .B(n37), .C(n10), .YC(n9), .YS(product[6]) );
  FAX1 U11 ( .A(n42), .B(n41), .C(n11), .YC(n10), .YS(product[5]) );
  FAX1 U12 ( .A(n68), .B(n43), .C(n12), .YC(n11), .YS(product[4]) );
  HAX1 U13 ( .A(n70), .B(n13), .YC(n12), .YS(product[3]) );
  HAX1 U14 ( .A(a[1]), .B(n71), .YC(n13), .YS(product[2]) );
  FAX1 U15 ( .A(a[6]), .B(n51), .C(n46), .YC(n14), .YS(n15) );
  FAX1 U16 ( .A(n52), .B(n47), .C(n20), .YC(n16), .YS(n17) );
  FAX1 U17 ( .A(n53), .B(n24), .C(n21), .YC(n18), .YS(n19) );
  FAX1 U18 ( .A(a[5]), .B(n57), .C(n48), .YC(n20), .YS(n21) );
  FAX1 U19 ( .A(n30), .B(n28), .C(n25), .YC(n22), .YS(n23) );
  FAX1 U20 ( .A(n58), .B(n49), .C(n54), .YC(n24), .YS(n25) );
  FAX1 U21 ( .A(n34), .B(n31), .C(n29), .YC(n26), .YS(n27) );
  FAX1 U22 ( .A(n62), .B(n50), .C(n59), .YC(n28), .YS(n29) );
  HAX1 U23 ( .A(a[4]), .B(n55), .YC(n30), .YS(n31) );
  FAX1 U24 ( .A(n60), .B(n38), .C(n35), .YC(n32), .YS(n33) );
  HAX1 U25 ( .A(n63), .B(n56), .YC(n34), .YS(n35) );
  FAX1 U26 ( .A(n64), .B(n61), .C(n40), .YC(n36), .YS(n37) );
  HAX1 U27 ( .A(a[3]), .B(n66), .YC(n38), .YS(n39) );
  HAX1 U28 ( .A(n67), .B(n65), .YC(n40), .YS(n41) );
  HAX1 U29 ( .A(a[2]), .B(n69), .YC(n42), .YS(n43) );
  AND2X2 U75 ( .A(b[7]), .B(b[0]), .Y(n50) );
  AND2X2 U76 ( .A(b[6]), .B(b[0]), .Y(n56) );
  AND2X2 U77 ( .A(b[5]), .B(b[0]), .Y(n61) );
  AND2X2 U78 ( .A(b[4]), .B(b[0]), .Y(n65) );
  AND2X2 U79 ( .A(b[3]), .B(b[0]), .Y(n68) );
  AND2X2 U80 ( .A(b[1]), .B(b[0]), .Y(n71) );
  AND2X1 U81 ( .A(b[3]), .B(b[1]), .Y(n67) );
  AND2X1 U82 ( .A(b[5]), .B(b[4]), .Y(n57) );
  AND2X1 U83 ( .A(b[5]), .B(b[3]), .Y(n58) );
  AND2X1 U84 ( .A(b[5]), .B(b[2]), .Y(n59) );
  AND2X1 U85 ( .A(b[6]), .B(b[5]), .Y(n51) );
  AND2X1 U86 ( .A(b[3]), .B(b[2]), .Y(n66) );
  AND2X1 U87 ( .A(b[4]), .B(b[3]), .Y(n62) );
  AND2X2 U88 ( .A(b[2]), .B(b[0]), .Y(n70) );
  AND2X2 U89 ( .A(b[7]), .B(b[5]), .Y(n45) );
  AND2X2 U90 ( .A(b[5]), .B(b[1]), .Y(n60) );
  AND2X1 U91 ( .A(b[7]), .B(b[2]), .Y(n48) );
  AND2X1 U92 ( .A(b[2]), .B(b[1]), .Y(n69) );
  AND2X1 U93 ( .A(b[4]), .B(b[1]), .Y(n64) );
  AND2X1 U94 ( .A(b[4]), .B(b[2]), .Y(n63) );
  AND2X1 U95 ( .A(b[6]), .B(b[1]), .Y(n55) );
  AND2X1 U96 ( .A(b[6]), .B(b[2]), .Y(n54) );
  AND2X1 U97 ( .A(b[6]), .B(b[3]), .Y(n53) );
  AND2X1 U98 ( .A(b[6]), .B(b[4]), .Y(n52) );
  AND2X1 U99 ( .A(b[7]), .B(b[1]), .Y(n49) );
  AND2X1 U100 ( .A(b[7]), .B(b[3]), .Y(n47) );
  AND2X1 U101 ( .A(b[7]), .B(b[4]), .Y(n46) );
  AND2X1 U102 ( .A(b[7]), .B(b[6]), .Y(n44) );
endmodule


module alu_DW_mult_uns_14 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n214, n215;

  FAX1 U2 ( .A(n99), .B(n15), .C(n2), .YC(product[15]), .YS(product[14]) );
  FAX1 U3 ( .A(n16), .B(n17), .C(n3), .YC(n2), .YS(product[13]) );
  FAX1 U4 ( .A(n18), .B(n21), .C(n4), .YC(n3), .YS(product[12]) );
  FAX1 U5 ( .A(n22), .B(n27), .C(n5), .YC(n4), .YS(product[11]) );
  FAX1 U6 ( .A(n35), .B(n28), .C(n6), .YC(n5), .YS(product[10]) );
  FAX1 U7 ( .A(n45), .B(n36), .C(n7), .YC(n6), .YS(product[9]) );
  FAX1 U8 ( .A(n57), .B(n46), .C(n8), .YC(n7), .YS(product[8]) );
  FAX1 U9 ( .A(n69), .B(n58), .C(n9), .YC(n8), .YS(product[7]) );
  FAX1 U10 ( .A(n79), .B(n70), .C(n10), .YC(n9), .YS(product[6]) );
  FAX1 U11 ( .A(n87), .B(n80), .C(n11), .YC(n10), .YS(product[5]) );
  FAX1 U12 ( .A(n93), .B(n88), .C(n12), .YC(n11), .YS(product[4]) );
  FAX1 U13 ( .A(n96), .B(n13), .C(n94), .YC(n12), .YS(product[3]) );
  FAX1 U14 ( .A(n146), .B(n14), .C(n98), .YC(n13), .YS(product[2]) );
  HAX1 U15 ( .A(n154), .B(n161), .YC(n14), .YS(product[1]) );
  FAX1 U16 ( .A(n107), .B(n100), .C(n19), .YC(n15), .YS(n16) );
  FAX1 U17 ( .A(n25), .B(n20), .C(n23), .YC(n17), .YS(n18) );
  FAX1 U18 ( .A(n115), .B(n101), .C(n108), .YC(n19), .YS(n20) );
  FAX1 U19 ( .A(n31), .B(n24), .C(n29), .YC(n21), .YS(n22) );
  FAX1 U20 ( .A(n116), .B(n33), .C(n26), .YC(n23), .YS(n24) );
  FAX1 U21 ( .A(n123), .B(n102), .C(n109), .YC(n25), .YS(n26) );
  FAX1 U22 ( .A(n39), .B(n37), .C(n30), .YC(n27), .YS(n28) );
  FAX1 U23 ( .A(n41), .B(n34), .C(n32), .YC(n29), .YS(n30) );
  FAX1 U24 ( .A(n124), .B(n117), .C(n43), .YC(n31), .YS(n32) );
  FAX1 U25 ( .A(n131), .B(n103), .C(n110), .YC(n33), .YS(n34) );
  FAX1 U26 ( .A(n40), .B(n47), .C(n38), .YC(n35), .YS(n36) );
  FAX1 U27 ( .A(n44), .B(n51), .C(n49), .YC(n37), .YS(n38) );
  FAX1 U28 ( .A(n55), .B(n53), .C(n42), .YC(n39), .YS(n40) );
  FAX1 U29 ( .A(n118), .B(n125), .C(n132), .YC(n41), .YS(n42) );
  FAX1 U30 ( .A(n139), .B(n104), .C(n111), .YC(n43), .YS(n44) );
  FAX1 U31 ( .A(n50), .B(n59), .C(n48), .YC(n45), .YS(n46) );
  FAX1 U32 ( .A(n54), .B(n52), .C(n61), .YC(n47), .YS(n48) );
  FAX1 U33 ( .A(n56), .B(n65), .C(n63), .YC(n49), .YS(n50) );
  FAX1 U34 ( .A(n140), .B(n133), .C(n67), .YC(n51), .YS(n52) );
  FAX1 U35 ( .A(n126), .B(n119), .C(n147), .YC(n53), .YS(n54) );
  HAX1 U36 ( .A(n112), .B(n105), .YC(n55), .YS(n56) );
  FAX1 U37 ( .A(n62), .B(n71), .C(n60), .YC(n57), .YS(n58) );
  FAX1 U38 ( .A(n64), .B(n66), .C(n73), .YC(n59), .YS(n60) );
  FAX1 U39 ( .A(n77), .B(n68), .C(n75), .YC(n61), .YS(n62) );
  FAX1 U40 ( .A(n141), .B(n127), .C(n134), .YC(n63), .YS(n64) );
  FAX1 U41 ( .A(n155), .B(n120), .C(n148), .YC(n65), .YS(n66) );
  HAX1 U42 ( .A(n113), .B(n106), .YC(n67), .YS(n68) );
  FAX1 U43 ( .A(n74), .B(n81), .C(n72), .YC(n69), .YS(n70) );
  FAX1 U44 ( .A(n78), .B(n83), .C(n76), .YC(n71), .YS(n72) );
  FAX1 U45 ( .A(n142), .B(n135), .C(n85), .YC(n73), .YS(n74) );
  FAX1 U46 ( .A(n156), .B(n128), .C(n149), .YC(n75), .YS(n76) );
  HAX1 U47 ( .A(n121), .B(n114), .YC(n77), .YS(n78) );
  FAX1 U48 ( .A(n89), .B(n84), .C(n82), .YC(n79), .YS(n80) );
  FAX1 U49 ( .A(n150), .B(n91), .C(n86), .YC(n81), .YS(n82) );
  FAX1 U50 ( .A(n157), .B(n136), .C(n143), .YC(n83), .YS(n84) );
  HAX1 U51 ( .A(n129), .B(n122), .YC(n85), .YS(n86) );
  FAX1 U52 ( .A(n95), .B(n92), .C(n90), .YC(n87), .YS(n88) );
  FAX1 U53 ( .A(n158), .B(n144), .C(n151), .YC(n89), .YS(n90) );
  HAX1 U54 ( .A(n137), .B(n130), .YC(n91), .YS(n92) );
  FAX1 U55 ( .A(n159), .B(n152), .C(n97), .YC(n93), .YS(n94) );
  HAX1 U56 ( .A(n145), .B(n138), .YC(n95), .YS(n96) );
  HAX1 U57 ( .A(n160), .B(n153), .YC(n97), .YS(n98) );
  BUFX2 U140 ( .A(b[1]), .Y(n214) );
  AND2X2 U141 ( .A(b[7]), .B(a[0]), .Y(n155) );
  AND2X2 U142 ( .A(b[6]), .B(a[0]), .Y(n156) );
  AND2X2 U143 ( .A(b[5]), .B(a[0]), .Y(n157) );
  AND2X2 U144 ( .A(b[2]), .B(a[0]), .Y(n160) );
  AND2X2 U145 ( .A(a[4]), .B(b[1]), .Y(n129) );
  AND2X2 U146 ( .A(a[2]), .B(n214), .Y(n145) );
  AND2X2 U147 ( .A(a[3]), .B(b[1]), .Y(n137) );
  AND2X2 U148 ( .A(b[1]), .B(a[0]), .Y(n161) );
  AND2X2 U149 ( .A(a[1]), .B(b[1]), .Y(n153) );
  AND2X1 U150 ( .A(a[6]), .B(b[2]), .Y(n112) );
  AND2X1 U151 ( .A(n215), .B(a[7]), .Y(n105) );
  AND2X1 U152 ( .A(a[5]), .B(b[5]), .Y(n117) );
  AND2X1 U153 ( .A(a[4]), .B(b[6]), .Y(n124) );
  AND2X1 U154 ( .A(a[5]), .B(b[6]), .Y(n116) );
  AND2X1 U155 ( .A(a[6]), .B(n215), .Y(n113) );
  AND2X1 U156 ( .A(a[7]), .B(b[0]), .Y(n106) );
  AND2X1 U157 ( .A(a[5]), .B(b[2]), .Y(n120) );
  AND2X1 U158 ( .A(a[1]), .B(b[6]), .Y(n148) );
  AND2X1 U159 ( .A(a[1]), .B(b[5]), .Y(n149) );
  AND2X1 U160 ( .A(a[4]), .B(b[2]), .Y(n128) );
  AND2X1 U161 ( .A(a[6]), .B(b[0]), .Y(n114) );
  AND2X1 U162 ( .A(a[5]), .B(n215), .Y(n121) );
  AND2X1 U163 ( .A(a[5]), .B(b[0]), .Y(n122) );
  AND2X1 U164 ( .A(a[2]), .B(b[3]), .Y(n143) );
  AND2X1 U165 ( .A(a[3]), .B(b[2]), .Y(n136) );
  AND2X1 U166 ( .A(a[4]), .B(b[0]), .Y(n130) );
  AND2X1 U167 ( .A(a[3]), .B(b[0]), .Y(n138) );
  AND2X1 U168 ( .A(b[7]), .B(a[7]), .Y(n99) );
  AND2X1 U169 ( .A(a[1]), .B(b[0]), .Y(n154) );
  AND2X2 U170 ( .A(b[3]), .B(a[0]), .Y(n159) );
  AND2X2 U171 ( .A(b[4]), .B(a[7]), .Y(n102) );
  AND2X2 U172 ( .A(a[6]), .B(b[4]), .Y(n110) );
  AND2X2 U173 ( .A(a[4]), .B(b[4]), .Y(n126) );
  AND2X2 U174 ( .A(a[3]), .B(b[4]), .Y(n134) );
  AND2X2 U175 ( .A(a[1]), .B(b[4]), .Y(n150) );
  AND2X2 U176 ( .A(b[4]), .B(a[0]), .Y(n158) );
  BUFX2 U177 ( .A(n214), .Y(n215) );
  AND2X2 U178 ( .A(a[2]), .B(b[4]), .Y(n142) );
  AND2X2 U179 ( .A(b[0]), .B(a[0]), .Y(product[0]) );
  AND2X2 U180 ( .A(a[2]), .B(b[0]), .Y(n146) );
  AND2X2 U181 ( .A(a[6]), .B(b[7]), .Y(n107) );
  AND2X2 U182 ( .A(a[5]), .B(b[7]), .Y(n115) );
  AND2X2 U183 ( .A(a[4]), .B(b[7]), .Y(n123) );
  AND2X2 U184 ( .A(a[3]), .B(b[7]), .Y(n131) );
  AND2X2 U185 ( .A(a[2]), .B(b[7]), .Y(n139) );
  AND2X2 U186 ( .A(a[1]), .B(b[7]), .Y(n147) );
  AND2X2 U187 ( .A(b[6]), .B(a[7]), .Y(n100) );
  AND2X2 U188 ( .A(a[6]), .B(b[6]), .Y(n108) );
  AND2X2 U189 ( .A(a[3]), .B(b[6]), .Y(n132) );
  AND2X2 U190 ( .A(a[2]), .B(b[6]), .Y(n140) );
  AND2X2 U191 ( .A(b[2]), .B(a[7]), .Y(n104) );
  AND2X2 U192 ( .A(a[1]), .B(b[2]), .Y(n152) );
  AND2X2 U193 ( .A(a[2]), .B(b[2]), .Y(n144) );
  AND2X2 U194 ( .A(b[5]), .B(a[7]), .Y(n101) );
  AND2X2 U195 ( .A(a[6]), .B(b[5]), .Y(n109) );
  AND2X2 U196 ( .A(a[4]), .B(b[5]), .Y(n125) );
  AND2X2 U197 ( .A(a[3]), .B(b[5]), .Y(n133) );
  AND2X2 U198 ( .A(a[2]), .B(b[5]), .Y(n141) );
  AND2X2 U199 ( .A(a[5]), .B(b[3]), .Y(n119) );
  AND2X2 U200 ( .A(a[5]), .B(b[4]), .Y(n118) );
  AND2X1 U201 ( .A(a[1]), .B(b[3]), .Y(n151) );
  AND2X1 U202 ( .A(a[3]), .B(b[3]), .Y(n135) );
  AND2X1 U203 ( .A(a[4]), .B(b[3]), .Y(n127) );
  AND2X1 U204 ( .A(a[6]), .B(b[3]), .Y(n111) );
  AND2X1 U205 ( .A(b[3]), .B(a[7]), .Y(n103) );
endmodule


module alu_DW_mult_uns_6 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161;

  FAX1 U2 ( .A(n99), .B(n15), .C(n2), .YC(product[15]), .YS(product[14]) );
  FAX1 U3 ( .A(n16), .B(n17), .C(n3), .YC(n2), .YS(product[13]) );
  FAX1 U4 ( .A(n18), .B(n21), .C(n4), .YC(n3), .YS(product[12]) );
  FAX1 U5 ( .A(n22), .B(n27), .C(n5), .YC(n4), .YS(product[11]) );
  FAX1 U6 ( .A(n35), .B(n28), .C(n6), .YC(n5), .YS(product[10]) );
  FAX1 U7 ( .A(n45), .B(n36), .C(n7), .YC(n6), .YS(product[9]) );
  FAX1 U8 ( .A(n57), .B(n46), .C(n8), .YC(n7), .YS(product[8]) );
  FAX1 U9 ( .A(n69), .B(n58), .C(n9), .YC(n8), .YS(product[7]) );
  FAX1 U10 ( .A(n79), .B(n70), .C(n10), .YC(n9), .YS(product[6]) );
  FAX1 U11 ( .A(n87), .B(n80), .C(n11), .YC(n10), .YS(product[5]) );
  FAX1 U12 ( .A(n93), .B(n88), .C(n12), .YC(n11), .YS(product[4]) );
  FAX1 U13 ( .A(n96), .B(n94), .C(n13), .YC(n12), .YS(product[3]) );
  FAX1 U14 ( .A(n146), .B(n14), .C(n98), .YC(n13), .YS(product[2]) );
  HAX1 U15 ( .A(n154), .B(n161), .YC(n14), .YS(product[1]) );
  FAX1 U16 ( .A(n107), .B(n100), .C(n19), .YC(n15), .YS(n16) );
  FAX1 U17 ( .A(n25), .B(n20), .C(n23), .YC(n17), .YS(n18) );
  FAX1 U18 ( .A(n115), .B(n101), .C(n108), .YC(n19), .YS(n20) );
  FAX1 U19 ( .A(n31), .B(n24), .C(n29), .YC(n21), .YS(n22) );
  FAX1 U20 ( .A(n116), .B(n33), .C(n26), .YC(n23), .YS(n24) );
  FAX1 U21 ( .A(n123), .B(n102), .C(n109), .YC(n25), .YS(n26) );
  FAX1 U22 ( .A(n39), .B(n37), .C(n30), .YC(n27), .YS(n28) );
  FAX1 U23 ( .A(n41), .B(n34), .C(n32), .YC(n29), .YS(n30) );
  FAX1 U24 ( .A(n124), .B(n117), .C(n43), .YC(n31), .YS(n32) );
  FAX1 U25 ( .A(n131), .B(n103), .C(n110), .YC(n33), .YS(n34) );
  FAX1 U26 ( .A(n40), .B(n47), .C(n38), .YC(n35), .YS(n36) );
  FAX1 U27 ( .A(n44), .B(n51), .C(n49), .YC(n37), .YS(n38) );
  FAX1 U28 ( .A(n55), .B(n53), .C(n42), .YC(n39), .YS(n40) );
  FAX1 U29 ( .A(n118), .B(n125), .C(n132), .YC(n41), .YS(n42) );
  FAX1 U30 ( .A(n139), .B(n104), .C(n111), .YC(n43), .YS(n44) );
  FAX1 U31 ( .A(n50), .B(n59), .C(n48), .YC(n45), .YS(n46) );
  FAX1 U32 ( .A(n54), .B(n52), .C(n61), .YC(n47), .YS(n48) );
  FAX1 U33 ( .A(n56), .B(n65), .C(n63), .YC(n49), .YS(n50) );
  FAX1 U34 ( .A(n140), .B(n133), .C(n67), .YC(n51), .YS(n52) );
  FAX1 U35 ( .A(n126), .B(n119), .C(n147), .YC(n53), .YS(n54) );
  HAX1 U36 ( .A(n112), .B(n105), .YC(n55), .YS(n56) );
  FAX1 U37 ( .A(n62), .B(n71), .C(n60), .YC(n57), .YS(n58) );
  FAX1 U38 ( .A(n64), .B(n66), .C(n73), .YC(n59), .YS(n60) );
  FAX1 U39 ( .A(n77), .B(n68), .C(n75), .YC(n61), .YS(n62) );
  FAX1 U40 ( .A(n141), .B(n127), .C(n134), .YC(n63), .YS(n64) );
  FAX1 U41 ( .A(n155), .B(n120), .C(n148), .YC(n65), .YS(n66) );
  HAX1 U42 ( .A(n113), .B(n106), .YC(n67), .YS(n68) );
  FAX1 U43 ( .A(n74), .B(n81), .C(n72), .YC(n69), .YS(n70) );
  FAX1 U44 ( .A(n78), .B(n83), .C(n76), .YC(n71), .YS(n72) );
  FAX1 U45 ( .A(n142), .B(n135), .C(n85), .YC(n73), .YS(n74) );
  FAX1 U46 ( .A(n156), .B(n128), .C(n149), .YC(n75), .YS(n76) );
  HAX1 U47 ( .A(n121), .B(n114), .YC(n77), .YS(n78) );
  FAX1 U48 ( .A(n89), .B(n84), .C(n82), .YC(n79), .YS(n80) );
  FAX1 U49 ( .A(n150), .B(n91), .C(n86), .YC(n81), .YS(n82) );
  FAX1 U50 ( .A(n157), .B(n136), .C(n143), .YC(n83), .YS(n84) );
  HAX1 U51 ( .A(n129), .B(n122), .YC(n85), .YS(n86) );
  FAX1 U52 ( .A(n95), .B(n92), .C(n90), .YC(n87), .YS(n88) );
  FAX1 U53 ( .A(n158), .B(n144), .C(n151), .YC(n89), .YS(n90) );
  HAX1 U54 ( .A(n137), .B(n130), .YC(n91), .YS(n92) );
  FAX1 U55 ( .A(n159), .B(n152), .C(n97), .YC(n93), .YS(n94) );
  HAX1 U56 ( .A(n145), .B(n138), .YC(n95), .YS(n96) );
  HAX1 U57 ( .A(n160), .B(n153), .YC(n97), .YS(n98) );
  AND2X1 U140 ( .A(a[6]), .B(b[6]), .Y(n108) );
  AND2X1 U141 ( .A(a[2]), .B(b[0]), .Y(n146) );
  AND2X1 U142 ( .A(a[3]), .B(b[6]), .Y(n132) );
  AND2X1 U143 ( .A(a[4]), .B(b[6]), .Y(n124) );
  AND2X1 U144 ( .A(a[5]), .B(b[6]), .Y(n116) );
  AND2X1 U145 ( .A(a[3]), .B(b[5]), .Y(n133) );
  AND2X1 U146 ( .A(a[2]), .B(b[6]), .Y(n140) );
  AND2X1 U147 ( .A(a[1]), .B(b[7]), .Y(n147) );
  AND2X1 U148 ( .A(a[3]), .B(b[4]), .Y(n134) );
  AND2X1 U149 ( .A(a[2]), .B(b[5]), .Y(n141) );
  AND2X1 U150 ( .A(a[1]), .B(b[6]), .Y(n148) );
  AND2X1 U151 ( .A(b[6]), .B(a[0]), .Y(n156) );
  AND2X1 U152 ( .A(a[1]), .B(b[5]), .Y(n149) );
  AND2X1 U153 ( .A(a[2]), .B(b[1]), .Y(n145) );
  AND2X1 U154 ( .A(a[3]), .B(b[0]), .Y(n138) );
  AND2X1 U155 ( .A(a[1]), .B(b[1]), .Y(n153) );
  AND2X1 U156 ( .A(b[6]), .B(a[7]), .Y(n100) );
  AND2X1 U157 ( .A(a[1]), .B(b[3]), .Y(n151) );
  AND2X1 U158 ( .A(a[2]), .B(b[2]), .Y(n144) );
  AND2X1 U159 ( .A(a[3]), .B(b[2]), .Y(n136) );
  AND2X1 U160 ( .A(a[2]), .B(b[3]), .Y(n143) );
  AND2X1 U161 ( .A(a[1]), .B(b[4]), .Y(n150) );
  AND2X1 U162 ( .A(a[3]), .B(b[3]), .Y(n135) );
  AND2X1 U163 ( .A(a[2]), .B(b[4]), .Y(n142) );
  AND2X1 U164 ( .A(a[1]), .B(b[0]), .Y(n154) );
  AND2X2 U165 ( .A(a[2]), .B(b[7]), .Y(n139) );
  AND2X2 U166 ( .A(a[1]), .B(b[2]), .Y(n152) );
  AND2X2 U167 ( .A(a[3]), .B(b[7]), .Y(n131) );
  AND2X2 U168 ( .A(a[3]), .B(b[1]), .Y(n137) );
  AND2X1 U169 ( .A(a[6]), .B(b[2]), .Y(n112) );
  AND2X1 U170 ( .A(b[1]), .B(a[0]), .Y(n161) );
  AND2X1 U171 ( .A(b[3]), .B(a[0]), .Y(n159) );
  AND2X1 U172 ( .A(a[6]), .B(b[1]), .Y(n113) );
  AND2X1 U173 ( .A(b[2]), .B(a[0]), .Y(n160) );
  AND2X1 U174 ( .A(b[4]), .B(a[0]), .Y(n158) );
  AND2X1 U175 ( .A(a[4]), .B(b[0]), .Y(n130) );
  AND2X1 U176 ( .A(b[0]), .B(a[0]), .Y(product[0]) );
  AND2X1 U177 ( .A(a[6]), .B(b[0]), .Y(n114) );
  AND2X1 U178 ( .A(a[5]), .B(b[1]), .Y(n121) );
  AND2X1 U179 ( .A(a[6]), .B(b[3]), .Y(n111) );
  AND2X1 U180 ( .A(a[6]), .B(b[7]), .Y(n107) );
  AND2X1 U181 ( .A(a[4]), .B(b[4]), .Y(n126) );
  AND2X1 U182 ( .A(a[5]), .B(b[3]), .Y(n119) );
  AND2X1 U183 ( .A(a[6]), .B(b[4]), .Y(n110) );
  AND2X1 U184 ( .A(b[7]), .B(a[0]), .Y(n155) );
  AND2X1 U185 ( .A(a[5]), .B(b[2]), .Y(n120) );
  AND2X1 U186 ( .A(a[4]), .B(b[1]), .Y(n129) );
  AND2X1 U187 ( .A(a[5]), .B(b[0]), .Y(n122) );
  AND2X1 U188 ( .A(a[5]), .B(b[5]), .Y(n117) );
  AND2X1 U189 ( .A(b[5]), .B(a[0]), .Y(n157) );
  AND2X1 U190 ( .A(a[4]), .B(b[3]), .Y(n127) );
  AND2X1 U191 ( .A(a[5]), .B(b[7]), .Y(n115) );
  AND2X1 U192 ( .A(a[4]), .B(b[2]), .Y(n128) );
  AND2X1 U193 ( .A(a[4]), .B(b[5]), .Y(n125) );
  AND2X1 U194 ( .A(a[5]), .B(b[4]), .Y(n118) );
  AND2X1 U195 ( .A(a[6]), .B(b[5]), .Y(n109) );
  AND2X1 U196 ( .A(a[4]), .B(b[7]), .Y(n123) );
  AND2X1 U197 ( .A(b[7]), .B(a[7]), .Y(n99) );
  AND2X1 U198 ( .A(a[7]), .B(b[0]), .Y(n106) );
  AND2X1 U199 ( .A(b[1]), .B(a[7]), .Y(n105) );
  AND2X1 U200 ( .A(b[2]), .B(a[7]), .Y(n104) );
  AND2X1 U201 ( .A(b[3]), .B(a[7]), .Y(n103) );
  AND2X1 U202 ( .A(b[4]), .B(a[7]), .Y(n102) );
  AND2X1 U203 ( .A(b[5]), .B(a[7]), .Y(n101) );
endmodule


module alu_DW_mult_uns_4 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161;

  FAX1 U2 ( .A(n99), .B(n15), .C(n2), .YC(product[15]), .YS(product[14]) );
  FAX1 U3 ( .A(n16), .B(n17), .C(n3), .YC(n2), .YS(product[13]) );
  FAX1 U4 ( .A(n18), .B(n21), .C(n4), .YC(n3), .YS(product[12]) );
  FAX1 U5 ( .A(n22), .B(n27), .C(n5), .YC(n4), .YS(product[11]) );
  FAX1 U6 ( .A(n35), .B(n28), .C(n6), .YC(n5), .YS(product[10]) );
  FAX1 U7 ( .A(n45), .B(n36), .C(n7), .YC(n6), .YS(product[9]) );
  FAX1 U8 ( .A(n57), .B(n46), .C(n8), .YC(n7), .YS(product[8]) );
  FAX1 U9 ( .A(n69), .B(n58), .C(n9), .YC(n8), .YS(product[7]) );
  FAX1 U10 ( .A(n79), .B(n70), .C(n10), .YC(n9), .YS(product[6]) );
  FAX1 U11 ( .A(n87), .B(n80), .C(n11), .YC(n10), .YS(product[5]) );
  FAX1 U12 ( .A(n93), .B(n88), .C(n12), .YC(n11), .YS(product[4]) );
  FAX1 U13 ( .A(n96), .B(n94), .C(n13), .YC(n12), .YS(product[3]) );
  FAX1 U14 ( .A(n146), .B(n14), .C(n98), .YC(n13), .YS(product[2]) );
  HAX1 U15 ( .A(n154), .B(n161), .YC(n14), .YS(product[1]) );
  FAX1 U16 ( .A(n107), .B(n100), .C(n19), .YC(n15), .YS(n16) );
  FAX1 U17 ( .A(n25), .B(n20), .C(n23), .YC(n17), .YS(n18) );
  FAX1 U18 ( .A(n115), .B(n101), .C(n108), .YC(n19), .YS(n20) );
  FAX1 U19 ( .A(n31), .B(n24), .C(n29), .YC(n21), .YS(n22) );
  FAX1 U20 ( .A(n116), .B(n33), .C(n26), .YC(n23), .YS(n24) );
  FAX1 U21 ( .A(n123), .B(n102), .C(n109), .YC(n25), .YS(n26) );
  FAX1 U22 ( .A(n39), .B(n37), .C(n30), .YC(n27), .YS(n28) );
  FAX1 U23 ( .A(n41), .B(n34), .C(n32), .YC(n29), .YS(n30) );
  FAX1 U24 ( .A(n124), .B(n117), .C(n43), .YC(n31), .YS(n32) );
  FAX1 U25 ( .A(n131), .B(n103), .C(n110), .YC(n33), .YS(n34) );
  FAX1 U26 ( .A(n40), .B(n47), .C(n38), .YC(n35), .YS(n36) );
  FAX1 U27 ( .A(n44), .B(n51), .C(n49), .YC(n37), .YS(n38) );
  FAX1 U28 ( .A(n55), .B(n53), .C(n42), .YC(n39), .YS(n40) );
  FAX1 U29 ( .A(n118), .B(n125), .C(n132), .YC(n41), .YS(n42) );
  FAX1 U30 ( .A(n139), .B(n104), .C(n111), .YC(n43), .YS(n44) );
  FAX1 U31 ( .A(n50), .B(n59), .C(n48), .YC(n45), .YS(n46) );
  FAX1 U32 ( .A(n54), .B(n52), .C(n61), .YC(n47), .YS(n48) );
  FAX1 U33 ( .A(n56), .B(n65), .C(n63), .YC(n49), .YS(n50) );
  FAX1 U34 ( .A(n140), .B(n133), .C(n67), .YC(n51), .YS(n52) );
  FAX1 U35 ( .A(n126), .B(n119), .C(n147), .YC(n53), .YS(n54) );
  HAX1 U36 ( .A(n112), .B(n105), .YC(n55), .YS(n56) );
  FAX1 U37 ( .A(n62), .B(n71), .C(n60), .YC(n57), .YS(n58) );
  FAX1 U38 ( .A(n64), .B(n66), .C(n73), .YC(n59), .YS(n60) );
  FAX1 U39 ( .A(n77), .B(n68), .C(n75), .YC(n61), .YS(n62) );
  FAX1 U40 ( .A(n141), .B(n127), .C(n134), .YC(n63), .YS(n64) );
  FAX1 U41 ( .A(n155), .B(n120), .C(n148), .YC(n65), .YS(n66) );
  HAX1 U42 ( .A(n113), .B(n106), .YC(n67), .YS(n68) );
  FAX1 U43 ( .A(n74), .B(n81), .C(n72), .YC(n69), .YS(n70) );
  FAX1 U44 ( .A(n78), .B(n83), .C(n76), .YC(n71), .YS(n72) );
  FAX1 U45 ( .A(n142), .B(n135), .C(n85), .YC(n73), .YS(n74) );
  FAX1 U46 ( .A(n156), .B(n128), .C(n149), .YC(n75), .YS(n76) );
  HAX1 U47 ( .A(n121), .B(n114), .YC(n77), .YS(n78) );
  FAX1 U48 ( .A(n89), .B(n84), .C(n82), .YC(n79), .YS(n80) );
  FAX1 U49 ( .A(n150), .B(n91), .C(n86), .YC(n81), .YS(n82) );
  FAX1 U50 ( .A(n157), .B(n136), .C(n143), .YC(n83), .YS(n84) );
  HAX1 U51 ( .A(n129), .B(n122), .YC(n85), .YS(n86) );
  FAX1 U52 ( .A(n95), .B(n92), .C(n90), .YC(n87), .YS(n88) );
  FAX1 U53 ( .A(n158), .B(n144), .C(n151), .YC(n89), .YS(n90) );
  HAX1 U54 ( .A(n137), .B(n130), .YC(n91), .YS(n92) );
  FAX1 U55 ( .A(n159), .B(n152), .C(n97), .YC(n93), .YS(n94) );
  HAX1 U56 ( .A(n145), .B(n138), .YC(n95), .YS(n96) );
  HAX1 U57 ( .A(n160), .B(n153), .YC(n97), .YS(n98) );
  AND2X2 U140 ( .A(a[7]), .B(b[0]), .Y(n106) );
  AND2X2 U141 ( .A(a[6]), .B(b[0]), .Y(n114) );
  AND2X2 U142 ( .A(a[3]), .B(b[0]), .Y(n138) );
  AND2X2 U143 ( .A(a[4]), .B(b[0]), .Y(n130) );
  AND2X2 U144 ( .A(a[2]), .B(b[0]), .Y(n146) );
  AND2X2 U145 ( .A(a[1]), .B(b[0]), .Y(n154) );
  AND2X1 U146 ( .A(a[5]), .B(b[4]), .Y(n118) );
  AND2X1 U147 ( .A(a[4]), .B(b[4]), .Y(n126) );
  AND2X1 U148 ( .A(a[5]), .B(b[3]), .Y(n119) );
  AND2X1 U149 ( .A(b[1]), .B(a[7]), .Y(n105) );
  AND2X1 U150 ( .A(b[5]), .B(a[0]), .Y(n157) );
  AND2X1 U151 ( .A(a[3]), .B(b[4]), .Y(n134) );
  AND2X1 U152 ( .A(b[7]), .B(a[0]), .Y(n155) );
  AND2X1 U153 ( .A(a[5]), .B(b[2]), .Y(n120) );
  AND2X1 U154 ( .A(b[6]), .B(a[0]), .Y(n156) );
  AND2X1 U155 ( .A(a[5]), .B(b[1]), .Y(n121) );
  AND2X1 U156 ( .A(a[6]), .B(b[1]), .Y(n113) );
  AND2X1 U157 ( .A(a[5]), .B(b[5]), .Y(n117) );
  AND2X1 U158 ( .A(a[5]), .B(b[6]), .Y(n116) );
  AND2X1 U159 ( .A(a[2]), .B(b[4]), .Y(n142) );
  AND2X1 U160 ( .A(b[4]), .B(a[0]), .Y(n158) );
  AND2X1 U161 ( .A(a[3]), .B(b[1]), .Y(n137) );
  AND2X1 U162 ( .A(a[2]), .B(b[1]), .Y(n145) );
  AND2X1 U163 ( .A(a[5]), .B(b[7]), .Y(n115) );
  AND2X1 U164 ( .A(b[3]), .B(a[0]), .Y(n159) );
  AND2X1 U165 ( .A(b[1]), .B(a[0]), .Y(n161) );
  AND2X2 U166 ( .A(a[4]), .B(b[1]), .Y(n129) );
  AND2X2 U167 ( .A(a[1]), .B(b[1]), .Y(n153) );
  AND2X2 U168 ( .A(b[0]), .B(a[0]), .Y(product[0]) );
  AND2X2 U169 ( .A(b[2]), .B(a[0]), .Y(n160) );
  AND2X2 U170 ( .A(a[5]), .B(b[0]), .Y(n122) );
  AND2X2 U171 ( .A(b[4]), .B(a[7]), .Y(n102) );
  AND2X2 U172 ( .A(a[6]), .B(b[4]), .Y(n110) );
  AND2X2 U173 ( .A(a[1]), .B(b[4]), .Y(n150) );
  AND2X1 U174 ( .A(a[3]), .B(b[3]), .Y(n135) );
  AND2X1 U175 ( .A(a[3]), .B(b[6]), .Y(n132) );
  AND2X1 U176 ( .A(a[3]), .B(b[5]), .Y(n133) );
  AND2X1 U177 ( .A(a[3]), .B(b[7]), .Y(n131) );
  AND2X1 U178 ( .A(a[3]), .B(b[2]), .Y(n136) );
  AND2X1 U179 ( .A(b[7]), .B(a[7]), .Y(n99) );
  AND2X1 U180 ( .A(a[1]), .B(b[2]), .Y(n152) );
  AND2X1 U181 ( .A(a[1]), .B(b[3]), .Y(n151) );
  AND2X1 U182 ( .A(a[1]), .B(b[5]), .Y(n149) );
  AND2X1 U183 ( .A(a[1]), .B(b[6]), .Y(n148) );
  AND2X1 U184 ( .A(a[1]), .B(b[7]), .Y(n147) );
  AND2X1 U185 ( .A(a[2]), .B(b[2]), .Y(n144) );
  AND2X1 U186 ( .A(a[2]), .B(b[3]), .Y(n143) );
  AND2X1 U187 ( .A(a[2]), .B(b[5]), .Y(n141) );
  AND2X1 U188 ( .A(a[2]), .B(b[6]), .Y(n140) );
  AND2X1 U189 ( .A(a[2]), .B(b[7]), .Y(n139) );
  AND2X1 U190 ( .A(a[4]), .B(b[2]), .Y(n128) );
  AND2X1 U191 ( .A(a[4]), .B(b[3]), .Y(n127) );
  AND2X1 U192 ( .A(a[4]), .B(b[5]), .Y(n125) );
  AND2X1 U193 ( .A(a[4]), .B(b[6]), .Y(n124) );
  AND2X1 U194 ( .A(a[4]), .B(b[7]), .Y(n123) );
  AND2X1 U195 ( .A(a[6]), .B(b[2]), .Y(n112) );
  AND2X1 U196 ( .A(a[6]), .B(b[3]), .Y(n111) );
  AND2X1 U197 ( .A(a[6]), .B(b[5]), .Y(n109) );
  AND2X1 U198 ( .A(a[6]), .B(b[6]), .Y(n108) );
  AND2X1 U199 ( .A(a[6]), .B(b[7]), .Y(n107) );
  AND2X1 U200 ( .A(b[2]), .B(a[7]), .Y(n104) );
  AND2X1 U201 ( .A(b[3]), .B(a[7]), .Y(n103) );
  AND2X1 U202 ( .A(b[5]), .B(a[7]), .Y(n101) );
  AND2X1 U203 ( .A(b[6]), .B(a[7]), .Y(n100) );
endmodule


module alu_DW_mult_uns_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161;

  FAX1 U2 ( .A(n99), .B(n15), .C(n2), .YC(product[15]), .YS(product[14]) );
  FAX1 U3 ( .A(n16), .B(n17), .C(n3), .YC(n2), .YS(product[13]) );
  FAX1 U4 ( .A(n18), .B(n21), .C(n4), .YC(n3), .YS(product[12]) );
  FAX1 U5 ( .A(n22), .B(n27), .C(n5), .YC(n4), .YS(product[11]) );
  FAX1 U6 ( .A(n35), .B(n28), .C(n6), .YC(n5), .YS(product[10]) );
  FAX1 U7 ( .A(n45), .B(n36), .C(n7), .YC(n6), .YS(product[9]) );
  FAX1 U8 ( .A(n57), .B(n46), .C(n8), .YC(n7), .YS(product[8]) );
  FAX1 U9 ( .A(n69), .B(n58), .C(n9), .YC(n8), .YS(product[7]) );
  FAX1 U10 ( .A(n79), .B(n70), .C(n10), .YC(n9), .YS(product[6]) );
  FAX1 U11 ( .A(n87), .B(n80), .C(n11), .YC(n10), .YS(product[5]) );
  FAX1 U12 ( .A(n93), .B(n88), .C(n12), .YC(n11), .YS(product[4]) );
  FAX1 U13 ( .A(n96), .B(n94), .C(n13), .YC(n12), .YS(product[3]) );
  FAX1 U14 ( .A(n146), .B(n14), .C(n98), .YC(n13), .YS(product[2]) );
  HAX1 U15 ( .A(n154), .B(n161), .YC(n14), .YS(product[1]) );
  FAX1 U16 ( .A(n107), .B(n100), .C(n19), .YC(n15), .YS(n16) );
  FAX1 U17 ( .A(n25), .B(n20), .C(n23), .YC(n17), .YS(n18) );
  FAX1 U18 ( .A(n115), .B(n101), .C(n108), .YC(n19), .YS(n20) );
  FAX1 U19 ( .A(n31), .B(n24), .C(n29), .YC(n21), .YS(n22) );
  FAX1 U20 ( .A(n116), .B(n33), .C(n26), .YC(n23), .YS(n24) );
  FAX1 U21 ( .A(n123), .B(n102), .C(n109), .YC(n25), .YS(n26) );
  FAX1 U22 ( .A(n39), .B(n37), .C(n30), .YC(n27), .YS(n28) );
  FAX1 U23 ( .A(n41), .B(n34), .C(n32), .YC(n29), .YS(n30) );
  FAX1 U24 ( .A(n124), .B(n117), .C(n43), .YC(n31), .YS(n32) );
  FAX1 U25 ( .A(n131), .B(n103), .C(n110), .YC(n33), .YS(n34) );
  FAX1 U26 ( .A(n40), .B(n47), .C(n38), .YC(n35), .YS(n36) );
  FAX1 U27 ( .A(n44), .B(n51), .C(n49), .YC(n37), .YS(n38) );
  FAX1 U28 ( .A(n55), .B(n53), .C(n42), .YC(n39), .YS(n40) );
  FAX1 U29 ( .A(n118), .B(n125), .C(n132), .YC(n41), .YS(n42) );
  FAX1 U30 ( .A(n139), .B(n104), .C(n111), .YC(n43), .YS(n44) );
  FAX1 U31 ( .A(n50), .B(n59), .C(n48), .YC(n45), .YS(n46) );
  FAX1 U32 ( .A(n54), .B(n52), .C(n61), .YC(n47), .YS(n48) );
  FAX1 U33 ( .A(n56), .B(n65), .C(n63), .YC(n49), .YS(n50) );
  FAX1 U34 ( .A(n140), .B(n133), .C(n67), .YC(n51), .YS(n52) );
  FAX1 U35 ( .A(n126), .B(n119), .C(n147), .YC(n53), .YS(n54) );
  HAX1 U36 ( .A(n112), .B(n105), .YC(n55), .YS(n56) );
  FAX1 U37 ( .A(n62), .B(n71), .C(n60), .YC(n57), .YS(n58) );
  FAX1 U38 ( .A(n64), .B(n66), .C(n73), .YC(n59), .YS(n60) );
  FAX1 U39 ( .A(n77), .B(n68), .C(n75), .YC(n61), .YS(n62) );
  FAX1 U40 ( .A(n141), .B(n127), .C(n134), .YC(n63), .YS(n64) );
  FAX1 U41 ( .A(n155), .B(n120), .C(n148), .YC(n65), .YS(n66) );
  HAX1 U42 ( .A(n113), .B(n106), .YC(n67), .YS(n68) );
  FAX1 U43 ( .A(n74), .B(n81), .C(n72), .YC(n69), .YS(n70) );
  FAX1 U44 ( .A(n78), .B(n83), .C(n76), .YC(n71), .YS(n72) );
  FAX1 U45 ( .A(n142), .B(n135), .C(n85), .YC(n73), .YS(n74) );
  FAX1 U46 ( .A(n156), .B(n128), .C(n149), .YC(n75), .YS(n76) );
  HAX1 U47 ( .A(n121), .B(n114), .YC(n77), .YS(n78) );
  FAX1 U48 ( .A(n89), .B(n84), .C(n82), .YC(n79), .YS(n80) );
  FAX1 U49 ( .A(n150), .B(n91), .C(n86), .YC(n81), .YS(n82) );
  FAX1 U50 ( .A(n157), .B(n136), .C(n143), .YC(n83), .YS(n84) );
  HAX1 U51 ( .A(n129), .B(n122), .YC(n85), .YS(n86) );
  FAX1 U52 ( .A(n95), .B(n92), .C(n90), .YC(n87), .YS(n88) );
  FAX1 U53 ( .A(n158), .B(n144), .C(n151), .YC(n89), .YS(n90) );
  HAX1 U54 ( .A(n137), .B(n130), .YC(n91), .YS(n92) );
  FAX1 U55 ( .A(n159), .B(n152), .C(n97), .YC(n93), .YS(n94) );
  HAX1 U56 ( .A(n145), .B(n138), .YC(n95), .YS(n96) );
  HAX1 U57 ( .A(n160), .B(n153), .YC(n97), .YS(n98) );
  AND2X2 U140 ( .A(b[5]), .B(a[0]), .Y(n157) );
  AND2X2 U141 ( .A(a[5]), .B(b[0]), .Y(n122) );
  AND2X2 U142 ( .A(a[5]), .B(b[1]), .Y(n121) );
  AND2X2 U143 ( .A(a[5]), .B(b[6]), .Y(n116) );
  AND2X2 U144 ( .A(a[5]), .B(b[2]), .Y(n120) );
  AND2X2 U145 ( .A(a[5]), .B(b[5]), .Y(n117) );
  AND2X2 U146 ( .A(a[5]), .B(b[3]), .Y(n119) );
  AND2X1 U147 ( .A(a[6]), .B(b[6]), .Y(n108) );
  AND2X1 U148 ( .A(a[6]), .B(b[3]), .Y(n111) );
  AND2X1 U149 ( .A(b[6]), .B(a[7]), .Y(n100) );
  AND2X1 U150 ( .A(a[4]), .B(b[5]), .Y(n125) );
  AND2X1 U151 ( .A(a[3]), .B(b[6]), .Y(n132) );
  AND2X1 U152 ( .A(a[1]), .B(b[7]), .Y(n147) );
  AND2X1 U153 ( .A(a[6]), .B(b[2]), .Y(n112) );
  AND2X1 U154 ( .A(b[1]), .B(a[7]), .Y(n105) );
  AND2X1 U155 ( .A(a[4]), .B(b[6]), .Y(n124) );
  AND2X1 U156 ( .A(a[2]), .B(b[5]), .Y(n141) );
  AND2X1 U157 ( .A(a[4]), .B(b[3]), .Y(n127) );
  AND2X1 U158 ( .A(b[7]), .B(a[0]), .Y(n155) );
  AND2X1 U159 ( .A(a[1]), .B(b[6]), .Y(n148) );
  AND2X1 U160 ( .A(a[7]), .B(b[0]), .Y(n106) );
  AND2X1 U161 ( .A(a[6]), .B(b[1]), .Y(n113) );
  AND2X1 U162 ( .A(a[3]), .B(b[1]), .Y(n137) );
  AND2X1 U163 ( .A(a[4]), .B(b[0]), .Y(n130) );
  AND2X1 U164 ( .A(a[1]), .B(b[5]), .Y(n149) );
  AND2X1 U165 ( .A(a[4]), .B(b[2]), .Y(n128) );
  AND2X1 U166 ( .A(b[6]), .B(a[0]), .Y(n156) );
  AND2X1 U167 ( .A(a[6]), .B(b[0]), .Y(n114) );
  AND2X1 U168 ( .A(a[4]), .B(b[1]), .Y(n129) );
  AND2X1 U169 ( .A(b[3]), .B(a[0]), .Y(n159) );
  AND2X1 U170 ( .A(a[1]), .B(b[2]), .Y(n152) );
  AND2X1 U171 ( .A(a[2]), .B(b[1]), .Y(n145) );
  AND2X1 U172 ( .A(a[3]), .B(b[0]), .Y(n138) );
  AND2X1 U173 ( .A(a[1]), .B(b[3]), .Y(n151) );
  AND2X1 U174 ( .A(b[7]), .B(a[7]), .Y(n99) );
  AND2X1 U175 ( .A(a[2]), .B(b[0]), .Y(n146) );
  AND2X2 U176 ( .A(a[3]), .B(b[7]), .Y(n131) );
  AND2X2 U177 ( .A(a[2]), .B(b[7]), .Y(n139) );
  AND2X2 U178 ( .A(a[1]), .B(b[0]), .Y(n154) );
  AND2X2 U179 ( .A(a[4]), .B(b[7]), .Y(n123) );
  AND2X2 U180 ( .A(b[0]), .B(a[0]), .Y(product[0]) );
  AND2X2 U181 ( .A(b[2]), .B(a[0]), .Y(n160) );
  AND2X2 U182 ( .A(b[4]), .B(a[7]), .Y(n102) );
  AND2X2 U183 ( .A(a[4]), .B(b[4]), .Y(n126) );
  AND2X2 U184 ( .A(a[3]), .B(b[4]), .Y(n134) );
  AND2X2 U185 ( .A(a[2]), .B(b[4]), .Y(n142) );
  AND2X2 U186 ( .A(a[1]), .B(b[4]), .Y(n150) );
  AND2X2 U187 ( .A(b[4]), .B(a[0]), .Y(n158) );
  AND2X2 U188 ( .A(b[5]), .B(a[7]), .Y(n101) );
  AND2X2 U189 ( .A(a[3]), .B(b[5]), .Y(n133) );
  AND2X2 U190 ( .A(a[5]), .B(b[7]), .Y(n115) );
  AND2X2 U191 ( .A(a[5]), .B(b[4]), .Y(n118) );
  AND2X2 U192 ( .A(a[6]), .B(b[7]), .Y(n107) );
  AND2X2 U193 ( .A(a[6]), .B(b[5]), .Y(n109) );
  AND2X2 U194 ( .A(a[6]), .B(b[4]), .Y(n110) );
  AND2X2 U195 ( .A(a[2]), .B(b[6]), .Y(n140) );
  AND2X2 U196 ( .A(b[1]), .B(a[0]), .Y(n161) );
  AND2X2 U197 ( .A(a[1]), .B(b[1]), .Y(n153) );
  AND2X1 U198 ( .A(a[3]), .B(b[3]), .Y(n135) );
  AND2X1 U199 ( .A(a[3]), .B(b[2]), .Y(n136) );
  AND2X1 U200 ( .A(b[3]), .B(a[7]), .Y(n103) );
  AND2X1 U201 ( .A(b[2]), .B(a[7]), .Y(n104) );
  AND2X1 U202 ( .A(a[2]), .B(b[2]), .Y(n144) );
  AND2X1 U203 ( .A(a[2]), .B(b[3]), .Y(n143) );
endmodule


module alu_DW_mult_uns_2 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n214, n215;

  FAX1 U2 ( .A(n99), .B(n15), .C(n2), .YC(product[15]), .YS(product[14]) );
  FAX1 U3 ( .A(n16), .B(n17), .C(n3), .YC(n2), .YS(product[13]) );
  FAX1 U4 ( .A(n18), .B(n21), .C(n4), .YC(n3), .YS(product[12]) );
  FAX1 U5 ( .A(n22), .B(n27), .C(n5), .YC(n4), .YS(product[11]) );
  FAX1 U6 ( .A(n35), .B(n28), .C(n6), .YC(n5), .YS(product[10]) );
  FAX1 U7 ( .A(n45), .B(n36), .C(n7), .YC(n6), .YS(product[9]) );
  FAX1 U8 ( .A(n57), .B(n46), .C(n8), .YC(n7), .YS(product[8]) );
  FAX1 U9 ( .A(n69), .B(n58), .C(n9), .YC(n8), .YS(product[7]) );
  FAX1 U10 ( .A(n79), .B(n70), .C(n10), .YC(n9), .YS(product[6]) );
  FAX1 U11 ( .A(n87), .B(n80), .C(n11), .YC(n10), .YS(product[5]) );
  FAX1 U12 ( .A(n93), .B(n88), .C(n12), .YC(n11), .YS(product[4]) );
  FAX1 U13 ( .A(n96), .B(n13), .C(n94), .YC(n12), .YS(product[3]) );
  FAX1 U14 ( .A(n146), .B(n14), .C(n98), .YC(n13), .YS(product[2]) );
  HAX1 U15 ( .A(n154), .B(n161), .YC(n14), .YS(product[1]) );
  FAX1 U16 ( .A(n107), .B(n100), .C(n19), .YC(n15), .YS(n16) );
  FAX1 U17 ( .A(n25), .B(n20), .C(n23), .YC(n17), .YS(n18) );
  FAX1 U18 ( .A(n115), .B(n101), .C(n108), .YC(n19), .YS(n20) );
  FAX1 U19 ( .A(n31), .B(n24), .C(n29), .YC(n21), .YS(n22) );
  FAX1 U20 ( .A(n116), .B(n33), .C(n26), .YC(n23), .YS(n24) );
  FAX1 U21 ( .A(n123), .B(n102), .C(n109), .YC(n25), .YS(n26) );
  FAX1 U22 ( .A(n39), .B(n37), .C(n30), .YC(n27), .YS(n28) );
  FAX1 U23 ( .A(n41), .B(n34), .C(n32), .YC(n29), .YS(n30) );
  FAX1 U24 ( .A(n124), .B(n117), .C(n43), .YC(n31), .YS(n32) );
  FAX1 U25 ( .A(n131), .B(n103), .C(n110), .YC(n33), .YS(n34) );
  FAX1 U26 ( .A(n40), .B(n47), .C(n38), .YC(n35), .YS(n36) );
  FAX1 U27 ( .A(n44), .B(n51), .C(n49), .YC(n37), .YS(n38) );
  FAX1 U28 ( .A(n55), .B(n53), .C(n42), .YC(n39), .YS(n40) );
  FAX1 U29 ( .A(n118), .B(n125), .C(n132), .YC(n41), .YS(n42) );
  FAX1 U30 ( .A(n139), .B(n104), .C(n111), .YC(n43), .YS(n44) );
  FAX1 U31 ( .A(n50), .B(n59), .C(n48), .YC(n45), .YS(n46) );
  FAX1 U32 ( .A(n54), .B(n52), .C(n61), .YC(n47), .YS(n48) );
  FAX1 U33 ( .A(n56), .B(n65), .C(n63), .YC(n49), .YS(n50) );
  FAX1 U34 ( .A(n140), .B(n133), .C(n67), .YC(n51), .YS(n52) );
  FAX1 U35 ( .A(n126), .B(n119), .C(n147), .YC(n53), .YS(n54) );
  HAX1 U36 ( .A(n112), .B(n105), .YC(n55), .YS(n56) );
  FAX1 U37 ( .A(n62), .B(n71), .C(n60), .YC(n57), .YS(n58) );
  FAX1 U38 ( .A(n64), .B(n66), .C(n73), .YC(n59), .YS(n60) );
  FAX1 U39 ( .A(n77), .B(n68), .C(n75), .YC(n61), .YS(n62) );
  FAX1 U40 ( .A(n141), .B(n127), .C(n134), .YC(n63), .YS(n64) );
  FAX1 U41 ( .A(n155), .B(n120), .C(n148), .YC(n65), .YS(n66) );
  HAX1 U42 ( .A(n113), .B(n106), .YC(n67), .YS(n68) );
  FAX1 U43 ( .A(n74), .B(n81), .C(n72), .YC(n69), .YS(n70) );
  FAX1 U44 ( .A(n78), .B(n83), .C(n76), .YC(n71), .YS(n72) );
  FAX1 U45 ( .A(n142), .B(n135), .C(n85), .YC(n73), .YS(n74) );
  FAX1 U46 ( .A(n156), .B(n128), .C(n149), .YC(n75), .YS(n76) );
  HAX1 U47 ( .A(n121), .B(n114), .YC(n77), .YS(n78) );
  FAX1 U48 ( .A(n89), .B(n84), .C(n82), .YC(n79), .YS(n80) );
  FAX1 U49 ( .A(n150), .B(n91), .C(n86), .YC(n81), .YS(n82) );
  FAX1 U50 ( .A(n157), .B(n136), .C(n143), .YC(n83), .YS(n84) );
  HAX1 U51 ( .A(n129), .B(n122), .YC(n85), .YS(n86) );
  FAX1 U52 ( .A(n95), .B(n92), .C(n90), .YC(n87), .YS(n88) );
  FAX1 U53 ( .A(n158), .B(n144), .C(n151), .YC(n89), .YS(n90) );
  HAX1 U54 ( .A(n137), .B(n130), .YC(n91), .YS(n92) );
  FAX1 U55 ( .A(n159), .B(n152), .C(n97), .YC(n93), .YS(n94) );
  HAX1 U56 ( .A(n145), .B(n138), .YC(n95), .YS(n96) );
  HAX1 U57 ( .A(n153), .B(n160), .YC(n97), .YS(n98) );
  BUFX2 U140 ( .A(a[0]), .Y(n214) );
  AND2X1 U141 ( .A(a[5]), .B(b[7]), .Y(n115) );
  AND2X1 U142 ( .A(a[5]), .B(b[0]), .Y(n122) );
  AND2X1 U143 ( .A(a[6]), .B(b[7]), .Y(n107) );
  AND2X1 U144 ( .A(b[0]), .B(n215), .Y(product[0]) );
  AND2X1 U145 ( .A(b[3]), .B(a[7]), .Y(n103) );
  AND2X1 U146 ( .A(a[3]), .B(b[7]), .Y(n131) );
  AND2X1 U147 ( .A(a[6]), .B(b[4]), .Y(n110) );
  AND2X1 U148 ( .A(a[2]), .B(b[7]), .Y(n139) );
  AND2X1 U149 ( .A(b[2]), .B(a[7]), .Y(n104) );
  AND2X1 U150 ( .A(a[6]), .B(b[3]), .Y(n111) );
  AND2X1 U151 ( .A(a[1]), .B(b[7]), .Y(n147) );
  AND2X1 U152 ( .A(a[5]), .B(b[3]), .Y(n119) );
  AND2X1 U153 ( .A(b[1]), .B(a[7]), .Y(n105) );
  AND2X1 U154 ( .A(a[6]), .B(b[2]), .Y(n112) );
  AND2X1 U155 ( .A(a[4]), .B(b[7]), .Y(n123) );
  AND2X1 U156 ( .A(b[4]), .B(a[7]), .Y(n102) );
  AND2X1 U157 ( .A(a[6]), .B(b[5]), .Y(n109) );
  AND2X1 U158 ( .A(a[7]), .B(b[0]), .Y(n106) );
  AND2X1 U159 ( .A(a[6]), .B(b[1]), .Y(n113) );
  AND2X1 U160 ( .A(a[5]), .B(b[2]), .Y(n120) );
  AND2X1 U161 ( .A(b[7]), .B(n215), .Y(n155) );
  AND2X1 U162 ( .A(a[4]), .B(b[3]), .Y(n127) );
  AND2X1 U163 ( .A(a[5]), .B(b[1]), .Y(n121) );
  AND2X1 U164 ( .A(a[6]), .B(b[0]), .Y(n114) );
  AND2X1 U165 ( .A(a[4]), .B(b[2]), .Y(n128) );
  AND2X1 U166 ( .A(a[2]), .B(b[3]), .Y(n143) );
  AND2X1 U167 ( .A(a[3]), .B(b[2]), .Y(n136) );
  AND2X1 U168 ( .A(a[2]), .B(b[2]), .Y(n144) );
  AND2X1 U169 ( .A(a[1]), .B(b[3]), .Y(n151) );
  AND2X1 U170 ( .A(b[4]), .B(a[0]), .Y(n158) );
  AND2X1 U171 ( .A(a[4]), .B(b[0]), .Y(n130) );
  AND2X1 U172 ( .A(a[3]), .B(b[1]), .Y(n137) );
  AND2X1 U173 ( .A(a[3]), .B(b[3]), .Y(n135) );
  AND2X1 U174 ( .A(a[2]), .B(b[1]), .Y(n145) );
  AND2X1 U175 ( .A(a[3]), .B(b[0]), .Y(n138) );
  AND2X1 U176 ( .A(a[1]), .B(b[1]), .Y(n153) );
  AND2X1 U177 ( .A(b[2]), .B(a[0]), .Y(n160) );
  AND2X1 U178 ( .A(b[7]), .B(a[7]), .Y(n99) );
  AND2X1 U179 ( .A(a[1]), .B(b[0]), .Y(n154) );
  AND2X1 U180 ( .A(b[1]), .B(n214), .Y(n161) );
  AND2X2 U181 ( .A(a[1]), .B(b[2]), .Y(n152) );
  AND2X2 U182 ( .A(a[6]), .B(b[6]), .Y(n108) );
  BUFX2 U183 ( .A(n214), .Y(n215) );
  AND2X2 U184 ( .A(b[3]), .B(n214), .Y(n159) );
  AND2X2 U185 ( .A(b[6]), .B(a[7]), .Y(n100) );
  AND2X2 U186 ( .A(b[5]), .B(a[7]), .Y(n101) );
  AND2X2 U187 ( .A(a[2]), .B(b[0]), .Y(n146) );
  AND2X2 U188 ( .A(a[4]), .B(b[1]), .Y(n129) );
  AND2X1 U189 ( .A(a[3]), .B(b[5]), .Y(n133) );
  AND2X1 U190 ( .A(b[5]), .B(n214), .Y(n157) );
  AND2X1 U191 ( .A(a[5]), .B(b[6]), .Y(n116) );
  AND2X1 U192 ( .A(a[3]), .B(b[4]), .Y(n134) );
  AND2X1 U193 ( .A(b[6]), .B(n214), .Y(n156) );
  AND2X1 U194 ( .A(a[3]), .B(b[6]), .Y(n132) );
  AND2X1 U195 ( .A(a[5]), .B(b[4]), .Y(n118) );
  AND2X1 U196 ( .A(a[5]), .B(b[5]), .Y(n117) );
  AND2X1 U197 ( .A(a[1]), .B(b[4]), .Y(n150) );
  AND2X1 U198 ( .A(a[1]), .B(b[5]), .Y(n149) );
  AND2X1 U199 ( .A(a[1]), .B(b[6]), .Y(n148) );
  AND2X1 U200 ( .A(a[2]), .B(b[4]), .Y(n142) );
  AND2X1 U201 ( .A(a[2]), .B(b[5]), .Y(n141) );
  AND2X1 U202 ( .A(a[2]), .B(b[6]), .Y(n140) );
  AND2X1 U203 ( .A(a[4]), .B(b[4]), .Y(n126) );
  AND2X1 U204 ( .A(a[4]), .B(b[5]), .Y(n125) );
  AND2X1 U205 ( .A(a[4]), .B(b[6]), .Y(n124) );
endmodule


module alu_DW01_sub_15 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n67, n68, n69, n73, n74, n75, n76, n77, n81,
         n82, n83, n84, n85, n89, n90, n91, n92, n93, n97, n98, n99, n100,
         n101, n105, n106, n107, n108, n109, n113, n114, n115, n116, n117,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n143, n144, n146,
         n147, n148, n149, n150, n151, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n171, n172,
         n173, n175, n176, n177, n178, n179, n180, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n196, n197, n198, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n309, n310, n311, n313, n314, n315, n316, n317, n318,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n334, n335, n336, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n399, n402, n404, n406, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053;

  XOR2X1 U1 ( .A(n61), .B(n1), .Y(DIFF[63]) );
  FAX1 U3 ( .A(n1053), .B(A[62]), .C(n62), .YC(n61), .YS(DIFF[62]) );
  FAX1 U4 ( .A(n1052), .B(A[61]), .C(n381), .YC(n62), .YS(DIFF[61]) );
  XNOR2X1 U6 ( .A(n68), .B(n961), .Y(DIFF[60]) );
  AOI21X1 U7 ( .A(n68), .B(n989), .C(n67), .Y(n63) );
  FAX1 U14 ( .A(n1050), .B(A[59]), .C(n382), .YC(n68), .YS(DIFF[59]) );
  XNOR2X1 U16 ( .A(n980), .B(n962), .Y(DIFF[58]) );
  AOI21X1 U17 ( .A(n74), .B(n985), .C(n73), .Y(n69) );
  XOR2X1 U24 ( .A(n719), .B(n791), .Y(DIFF[57]) );
  OAI21X1 U25 ( .A(n737), .B(n875), .C(n824), .Y(n74) );
  XNOR2X1 U30 ( .A(n718), .B(n943), .Y(DIFF[56]) );
  AOI21X1 U31 ( .A(n82), .B(n984), .C(n81), .Y(n77) );
  XOR2X1 U38 ( .A(n873), .B(n790), .Y(DIFF[55]) );
  OAI21X1 U39 ( .A(n825), .B(n873), .C(n823), .Y(n82) );
  XNOR2X1 U44 ( .A(n713), .B(n773), .Y(DIFF[54]) );
  AOI21X1 U45 ( .A(n90), .B(n983), .C(n89), .Y(n85) );
  XOR2X1 U52 ( .A(n716), .B(n789), .Y(DIFF[53]) );
  OAI21X1 U53 ( .A(n736), .B(n871), .C(n822), .Y(n90) );
  XNOR2X1 U58 ( .A(n712), .B(n921), .Y(DIFF[52]) );
  AOI21X1 U59 ( .A(n98), .B(n990), .C(n97), .Y(n93) );
  XOR2X1 U66 ( .A(n869), .B(n788), .Y(DIFF[51]) );
  OAI21X1 U67 ( .A(n735), .B(n738), .C(n821), .Y(n98) );
  XNOR2X1 U72 ( .A(n706), .B(n772), .Y(DIFF[50]) );
  AOI21X1 U73 ( .A(n106), .B(n988), .C(n105), .Y(n101) );
  XOR2X1 U80 ( .A(n867), .B(n787), .Y(DIFF[49]) );
  OAI21X1 U81 ( .A(n734), .B(n868), .C(n820), .Y(n106) );
  XNOR2X1 U86 ( .A(n979), .B(n771), .Y(DIFF[48]) );
  AOI21X1 U87 ( .A(n114), .B(n986), .C(n113), .Y(n109) );
  XOR2X1 U94 ( .A(n864), .B(n786), .Y(DIFF[47]) );
  OAI21X1 U95 ( .A(n733), .B(n865), .C(n819), .Y(n114) );
  XNOR2X1 U100 ( .A(n705), .B(n770), .Y(DIFF[46]) );
  AOI21X1 U101 ( .A(n122), .B(n982), .C(n121), .Y(n117) );
  XOR2X1 U108 ( .A(n861), .B(n785), .Y(DIFF[45]) );
  OAI21X1 U109 ( .A(n732), .B(n862), .C(n818), .Y(n122) );
  XNOR2X1 U114 ( .A(n130), .B(n769), .Y(DIFF[44]) );
  AOI21X1 U115 ( .A(n209), .B(n728), .C(n127), .Y(n125) );
  OAI21X1 U117 ( .A(n884), .B(n731), .C(n817), .Y(n127) );
  XNOR2X1 U122 ( .A(n137), .B(n768), .Y(DIFF[43]) );
  OAI21X1 U123 ( .A(n852), .B(n208), .C(n708), .Y(n130) );
  AOI21X1 U125 ( .A(n161), .B(n715), .C(n134), .Y(n132) );
  OAI21X1 U127 ( .A(n883), .B(n849), .C(n816), .Y(n134) );
  XNOR2X1 U132 ( .A(n144), .B(n901), .Y(DIFF[42]) );
  OAI21X1 U133 ( .A(n726), .B(n156), .C(n849), .Y(n137) );
  AOI21X1 U135 ( .A(n148), .B(n987), .C(n143), .Y(n139) );
  XOR2X1 U142 ( .A(n904), .B(n903), .Y(DIFF[41]) );
  OAI21X1 U143 ( .A(n147), .B(n156), .C(n146), .Y(n144) );
  OAI21X1 U147 ( .A(n954), .B(n973), .C(n938), .Y(n148) );
  XOR2X1 U152 ( .A(n156), .B(n913), .Y(DIFF[40]) );
  AOI21X1 U153 ( .A(n157), .B(n402), .C(n155), .Y(n151) );
  XOR2X1 U160 ( .A(n753), .B(n784), .Y(DIFF[39]) );
  OAI21X1 U162 ( .A(n158), .B(n208), .C(n159), .Y(n157) );
  OAI21X1 U166 ( .A(n717), .B(n847), .C(n747), .Y(n161) );
  AOI21X1 U168 ( .A(n177), .B(n842), .C(n165), .Y(n163) );
  OAI21X1 U170 ( .A(n953), .B(n972), .C(n815), .Y(n165) );
  XNOR2X1 U175 ( .A(n173), .B(n922), .Y(DIFF[38]) );
  AOI21X1 U176 ( .A(n173), .B(n404), .C(n172), .Y(n168) );
  XOR2X1 U183 ( .A(n752), .B(n783), .Y(DIFF[37]) );
  OAI21X1 U184 ( .A(n176), .B(n185), .C(n175), .Y(n173) );
  OAI21X1 U188 ( .A(n949), .B(n978), .C(n936), .Y(n177) );
  XOR2X1 U193 ( .A(n185), .B(n912), .Y(DIFF[36]) );
  AOI21X1 U194 ( .A(n186), .B(n406), .C(n184), .Y(n180) );
  XOR2X1 U201 ( .A(n751), .B(n782), .Y(DIFF[35]) );
  OAI21X1 U203 ( .A(n851), .B(n208), .C(n707), .Y(n186) );
  AOI21X1 U205 ( .A(n835), .B(n202), .C(n190), .Y(n188) );
  OAI21X1 U207 ( .A(n952), .B(n714), .C(n814), .Y(n190) );
  XNOR2X1 U212 ( .A(n198), .B(n909), .Y(DIFF[34]) );
  AOI21X1 U213 ( .A(n198), .B(n196), .C(n197), .Y(n193) );
  XNOR2X1 U220 ( .A(n205), .B(n902), .Y(DIFF[33]) );
  OAI21X1 U221 ( .A(n792), .B(n208), .C(n200), .Y(n198) );
  OAI21X1 U225 ( .A(n960), .B(n941), .C(n803), .Y(n202) );
  XOR2X1 U230 ( .A(n208), .B(n924), .Y(DIFF[32]) );
  OAI21X1 U231 ( .A(n964), .B(n208), .C(n960), .Y(n205) );
  XNOR2X1 U236 ( .A(n220), .B(n767), .Y(DIFF[31]) );
  OAI21X1 U238 ( .A(n729), .B(n739), .C(n746), .Y(n209) );
  AOI21X1 U240 ( .A(n255), .B(n725), .C(n213), .Y(n211) );
  OAI21X1 U242 ( .A(n854), .B(n831), .C(n744), .Y(n213) );
  AOI21X1 U244 ( .A(n225), .B(n724), .C(n217), .Y(n215) );
  OAI21X1 U246 ( .A(n893), .B(n879), .C(n813), .Y(n217) );
  XOR2X1 U251 ( .A(n859), .B(n781), .Y(DIFF[30]) );
  OAI21X1 U252 ( .A(n882), .B(n859), .C(n893), .Y(n220) );
  XNOR2X1 U257 ( .A(n228), .B(n766), .Y(DIFF[29]) );
  AOI21X1 U258 ( .A(n231), .B(n834), .C(n225), .Y(n223) );
  OAI21X1 U260 ( .A(n892), .B(n956), .C(n812), .Y(n225) );
  XNOR2X1 U265 ( .A(n231), .B(n765), .Y(DIFF[28]) );
  OAI21X1 U266 ( .A(n975), .B(n832), .C(n892), .Y(n228) );
  XNOR2X1 U271 ( .A(n241), .B(n764), .Y(DIFF[27]) );
  AOI21X1 U273 ( .A(n252), .B(n233), .C(n830), .Y(n232) );
  AOI21X1 U277 ( .A(n246), .B(n841), .C(n238), .Y(n236) );
  OAI21X1 U279 ( .A(n891), .B(n977), .C(n811), .Y(n238) );
  XOR2X1 U284 ( .A(n858), .B(n780), .Y(DIFF[26]) );
  OAI21X1 U285 ( .A(n955), .B(n858), .C(n891), .Y(n241) );
  XNOR2X1 U290 ( .A(n249), .B(n763), .Y(DIFF[25]) );
  AOI21X1 U291 ( .A(n252), .B(n838), .C(n246), .Y(n244) );
  OAI21X1 U293 ( .A(n890), .B(n968), .C(n810), .Y(n246) );
  XNOR2X1 U298 ( .A(n252), .B(n762), .Y(DIFF[24]) );
  OAI21X1 U299 ( .A(n957), .B(n829), .C(n890), .Y(n249) );
  XNOR2X1 U304 ( .A(n262), .B(n761), .Y(DIFF[23]) );
  AOI21X1 U306 ( .A(n296), .B(n840), .C(n255), .Y(n253) );
  OAI21X1 U308 ( .A(n853), .B(n827), .C(n743), .Y(n255) );
  AOI21X1 U310 ( .A(n267), .B(n722), .C(n259), .Y(n257) );
  OAI21X1 U312 ( .A(n889), .B(n878), .C(n809), .Y(n259) );
  XOR2X1 U317 ( .A(n857), .B(n779), .Y(DIFF[22]) );
  OAI21X1 U318 ( .A(n881), .B(n857), .C(n889), .Y(n262) );
  XNOR2X1 U323 ( .A(n270), .B(n760), .Y(DIFF[21]) );
  AOI21X1 U324 ( .A(n273), .B(n720), .C(n267), .Y(n265) );
  OAI21X1 U326 ( .A(n888), .B(n877), .C(n808), .Y(n267) );
  XNOR2X1 U331 ( .A(n273), .B(n759), .Y(DIFF[20]) );
  OAI21X1 U332 ( .A(n880), .B(n828), .C(n888), .Y(n270) );
  XNOR2X1 U337 ( .A(n283), .B(n758), .Y(DIFF[19]) );
  AOI21X1 U339 ( .A(n296), .B(n277), .C(n826), .Y(n274) );
  AOI21X1 U343 ( .A(n288), .B(n837), .C(n280), .Y(n278) );
  OAI21X1 U345 ( .A(n887), .B(n885), .C(n807), .Y(n280) );
  XOR2X1 U350 ( .A(n856), .B(n778), .Y(DIFF[18]) );
  OAI21X1 U351 ( .A(n876), .B(n856), .C(n887), .Y(n283) );
  XOR2X1 U356 ( .A(n750), .B(n777), .Y(DIFF[17]) );
  AOI21X1 U357 ( .A(n296), .B(n839), .C(n288), .Y(n286) );
  OAI21X1 U359 ( .A(n950), .B(n971), .C(n937), .Y(n288) );
  XNOR2X1 U364 ( .A(n296), .B(n757), .Y(DIFF[16]) );
  AOI21X1 U365 ( .A(n296), .B(n294), .C(n295), .Y(n291) );
  XOR2X1 U372 ( .A(n897), .B(n896), .Y(DIFF[15]) );
  AOI21X1 U374 ( .A(n347), .B(n727), .C(n299), .Y(n297) );
  OAI21X1 U376 ( .A(n721), .B(n845), .C(n742), .Y(n299) );
  AOI21X1 U378 ( .A(n315), .B(n919), .C(n303), .Y(n301) );
  OAI21X1 U380 ( .A(n946), .B(n970), .C(n802), .Y(n303) );
  XNOR2X1 U385 ( .A(n311), .B(n911), .Y(DIFF[14]) );
  AOI21X1 U386 ( .A(n311), .B(n309), .C(n310), .Y(n306) );
  XOR2X1 U393 ( .A(n749), .B(n776), .Y(DIFF[13]) );
  OAI21X1 U394 ( .A(n314), .B(n323), .C(n313), .Y(n311) );
  OAI21X1 U398 ( .A(n947), .B(n967), .C(n934), .Y(n315) );
  XOR2X1 U403 ( .A(n323), .B(n914), .Y(DIFF[12]) );
  AOI21X1 U404 ( .A(n324), .B(n321), .C(n322), .Y(n318) );
  XOR2X1 U411 ( .A(n926), .B(n925), .Y(DIFF[11]) );
  OAI21X1 U413 ( .A(n850), .B(n346), .C(n845), .Y(n324) );
  AOI21X1 U415 ( .A(n340), .B(n833), .C(n328), .Y(n326) );
  OAI21X1 U417 ( .A(n951), .B(n976), .C(n915), .Y(n328) );
  XNOR2X1 U422 ( .A(n336), .B(n756), .Y(DIFF[10]) );
  AOI21X1 U423 ( .A(n336), .B(n981), .C(n335), .Y(n331) );
  XNOR2X1 U430 ( .A(n343), .B(n894), .Y(DIFF[9]) );
  OAI21X1 U431 ( .A(n339), .B(n346), .C(n338), .Y(n336) );
  OAI21X1 U435 ( .A(n942), .B(n969), .C(n906), .Y(n340) );
  XOR2X1 U440 ( .A(n346), .B(n775), .Y(DIFF[8]) );
  OAI21X1 U441 ( .A(n920), .B(n346), .C(n942), .Y(n343) );
  XNOR2X1 U446 ( .A(n354), .B(n755), .Y(DIFF[7]) );
  OAI21X1 U448 ( .A(n748), .B(n907), .C(n741), .Y(n347) );
  AOI21X1 U450 ( .A(n359), .B(n939), .C(n351), .Y(n349) );
  OAI21X1 U452 ( .A(n886), .B(n965), .C(n806), .Y(n351) );
  XOR2X1 U457 ( .A(n855), .B(n774), .Y(DIFF[6]) );
  OAI21X1 U458 ( .A(n958), .B(n855), .C(n886), .Y(n354) );
  XOR2X1 U463 ( .A(n900), .B(n899), .Y(DIFF[5]) );
  AOI21X1 U464 ( .A(n367), .B(n918), .C(n359), .Y(n357) );
  OAI21X1 U466 ( .A(n948), .B(n966), .C(n935), .Y(n359) );
  XNOR2X1 U471 ( .A(n367), .B(n910), .Y(DIFF[4]) );
  AOI21X1 U472 ( .A(n367), .B(n365), .C(n366), .Y(n362) );
  XNOR2X1 U479 ( .A(n373), .B(n895), .Y(DIFF[3]) );
  AOI21X1 U481 ( .A(n377), .B(n908), .C(n370), .Y(n368) );
  OAI21X1 U483 ( .A(n959), .B(n940), .C(n916), .Y(n370) );
  XOR2X1 U488 ( .A(n376), .B(n923), .Y(DIFF[2]) );
  OAI21X1 U489 ( .A(n974), .B(n376), .C(n959), .Y(n373) );
  XOR2X1 U494 ( .A(n754), .B(n963), .Y(DIFF[1]) );
  OAI21X1 U496 ( .A(n963), .B(n917), .C(n898), .Y(n377) );
  XNOR2X1 U501 ( .A(n992), .B(A[0]), .Y(DIFF[0]) );
  INVX2 U570 ( .A(n872), .Y(n873) );
  AND2X2 U571 ( .A(n814), .B(n191), .Y(n26) );
  BUFX2 U572 ( .A(A[35]), .Y(n704) );
  BUFX2 U573 ( .A(n122), .Y(n705) );
  INVX1 U574 ( .A(B[31]), .Y(n1023) );
  AND2X1 U575 ( .A(n803), .B(n203), .Y(n28) );
  OR2X1 U576 ( .A(n878), .B(n881), .Y(n258) );
  OR2X1 U577 ( .A(n805), .B(n972), .Y(n164) );
  OR2X1 U578 ( .A(n714), .B(n928), .Y(n189) );
  OR2X1 U579 ( .A(n879), .B(n882), .Y(n216) );
  AND2X1 U580 ( .A(n1023), .B(A[31]), .Y(n219) );
  OR2X1 U581 ( .A(n804), .B(n853), .Y(n254) );
  AND2X1 U582 ( .A(n905), .B(n919), .Y(n300) );
  AND2X1 U583 ( .A(n802), .B(n304), .Y(n46) );
  AND2X1 U584 ( .A(n833), .B(n797), .Y(n325) );
  AND2X1 U585 ( .A(n843), .B(n730), .Y(n131) );
  AND2X1 U586 ( .A(n1034), .B(A[43]), .Y(n136) );
  AND2X1 U587 ( .A(n840), .B(n725), .Y(n210) );
  OR2X1 U588 ( .A(n956), .B(n975), .Y(n224) );
  AND2X1 U589 ( .A(n841), .B(n838), .Y(n235) );
  INVX1 U590 ( .A(B[28]), .Y(n1020) );
  AND2X1 U591 ( .A(n1017), .B(A[25]), .Y(n248) );
  OR2X1 U592 ( .A(n877), .B(n880), .Y(n266) );
  AND2X1 U593 ( .A(n1009), .B(A[17]), .Y(n290) );
  AND2X1 U594 ( .A(n1003), .B(A[11]), .Y(n330) );
  OR2X1 U595 ( .A(n997), .B(A[5]), .Y(n360) );
  AND2X1 U596 ( .A(A[3]), .B(n995), .Y(n372) );
  OR2X1 U597 ( .A(n993), .B(A[1]), .Y(n378) );
  AND2X1 U598 ( .A(A[1]), .B(n993), .Y(n379) );
  AND2X1 U599 ( .A(n945), .B(n985), .Y(n3) );
  AND2X1 U600 ( .A(n796), .B(n984), .Y(n5) );
  AND2X1 U601 ( .A(n795), .B(n990), .Y(n9) );
  OR2X1 U602 ( .A(n852), .B(n884), .Y(n126) );
  AND2X1 U603 ( .A(n1035), .B(A[44]), .Y(n129) );
  AND2X1 U604 ( .A(n987), .B(n711), .Y(n138) );
  AND2X1 U605 ( .A(n794), .B(n987), .Y(n19) );
  AND2X1 U606 ( .A(n1030), .B(A[39]), .Y(n167) );
  OR2X1 U607 ( .A(n1027), .B(A[36]), .Y(n183) );
  AND2X1 U608 ( .A(A[33]), .B(n1024), .Y(n204) );
  AND2X1 U609 ( .A(n1021), .B(A[29]), .Y(n227) );
  AND2X1 U610 ( .A(n1012), .B(A[20]), .Y(n272) );
  AND2X1 U611 ( .A(A[18]), .B(n1010), .Y(n285) );
  AND2X1 U612 ( .A(n915), .B(n329), .Y(n50) );
  AND2X1 U613 ( .A(A[5]), .B(n997), .Y(n361) );
  OR2X1 U614 ( .A(n996), .B(A[4]), .Y(n365) );
  AND2X1 U615 ( .A(A[2]), .B(n994), .Y(n375) );
  AND2X1 U616 ( .A(n944), .B(n989), .Y(n2) );
  AND2X1 U617 ( .A(A[38]), .B(n1029), .Y(n172) );
  BUFX2 U618 ( .A(n106), .Y(n706) );
  OR2X2 U619 ( .A(n1026), .B(A[35]), .Y(n191) );
  BUFX2 U620 ( .A(n847), .Y(n707) );
  BUFX2 U621 ( .A(n731), .Y(n708) );
  INVX1 U622 ( .A(n865), .Y(n709) );
  INVX1 U623 ( .A(n868), .Y(n710) );
  OR2X2 U624 ( .A(n851), .B(n717), .Y(n160) );
  AND2X2 U625 ( .A(n842), .B(n740), .Y(n162) );
  AND2X2 U626 ( .A(n149), .B(n154), .Y(n711) );
  INVX1 U627 ( .A(n711), .Y(n147) );
  AND2X1 U628 ( .A(n1045), .B(A[54]), .Y(n89) );
  OR2X1 U629 ( .A(A[44]), .B(n1035), .Y(n128) );
  AND2X1 U630 ( .A(n1047), .B(A[56]), .Y(n81) );
  OR2X1 U631 ( .A(A[31]), .B(n1023), .Y(n218) );
  OR2X1 U632 ( .A(A[25]), .B(n1017), .Y(n247) );
  OR2X1 U633 ( .A(A[17]), .B(n1009), .Y(n289) );
  OR2X1 U634 ( .A(n1010), .B(A[18]), .Y(n284) );
  OR2X1 U635 ( .A(n967), .B(n930), .Y(n314) );
  OR2X1 U636 ( .A(n927), .B(n978), .Y(n176) );
  OR2X1 U637 ( .A(n334), .B(n976), .Y(n327) );
  AND2X1 U638 ( .A(n1031), .B(A[40]), .Y(n155) );
  OR2X1 U639 ( .A(n994), .B(A[2]), .Y(n374) );
  OR2X1 U640 ( .A(n991), .B(A[32]), .Y(n206) );
  OR2X1 U641 ( .A(n1024), .B(A[33]), .Y(n203) );
  AND2X1 U642 ( .A(A[4]), .B(n996), .Y(n366) );
  OR2X1 U643 ( .A(n995), .B(A[3]), .Y(n371) );
  OAI21X1 U644 ( .A(n735), .B(n738), .C(n821), .Y(n712) );
  BUFX2 U645 ( .A(n90), .Y(n713) );
  INVX2 U646 ( .A(n191), .Y(n714) );
  AND2X1 U647 ( .A(A[36]), .B(n1027), .Y(n184) );
  AND2X2 U648 ( .A(A[32]), .B(n991), .Y(n207) );
  INVX1 U649 ( .A(n133), .Y(n715) );
  AND2X2 U650 ( .A(n834), .B(n724), .Y(n214) );
  OR2X2 U651 ( .A(A[56]), .B(n1047), .Y(n984) );
  OR2X1 U652 ( .A(A[43]), .B(n1034), .Y(n135) );
  OR2X1 U653 ( .A(A[29]), .B(n1021), .Y(n226) );
  BUFX2 U654 ( .A(n871), .Y(n716) );
  INVX1 U655 ( .A(n870), .Y(n871) );
  INVX1 U656 ( .A(n162), .Y(n717) );
  OAI21X1 U657 ( .A(n825), .B(n873), .C(n823), .Y(n718) );
  BUFX2 U658 ( .A(n875), .Y(n719) );
  INVX1 U659 ( .A(n874), .Y(n875) );
  AND2X2 U660 ( .A(n720), .B(n722), .Y(n256) );
  AND2X2 U661 ( .A(n1033), .B(A[42]), .Y(n143) );
  OR2X2 U662 ( .A(A[42]), .B(n1033), .Y(n987) );
  INVX2 U663 ( .A(B[20]), .Y(n1012) );
  OR2X1 U664 ( .A(A[10]), .B(n1002), .Y(n981) );
  OR2X2 U665 ( .A(A[54]), .B(n1045), .Y(n983) );
  INVX1 U666 ( .A(n266), .Y(n720) );
  INVX1 U667 ( .A(n300), .Y(n721) );
  INVX1 U668 ( .A(n258), .Y(n722) );
  INVX1 U669 ( .A(n235), .Y(n723) );
  INVX1 U670 ( .A(n216), .Y(n724) );
  OR2X2 U671 ( .A(n723), .B(n854), .Y(n212) );
  INVX1 U672 ( .A(n212), .Y(n725) );
  INVX1 U673 ( .A(n138), .Y(n726) );
  OR2X2 U674 ( .A(n850), .B(n721), .Y(n298) );
  INVX1 U675 ( .A(n298), .Y(n727) );
  INVX1 U676 ( .A(n126), .Y(n728) );
  INVX1 U677 ( .A(n210), .Y(n729) );
  INVX1 U678 ( .A(n160), .Y(n730) );
  BUFX2 U679 ( .A(n132), .Y(n731) );
  OR2X1 U680 ( .A(A[45]), .B(n1036), .Y(n123) );
  INVX1 U681 ( .A(n123), .Y(n732) );
  OR2X1 U682 ( .A(A[47]), .B(n1038), .Y(n115) );
  INVX1 U683 ( .A(n115), .Y(n733) );
  OR2X1 U684 ( .A(A[49]), .B(n1040), .Y(n107) );
  INVX1 U685 ( .A(n107), .Y(n734) );
  OR2X1 U686 ( .A(A[51]), .B(n1042), .Y(n99) );
  INVX1 U687 ( .A(n99), .Y(n735) );
  OR2X1 U688 ( .A(A[53]), .B(n1044), .Y(n91) );
  INVX1 U689 ( .A(n91), .Y(n736) );
  OR2X1 U690 ( .A(A[57]), .B(n1048), .Y(n75) );
  INVX1 U691 ( .A(n75), .Y(n737) );
  BUFX2 U692 ( .A(n101), .Y(n738) );
  BUFX2 U693 ( .A(n297), .Y(n739) );
  OR2X2 U694 ( .A(n955), .B(n977), .Y(n237) );
  INVX1 U695 ( .A(n176), .Y(n740) );
  BUFX2 U696 ( .A(n349), .Y(n741) );
  BUFX2 U697 ( .A(n301), .Y(n742) );
  BUFX2 U698 ( .A(n257), .Y(n743) );
  BUFX2 U699 ( .A(n215), .Y(n744) );
  INVX1 U700 ( .A(n211), .Y(n745) );
  INVX1 U701 ( .A(n745), .Y(n746) );
  BUFX2 U702 ( .A(n163), .Y(n747) );
  AND2X1 U703 ( .A(n939), .B(n918), .Y(n348) );
  INVX1 U704 ( .A(n348), .Y(n748) );
  BUFX2 U705 ( .A(n318), .Y(n749) );
  BUFX2 U706 ( .A(n291), .Y(n750) );
  BUFX2 U707 ( .A(n193), .Y(n751) );
  BUFX2 U708 ( .A(n180), .Y(n752) );
  BUFX2 U709 ( .A(n168), .Y(n753) );
  AND2X1 U710 ( .A(n898), .B(n378), .Y(n60) );
  INVX1 U711 ( .A(n60), .Y(n754) );
  AND2X1 U712 ( .A(n806), .B(n352), .Y(n54) );
  INVX1 U713 ( .A(n54), .Y(n755) );
  AND2X1 U714 ( .A(n951), .B(n981), .Y(n51) );
  INVX1 U715 ( .A(n51), .Y(n756) );
  AND2X1 U716 ( .A(n950), .B(n294), .Y(n45) );
  INVX1 U717 ( .A(n45), .Y(n757) );
  AND2X1 U718 ( .A(n807), .B(n281), .Y(n42) );
  INVX1 U719 ( .A(n42), .Y(n758) );
  AND2X1 U720 ( .A(n888), .B(n271), .Y(n41) );
  INVX1 U721 ( .A(n41), .Y(n759) );
  AND2X1 U722 ( .A(n808), .B(n268), .Y(n40) );
  INVX1 U723 ( .A(n40), .Y(n760) );
  AND2X1 U724 ( .A(n809), .B(n260), .Y(n38) );
  INVX1 U725 ( .A(n38), .Y(n761) );
  AND2X1 U726 ( .A(n890), .B(n250), .Y(n37) );
  INVX1 U727 ( .A(n37), .Y(n762) );
  AND2X1 U728 ( .A(n810), .B(n247), .Y(n36) );
  INVX1 U729 ( .A(n36), .Y(n763) );
  AND2X1 U730 ( .A(n811), .B(n239), .Y(n34) );
  INVX1 U731 ( .A(n34), .Y(n764) );
  AND2X1 U732 ( .A(n892), .B(n229), .Y(n33) );
  INVX1 U733 ( .A(n33), .Y(n765) );
  AND2X1 U734 ( .A(n812), .B(n226), .Y(n32) );
  INVX1 U735 ( .A(n32), .Y(n766) );
  AND2X1 U736 ( .A(n813), .B(n218), .Y(n30) );
  INVX1 U737 ( .A(n30), .Y(n767) );
  AND2X1 U738 ( .A(n816), .B(n399), .Y(n18) );
  INVX1 U739 ( .A(n18), .Y(n768) );
  AND2X1 U740 ( .A(n817), .B(n128), .Y(n17) );
  INVX1 U741 ( .A(n17), .Y(n769) );
  AND2X1 U742 ( .A(n798), .B(n982), .Y(n15) );
  INVX1 U743 ( .A(n15), .Y(n770) );
  AND2X1 U744 ( .A(n799), .B(n986), .Y(n13) );
  INVX1 U745 ( .A(n13), .Y(n771) );
  AND2X1 U746 ( .A(n800), .B(n988), .Y(n11) );
  INVX1 U747 ( .A(n11), .Y(n772) );
  AND2X1 U748 ( .A(n801), .B(n983), .Y(n7) );
  INVX1 U749 ( .A(n7), .Y(n773) );
  AND2X1 U750 ( .A(n886), .B(n355), .Y(n55) );
  INVX1 U751 ( .A(n55), .Y(n774) );
  AND2X1 U752 ( .A(n942), .B(n344), .Y(n53) );
  INVX1 U753 ( .A(n53), .Y(n775) );
  AND2X1 U754 ( .A(n934), .B(n316), .Y(n48) );
  INVX1 U755 ( .A(n48), .Y(n776) );
  AND2X1 U756 ( .A(n937), .B(n289), .Y(n44) );
  INVX1 U757 ( .A(n44), .Y(n777) );
  AND2X1 U758 ( .A(n887), .B(n284), .Y(n43) );
  INVX1 U759 ( .A(n43), .Y(n778) );
  AND2X1 U760 ( .A(n889), .B(n263), .Y(n39) );
  INVX1 U761 ( .A(n39), .Y(n779) );
  AND2X1 U762 ( .A(n891), .B(n242), .Y(n35) );
  INVX1 U763 ( .A(n35), .Y(n780) );
  AND2X1 U764 ( .A(n893), .B(n221), .Y(n31) );
  INVX1 U765 ( .A(n31), .Y(n781) );
  INVX1 U766 ( .A(n26), .Y(n782) );
  AND2X1 U767 ( .A(n936), .B(n178), .Y(n24) );
  INVX1 U768 ( .A(n24), .Y(n783) );
  AND2X1 U769 ( .A(n815), .B(n166), .Y(n22) );
  INVX1 U770 ( .A(n22), .Y(n784) );
  AND2X1 U771 ( .A(n818), .B(n123), .Y(n16) );
  INVX1 U772 ( .A(n16), .Y(n785) );
  AND2X1 U773 ( .A(n819), .B(n115), .Y(n14) );
  INVX1 U774 ( .A(n14), .Y(n786) );
  AND2X1 U775 ( .A(n820), .B(n107), .Y(n12) );
  INVX1 U776 ( .A(n12), .Y(n787) );
  AND2X1 U777 ( .A(n821), .B(n99), .Y(n10) );
  INVX1 U778 ( .A(n10), .Y(n788) );
  AND2X1 U779 ( .A(n822), .B(n91), .Y(n8) );
  INVX1 U780 ( .A(n8), .Y(n789) );
  AND2X1 U781 ( .A(n823), .B(n83), .Y(n6) );
  INVX1 U782 ( .A(n6), .Y(n790) );
  AND2X1 U783 ( .A(n824), .B(n75), .Y(n4) );
  INVX1 U784 ( .A(n4), .Y(n791) );
  INVX1 U785 ( .A(n793), .Y(n792) );
  OR2X1 U786 ( .A(n964), .B(n941), .Y(n201) );
  INVX1 U787 ( .A(n201), .Y(n793) );
  INVX1 U788 ( .A(n143), .Y(n794) );
  AND2X1 U789 ( .A(n1043), .B(A[52]), .Y(n97) );
  INVX1 U790 ( .A(n97), .Y(n795) );
  INVX1 U791 ( .A(n81), .Y(n796) );
  OR2X1 U792 ( .A(n969), .B(n920), .Y(n339) );
  INVX1 U793 ( .A(n339), .Y(n797) );
  AND2X1 U794 ( .A(n1037), .B(A[46]), .Y(n121) );
  INVX1 U795 ( .A(n121), .Y(n798) );
  AND2X1 U796 ( .A(A[48]), .B(n1039), .Y(n113) );
  INVX1 U797 ( .A(n113), .Y(n799) );
  AND2X1 U798 ( .A(A[50]), .B(n1041), .Y(n105) );
  INVX1 U799 ( .A(n105), .Y(n800) );
  INVX1 U800 ( .A(n89), .Y(n801) );
  AND2X1 U801 ( .A(n1007), .B(A[15]), .Y(n305) );
  INVX1 U802 ( .A(n305), .Y(n802) );
  INVX1 U803 ( .A(n204), .Y(n803) );
  AND2X1 U804 ( .A(n839), .B(n837), .Y(n277) );
  INVX1 U805 ( .A(n277), .Y(n804) );
  OR2X1 U806 ( .A(A[38]), .B(n1029), .Y(n171) );
  INVX1 U807 ( .A(n171), .Y(n805) );
  AND2X1 U808 ( .A(n999), .B(A[7]), .Y(n353) );
  INVX1 U809 ( .A(n353), .Y(n806) );
  AND2X1 U810 ( .A(n1011), .B(A[19]), .Y(n282) );
  INVX1 U811 ( .A(n282), .Y(n807) );
  AND2X1 U812 ( .A(n1013), .B(A[21]), .Y(n269) );
  INVX1 U813 ( .A(n269), .Y(n808) );
  AND2X1 U814 ( .A(n1015), .B(A[23]), .Y(n261) );
  INVX1 U815 ( .A(n261), .Y(n809) );
  INVX1 U816 ( .A(n248), .Y(n810) );
  AND2X1 U817 ( .A(n1019), .B(A[27]), .Y(n240) );
  INVX1 U818 ( .A(n240), .Y(n811) );
  INVX1 U819 ( .A(n227), .Y(n812) );
  INVX1 U820 ( .A(n219), .Y(n813) );
  AND2X1 U821 ( .A(n704), .B(n1026), .Y(n192) );
  INVX1 U822 ( .A(n192), .Y(n814) );
  INVX1 U823 ( .A(n167), .Y(n815) );
  INVX1 U824 ( .A(n136), .Y(n816) );
  INVX1 U825 ( .A(n129), .Y(n817) );
  AND2X1 U826 ( .A(n1036), .B(A[45]), .Y(n124) );
  INVX1 U827 ( .A(n124), .Y(n818) );
  AND2X1 U828 ( .A(n1038), .B(A[47]), .Y(n116) );
  INVX1 U829 ( .A(n116), .Y(n819) );
  AND2X1 U830 ( .A(n1040), .B(A[49]), .Y(n108) );
  INVX1 U831 ( .A(n108), .Y(n820) );
  AND2X1 U832 ( .A(n1042), .B(A[51]), .Y(n100) );
  INVX1 U833 ( .A(n100), .Y(n821) );
  AND2X1 U834 ( .A(n1044), .B(A[53]), .Y(n92) );
  INVX1 U835 ( .A(n92), .Y(n822) );
  AND2X1 U836 ( .A(n1046), .B(A[55]), .Y(n84) );
  INVX1 U837 ( .A(n84), .Y(n823) );
  AND2X1 U838 ( .A(n1048), .B(A[57]), .Y(n76) );
  INVX1 U839 ( .A(n76), .Y(n824) );
  INVX1 U840 ( .A(n83), .Y(n825) );
  OR2X1 U841 ( .A(A[55]), .B(n1046), .Y(n83) );
  INVX1 U842 ( .A(n827), .Y(n826) );
  BUFX2 U843 ( .A(n278), .Y(n827) );
  BUFX2 U844 ( .A(n274), .Y(n828) );
  BUFX2 U845 ( .A(n253), .Y(n829) );
  INVX1 U846 ( .A(n831), .Y(n830) );
  BUFX2 U847 ( .A(n236), .Y(n831) );
  BUFX2 U848 ( .A(n232), .Y(n832) );
  INVX1 U849 ( .A(n327), .Y(n833) );
  INVX1 U850 ( .A(n224), .Y(n834) );
  INVX1 U851 ( .A(n189), .Y(n835) );
  INVX1 U852 ( .A(n189), .Y(n836) );
  OR2X1 U853 ( .A(n876), .B(n885), .Y(n279) );
  INVX1 U854 ( .A(n279), .Y(n837) );
  OR2X1 U855 ( .A(n968), .B(n957), .Y(n245) );
  INVX1 U856 ( .A(n245), .Y(n838) );
  OR2X1 U857 ( .A(n971), .B(n932), .Y(n287) );
  INVX1 U858 ( .A(n287), .Y(n839) );
  INVX1 U859 ( .A(n254), .Y(n840) );
  INVX1 U860 ( .A(n237), .Y(n841) );
  INVX1 U861 ( .A(n164), .Y(n842) );
  OR2X2 U862 ( .A(n726), .B(n883), .Y(n133) );
  INVX1 U863 ( .A(n133), .Y(n843) );
  INVX1 U864 ( .A(n326), .Y(n844) );
  INVX1 U865 ( .A(n844), .Y(n845) );
  INVX1 U866 ( .A(n188), .Y(n846) );
  INVX1 U867 ( .A(n846), .Y(n847) );
  INVX1 U868 ( .A(n139), .Y(n848) );
  INVX1 U869 ( .A(n848), .Y(n849) );
  INVX1 U870 ( .A(n325), .Y(n850) );
  AND2X2 U871 ( .A(n793), .B(n836), .Y(n187) );
  INVX1 U872 ( .A(n187), .Y(n851) );
  INVX1 U873 ( .A(n131), .Y(n852) );
  INVX1 U874 ( .A(n256), .Y(n853) );
  INVX1 U875 ( .A(n214), .Y(n854) );
  BUFX2 U876 ( .A(n357), .Y(n855) );
  BUFX2 U877 ( .A(n286), .Y(n856) );
  BUFX2 U878 ( .A(n265), .Y(n857) );
  BUFX2 U879 ( .A(n244), .Y(n858) );
  BUFX2 U880 ( .A(n223), .Y(n859) );
  INVX1 U881 ( .A(n125), .Y(n860) );
  INVX1 U882 ( .A(n860), .Y(n861) );
  INVX1 U883 ( .A(n860), .Y(n862) );
  INVX1 U884 ( .A(n117), .Y(n863) );
  INVX1 U885 ( .A(n709), .Y(n864) );
  INVX1 U886 ( .A(n863), .Y(n865) );
  INVX1 U887 ( .A(n109), .Y(n866) );
  INVX1 U888 ( .A(n710), .Y(n867) );
  INVX1 U889 ( .A(n866), .Y(n868) );
  BUFX2 U890 ( .A(n738), .Y(n869) );
  INVX1 U891 ( .A(n93), .Y(n870) );
  INVX1 U892 ( .A(n85), .Y(n872) );
  INVX1 U893 ( .A(n77), .Y(n874) );
  INVX1 U894 ( .A(n284), .Y(n876) );
  INVX1 U895 ( .A(n268), .Y(n877) );
  OR2X1 U896 ( .A(A[21]), .B(n1013), .Y(n268) );
  INVX1 U897 ( .A(n260), .Y(n878) );
  OR2X1 U898 ( .A(A[23]), .B(n1015), .Y(n260) );
  INVX1 U899 ( .A(n218), .Y(n879) );
  OR2X1 U900 ( .A(A[20]), .B(n1012), .Y(n271) );
  INVX1 U901 ( .A(n271), .Y(n880) );
  OR2X1 U902 ( .A(A[22]), .B(n1014), .Y(n263) );
  INVX1 U903 ( .A(n263), .Y(n881) );
  OR2X1 U904 ( .A(A[30]), .B(n1022), .Y(n221) );
  INVX1 U905 ( .A(n221), .Y(n882) );
  INVX1 U906 ( .A(n135), .Y(n883) );
  INVX1 U907 ( .A(n128), .Y(n884) );
  OR2X1 U908 ( .A(A[19]), .B(n1011), .Y(n281) );
  INVX1 U909 ( .A(n281), .Y(n885) );
  AND2X1 U910 ( .A(n998), .B(A[6]), .Y(n356) );
  INVX1 U911 ( .A(n356), .Y(n886) );
  INVX1 U912 ( .A(n285), .Y(n887) );
  INVX1 U913 ( .A(n272), .Y(n888) );
  AND2X1 U914 ( .A(n1014), .B(A[22]), .Y(n264) );
  INVX1 U915 ( .A(n264), .Y(n889) );
  AND2X1 U916 ( .A(n1016), .B(A[24]), .Y(n251) );
  INVX1 U917 ( .A(n251), .Y(n890) );
  AND2X1 U918 ( .A(n1018), .B(A[26]), .Y(n243) );
  INVX1 U919 ( .A(n243), .Y(n891) );
  AND2X1 U920 ( .A(n1020), .B(A[28]), .Y(n230) );
  INVX1 U921 ( .A(n230), .Y(n892) );
  AND2X1 U922 ( .A(n1022), .B(A[30]), .Y(n222) );
  INVX1 U923 ( .A(n222), .Y(n893) );
  INVX1 U924 ( .A(B[10]), .Y(n1002) );
  AND2X1 U925 ( .A(n906), .B(n341), .Y(n52) );
  INVX1 U926 ( .A(n52), .Y(n894) );
  AND2X1 U927 ( .A(n916), .B(n371), .Y(n58) );
  INVX1 U928 ( .A(n58), .Y(n895) );
  INVX1 U929 ( .A(n46), .Y(n896) );
  BUFX2 U930 ( .A(n306), .Y(n897) );
  INVX1 U931 ( .A(n379), .Y(n898) );
  AND2X1 U932 ( .A(n935), .B(n360), .Y(n56) );
  INVX1 U933 ( .A(n56), .Y(n899) );
  BUFX2 U934 ( .A(n362), .Y(n900) );
  INVX1 U935 ( .A(n19), .Y(n901) );
  INVX1 U936 ( .A(n28), .Y(n902) );
  AND2X1 U937 ( .A(n938), .B(n149), .Y(n20) );
  INVX1 U938 ( .A(n20), .Y(n903) );
  BUFX2 U939 ( .A(n151), .Y(n904) );
  INVX1 U940 ( .A(n314), .Y(n905) );
  AND2X1 U941 ( .A(n1001), .B(A[9]), .Y(n342) );
  INVX1 U942 ( .A(n342), .Y(n906) );
  BUFX2 U943 ( .A(n368), .Y(n907) );
  OR2X1 U944 ( .A(n940), .B(n974), .Y(n369) );
  INVX1 U945 ( .A(n369), .Y(n908) );
  AND2X1 U946 ( .A(n952), .B(n196), .Y(n27) );
  INVX1 U947 ( .A(n27), .Y(n909) );
  AND2X1 U948 ( .A(n948), .B(n365), .Y(n57) );
  INVX1 U949 ( .A(n57), .Y(n910) );
  AND2X1 U950 ( .A(n946), .B(n309), .Y(n47) );
  INVX1 U951 ( .A(n47), .Y(n911) );
  AND2X1 U952 ( .A(n949), .B(n406), .Y(n25) );
  INVX1 U953 ( .A(n25), .Y(n912) );
  AND2X1 U954 ( .A(n954), .B(n402), .Y(n21) );
  INVX1 U955 ( .A(n21), .Y(n913) );
  AND2X1 U956 ( .A(n947), .B(n321), .Y(n49) );
  INVX1 U957 ( .A(n49), .Y(n914) );
  INVX1 U958 ( .A(n330), .Y(n915) );
  INVX1 U959 ( .A(n372), .Y(n916) );
  INVX1 U960 ( .A(n378), .Y(n917) );
  OR2X1 U961 ( .A(n966), .B(n929), .Y(n358) );
  INVX1 U962 ( .A(n358), .Y(n918) );
  OR2X1 U963 ( .A(n970), .B(n931), .Y(n302) );
  INVX1 U964 ( .A(n302), .Y(n919) );
  OR2X1 U965 ( .A(A[8]), .B(n1000), .Y(n344) );
  INVX1 U966 ( .A(n344), .Y(n920) );
  INVX1 U967 ( .A(n9), .Y(n921) );
  AND2X1 U968 ( .A(n953), .B(n404), .Y(n23) );
  INVX1 U969 ( .A(n23), .Y(n922) );
  AND2X1 U970 ( .A(n959), .B(n374), .Y(n59) );
  INVX1 U971 ( .A(n59), .Y(n923) );
  AND2X1 U972 ( .A(n960), .B(n206), .Y(n29) );
  INVX1 U973 ( .A(n29), .Y(n924) );
  INVX1 U974 ( .A(n50), .Y(n925) );
  BUFX2 U975 ( .A(n331), .Y(n926) );
  INVX1 U976 ( .A(n183), .Y(n927) );
  OR2X1 U977 ( .A(n1025), .B(A[34]), .Y(n196) );
  INVX1 U978 ( .A(n196), .Y(n928) );
  INVX1 U979 ( .A(n365), .Y(n929) );
  OR2X1 U980 ( .A(A[12]), .B(n1004), .Y(n321) );
  INVX1 U981 ( .A(n321), .Y(n930) );
  OR2X1 U982 ( .A(A[14]), .B(n1006), .Y(n309) );
  INVX1 U983 ( .A(n309), .Y(n931) );
  OR2X1 U984 ( .A(A[16]), .B(n1008), .Y(n294) );
  INVX1 U985 ( .A(n294), .Y(n932) );
  OR2X1 U986 ( .A(A[40]), .B(n1031), .Y(n154) );
  INVX1 U987 ( .A(n154), .Y(n933) );
  AND2X1 U988 ( .A(n1005), .B(A[13]), .Y(n317) );
  INVX1 U989 ( .A(n317), .Y(n934) );
  INVX1 U990 ( .A(n361), .Y(n935) );
  AND2X1 U991 ( .A(n1028), .B(A[37]), .Y(n179) );
  INVX1 U992 ( .A(n179), .Y(n936) );
  INVX1 U993 ( .A(n290), .Y(n937) );
  AND2X1 U994 ( .A(n1032), .B(A[41]), .Y(n150) );
  INVX1 U995 ( .A(n150), .Y(n938) );
  OR2X1 U996 ( .A(n965), .B(n958), .Y(n350) );
  INVX1 U997 ( .A(n350), .Y(n939) );
  INVX1 U998 ( .A(n371), .Y(n940) );
  INVX1 U999 ( .A(n203), .Y(n941) );
  AND2X1 U1000 ( .A(n1000), .B(A[8]), .Y(n345) );
  INVX1 U1001 ( .A(n345), .Y(n942) );
  INVX1 U1002 ( .A(n5), .Y(n943) );
  AND2X1 U1003 ( .A(n1051), .B(A[60]), .Y(n67) );
  INVX1 U1004 ( .A(n67), .Y(n944) );
  AND2X1 U1005 ( .A(n1049), .B(A[58]), .Y(n73) );
  INVX1 U1006 ( .A(n73), .Y(n945) );
  AND2X1 U1007 ( .A(n1006), .B(A[14]), .Y(n310) );
  INVX1 U1008 ( .A(n310), .Y(n946) );
  AND2X1 U1009 ( .A(n1004), .B(A[12]), .Y(n322) );
  INVX1 U1010 ( .A(n322), .Y(n947) );
  INVX1 U1011 ( .A(n366), .Y(n948) );
  INVX1 U1012 ( .A(n184), .Y(n949) );
  AND2X1 U1013 ( .A(n1008), .B(A[16]), .Y(n295) );
  INVX1 U1014 ( .A(n295), .Y(n950) );
  AND2X1 U1015 ( .A(n1002), .B(A[10]), .Y(n335) );
  INVX1 U1016 ( .A(n335), .Y(n951) );
  AND2X1 U1017 ( .A(A[34]), .B(n1025), .Y(n197) );
  INVX1 U1018 ( .A(n197), .Y(n952) );
  INVX1 U1019 ( .A(n172), .Y(n953) );
  INVX1 U1020 ( .A(n155), .Y(n954) );
  OR2X1 U1021 ( .A(A[26]), .B(n1018), .Y(n242) );
  INVX1 U1022 ( .A(n242), .Y(n955) );
  INVX1 U1023 ( .A(n226), .Y(n956) );
  OR2X1 U1024 ( .A(A[24]), .B(n1016), .Y(n250) );
  INVX1 U1025 ( .A(n250), .Y(n957) );
  OR2X1 U1026 ( .A(A[6]), .B(n998), .Y(n355) );
  INVX1 U1027 ( .A(n355), .Y(n958) );
  INVX1 U1028 ( .A(n375), .Y(n959) );
  INVX1 U1029 ( .A(n207), .Y(n960) );
  INVX1 U1030 ( .A(n2), .Y(n961) );
  INVX1 U1031 ( .A(n3), .Y(n962) );
  OR2X1 U1032 ( .A(n992), .B(A[0]), .Y(n380) );
  INVX1 U1033 ( .A(n380), .Y(n963) );
  INVX1 U1034 ( .A(n206), .Y(n964) );
  OR2X1 U1035 ( .A(A[7]), .B(n999), .Y(n352) );
  INVX1 U1036 ( .A(n352), .Y(n965) );
  INVX1 U1037 ( .A(n360), .Y(n966) );
  OR2X1 U1038 ( .A(A[13]), .B(n1005), .Y(n316) );
  INVX1 U1039 ( .A(n316), .Y(n967) );
  INVX1 U1040 ( .A(n247), .Y(n968) );
  OR2X1 U1041 ( .A(A[9]), .B(n1001), .Y(n341) );
  INVX1 U1042 ( .A(n341), .Y(n969) );
  OR2X1 U1043 ( .A(A[15]), .B(n1007), .Y(n304) );
  INVX1 U1044 ( .A(n304), .Y(n970) );
  INVX1 U1045 ( .A(n289), .Y(n971) );
  OR2X1 U1046 ( .A(A[39]), .B(n1030), .Y(n166) );
  INVX1 U1047 ( .A(n166), .Y(n972) );
  OR2X1 U1048 ( .A(A[41]), .B(n1032), .Y(n149) );
  INVX1 U1049 ( .A(n149), .Y(n973) );
  INVX1 U1050 ( .A(n374), .Y(n974) );
  OR2X1 U1051 ( .A(A[28]), .B(n1020), .Y(n229) );
  INVX1 U1052 ( .A(n229), .Y(n975) );
  OR2X1 U1053 ( .A(A[11]), .B(n1003), .Y(n329) );
  INVX1 U1054 ( .A(n329), .Y(n976) );
  OR2X1 U1055 ( .A(A[27]), .B(n1019), .Y(n239) );
  INVX1 U1056 ( .A(n239), .Y(n977) );
  OR2X1 U1057 ( .A(A[37]), .B(n1028), .Y(n178) );
  INVX1 U1058 ( .A(n178), .Y(n978) );
  BUFX2 U1059 ( .A(n114), .Y(n979) );
  BUFX2 U1060 ( .A(n74), .Y(n980) );
  INVX1 U1061 ( .A(n981), .Y(n334) );
  INVX1 U1062 ( .A(n209), .Y(n208) );
  INVX1 U1063 ( .A(n739), .Y(n296) );
  INVX1 U1064 ( .A(n157), .Y(n156) );
  INVX1 U1065 ( .A(n186), .Y(n185) );
  INVX1 U1066 ( .A(n324), .Y(n323) );
  INVX1 U1067 ( .A(n829), .Y(n252) );
  INVX1 U1068 ( .A(n828), .Y(n273) );
  INVX1 U1069 ( .A(n832), .Y(n231) );
  INVX1 U1070 ( .A(n177), .Y(n175) );
  INVX1 U1071 ( .A(n202), .Y(n200) );
  INVX1 U1072 ( .A(n315), .Y(n313) );
  INVX1 U1073 ( .A(n730), .Y(n158) );
  INVX1 U1074 ( .A(n161), .Y(n159) );
  INVX1 U1075 ( .A(n723), .Y(n233) );
  INVX1 U1076 ( .A(n347), .Y(n346) );
  INVX1 U1077 ( .A(n340), .Y(n338) );
  INVX1 U1078 ( .A(n377), .Y(n376) );
  INVX1 U1079 ( .A(n907), .Y(n367) );
  INVX1 U1080 ( .A(n148), .Y(n146) );
  INVX1 U1081 ( .A(n805), .Y(n404) );
  INVX1 U1082 ( .A(n933), .Y(n402) );
  OR2X1 U1083 ( .A(A[46]), .B(n1037), .Y(n982) );
  INVX1 U1084 ( .A(B[34]), .Y(n1025) );
  INVX1 U1085 ( .A(B[35]), .Y(n1026) );
  INVX1 U1086 ( .A(n883), .Y(n399) );
  INVX1 U1087 ( .A(n927), .Y(n406) );
  INVX1 U1088 ( .A(B[50]), .Y(n1041) );
  INVX1 U1089 ( .A(B[18]), .Y(n1010) );
  INVX1 U1090 ( .A(B[33]), .Y(n1024) );
  INVX1 U1091 ( .A(B[51]), .Y(n1042) );
  INVX1 U1092 ( .A(B[19]), .Y(n1011) );
  OR2X1 U1093 ( .A(A[58]), .B(n1049), .Y(n985) );
  INVX1 U1094 ( .A(B[58]), .Y(n1049) );
  INVX1 U1095 ( .A(B[26]), .Y(n1018) );
  INVX1 U1096 ( .A(B[42]), .Y(n1033) );
  INVX1 U1097 ( .A(B[36]), .Y(n1027) );
  INVX1 U1098 ( .A(B[57]), .Y(n1048) );
  INVX1 U1099 ( .A(B[24]), .Y(n1016) );
  INVX1 U1100 ( .A(B[40]), .Y(n1031) );
  INVX1 U1101 ( .A(B[25]), .Y(n1017) );
  INVX1 U1102 ( .A(B[41]), .Y(n1032) );
  INVX1 U1103 ( .A(B[56]), .Y(n1047) );
  INVX1 U1104 ( .A(B[49]), .Y(n1040) );
  INVX1 U1105 ( .A(B[16]), .Y(n1008) );
  INVX1 U1106 ( .A(B[48]), .Y(n1039) );
  INVX1 U1107 ( .A(B[9]), .Y(n1001) );
  OR2X1 U1108 ( .A(n1039), .B(A[48]), .Y(n986) );
  INVX1 U1109 ( .A(B[46]), .Y(n1037) );
  INVX1 U1110 ( .A(B[6]), .Y(n998) );
  INVX1 U1111 ( .A(B[38]), .Y(n1029) );
  INVX1 U1112 ( .A(B[2]), .Y(n994) );
  OR2X1 U1113 ( .A(n1041), .B(A[50]), .Y(n988) );
  INVX1 U1114 ( .A(B[3]), .Y(n995) );
  INVX1 U1115 ( .A(B[1]), .Y(n993) );
  INVX1 U1116 ( .A(B[4]), .Y(n996) );
  OR2X1 U1117 ( .A(A[60]), .B(n1051), .Y(n989) );
  INVX1 U1118 ( .A(B[61]), .Y(n1052) );
  INVX1 U1119 ( .A(n63), .Y(n381) );
  INVX1 U1120 ( .A(B[59]), .Y(n1050) );
  INVX1 U1121 ( .A(n69), .Y(n382) );
  XNOR2X1 U1122 ( .A(A[63]), .B(B[63]), .Y(n1) );
  INVX1 U1123 ( .A(B[32]), .Y(n991) );
  INVX1 U1124 ( .A(B[62]), .Y(n1053) );
  OR2X1 U1125 ( .A(A[52]), .B(n1043), .Y(n990) );
  INVX1 U1126 ( .A(B[30]), .Y(n1022) );
  INVX1 U1127 ( .A(B[29]), .Y(n1021) );
  INVX1 U1128 ( .A(B[27]), .Y(n1019) );
  INVX1 U1129 ( .A(B[12]), .Y(n1004) );
  INVX1 U1130 ( .A(B[13]), .Y(n1005) );
  INVX1 U1131 ( .A(B[14]), .Y(n1006) );
  INVX1 U1132 ( .A(B[11]), .Y(n1003) );
  INVX1 U1133 ( .A(B[44]), .Y(n1035) );
  INVX1 U1134 ( .A(B[45]), .Y(n1036) );
  INVX1 U1135 ( .A(B[43]), .Y(n1034) );
  INVX1 U1136 ( .A(B[7]), .Y(n999) );
  INVX1 U1137 ( .A(B[39]), .Y(n1030) );
  INVX1 U1138 ( .A(B[23]), .Y(n1015) );
  INVX1 U1139 ( .A(B[22]), .Y(n1014) );
  INVX1 U1140 ( .A(B[21]), .Y(n1013) );
  INVX1 U1141 ( .A(B[52]), .Y(n1043) );
  INVX1 U1142 ( .A(B[54]), .Y(n1045) );
  INVX1 U1143 ( .A(B[55]), .Y(n1046) );
  INVX1 U1144 ( .A(B[53]), .Y(n1044) );
  INVX1 U1145 ( .A(B[15]), .Y(n1007) );
  INVX1 U1146 ( .A(B[47]), .Y(n1038) );
  INVX1 U1147 ( .A(B[37]), .Y(n1028) );
  INVX1 U1148 ( .A(B[60]), .Y(n1051) );
  INVX1 U1149 ( .A(B[5]), .Y(n997) );
  INVX1 U1150 ( .A(B[0]), .Y(n992) );
  INVX1 U1151 ( .A(B[17]), .Y(n1009) );
  INVX1 U1152 ( .A(B[8]), .Y(n1000) );
endmodule


module alu_DW01_add_15 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n61, n62, n63, n64, n65, n69, n70, n71, n72, n73, n77, n78, n79,
         n80, n81, n85, n86, n87, n88, n89, n93, n94, n95, n96, n97, n101,
         n102, n103, n104, n105, n109, n110, n111, n112, n113, n117, n118,
         n119, n120, n121, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n139, n140, n142, n143, n144, n145,
         n146, n147, n150, n151, n152, n153, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n192, n193, n194, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n305, n306, n307,
         n309, n310, n311, n312, n313, n314, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n330, n331, n332, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n377, n378, n396, n397, n399, n400,
         n403, n408, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935;

  FAX1 U3 ( .A(B[62]), .B(A[62]), .C(n62), .YC(n61), .YS(SUM[62]) );
  FAX1 U4 ( .A(B[61]), .B(A[61]), .C(n63), .YC(n62), .YS(SUM[61]) );
  FAX1 U5 ( .A(B[60]), .B(A[60]), .C(n64), .YC(n63), .YS(SUM[60]) );
  FAX1 U6 ( .A(B[59]), .B(A[59]), .C(n378), .YC(n64), .YS(SUM[59]) );
  XNOR2X1 U8 ( .A(n658), .B(n894), .Y(SUM[58]) );
  AOI21X1 U9 ( .A(n70), .B(n930), .C(n69), .Y(n65) );
  XOR2X1 U16 ( .A(n839), .B(n741), .Y(SUM[57]) );
  OAI21X1 U17 ( .A(n671), .B(n673), .C(n783), .Y(n70) );
  XNOR2X1 U22 ( .A(n923), .B(n911), .Y(SUM[56]) );
  AOI21X1 U23 ( .A(n78), .B(n929), .C(n77), .Y(n73) );
  XOR2X1 U30 ( .A(n655), .B(n740), .Y(SUM[55]) );
  OAI21X1 U31 ( .A(n787), .B(n838), .C(n782), .Y(n78) );
  XNOR2X1 U36 ( .A(n924), .B(n719), .Y(SUM[54]) );
  AOI21X1 U37 ( .A(n86), .B(n934), .C(n85), .Y(n81) );
  XOR2X1 U44 ( .A(n652), .B(n739), .Y(SUM[53]) );
  OAI21X1 U45 ( .A(n786), .B(n836), .C(n781), .Y(n86) );
  XNOR2X1 U50 ( .A(n921), .B(n910), .Y(SUM[52]) );
  AOI21X1 U51 ( .A(n94), .B(n933), .C(n93), .Y(n89) );
  XOR2X1 U58 ( .A(n833), .B(n738), .Y(SUM[51]) );
  OAI21X1 U59 ( .A(n670), .B(n834), .C(n780), .Y(n94) );
  XNOR2X1 U64 ( .A(n659), .B(n718), .Y(SUM[50]) );
  AOI21X1 U65 ( .A(n102), .B(n931), .C(n101), .Y(n97) );
  XOR2X1 U72 ( .A(n657), .B(n737), .Y(SUM[49]) );
  OAI21X1 U73 ( .A(n669), .B(n672), .C(n779), .Y(n102) );
  XNOR2X1 U78 ( .A(n935), .B(n717), .Y(SUM[48]) );
  AOI21X1 U79 ( .A(n110), .B(n926), .C(n109), .Y(n105) );
  XOR2X1 U86 ( .A(n830), .B(n736), .Y(SUM[47]) );
  OAI21X1 U87 ( .A(n785), .B(n831), .C(n778), .Y(n110) );
  XNOR2X1 U92 ( .A(n922), .B(n908), .Y(SUM[46]) );
  AOI21X1 U93 ( .A(n118), .B(n928), .C(n117), .Y(n113) );
  XOR2X1 U100 ( .A(n827), .B(n735), .Y(SUM[45]) );
  OAI21X1 U101 ( .A(n784), .B(n828), .C(n777), .Y(n118) );
  XNOR2X1 U106 ( .A(n126), .B(n716), .Y(SUM[44]) );
  AOI21X1 U107 ( .A(n205), .B(n662), .C(n123), .Y(n121) );
  OAI21X1 U109 ( .A(n914), .B(n814), .C(n776), .Y(n123) );
  XNOR2X1 U114 ( .A(n133), .B(n715), .Y(SUM[43]) );
  OAI21X1 U115 ( .A(n818), .B(n204), .C(n661), .Y(n126) );
  AOI21X1 U117 ( .A(n641), .B(n799), .C(n130), .Y(n128) );
  OAI21X1 U119 ( .A(n916), .B(n812), .C(n775), .Y(n130) );
  XNOR2X1 U124 ( .A(n140), .B(n909), .Y(SUM[42]) );
  OAI21X1 U125 ( .A(n817), .B(n152), .C(n645), .Y(n133) );
  AOI21X1 U127 ( .A(n639), .B(n927), .C(n139), .Y(n135) );
  XOR2X1 U134 ( .A(n696), .B(n734), .Y(SUM[41]) );
  OAI21X1 U135 ( .A(n143), .B(n152), .C(n142), .Y(n140) );
  OAI21X1 U139 ( .A(n846), .B(n860), .C(n774), .Y(n144) );
  XOR2X1 U144 ( .A(n152), .B(n733), .Y(SUM[40]) );
  AOI21X1 U145 ( .A(n153), .B(n397), .C(n151), .Y(n147) );
  XOR2X1 U152 ( .A(n695), .B(n732), .Y(SUM[39]) );
  OAI21X1 U154 ( .A(n156), .B(n204), .C(n155), .Y(n153) );
  OAI21X1 U158 ( .A(n820), .B(n668), .C(n684), .Y(n157) );
  AOI21X1 U160 ( .A(n173), .B(n677), .C(n161), .Y(n159) );
  OAI21X1 U162 ( .A(n845), .B(n859), .C(n773), .Y(n161) );
  XNOR2X1 U167 ( .A(n169), .B(n714), .Y(SUM[38]) );
  AOI21X1 U168 ( .A(n169), .B(n399), .C(n168), .Y(n164) );
  XOR2X1 U175 ( .A(n694), .B(n731), .Y(SUM[37]) );
  OAI21X1 U176 ( .A(n170), .B(n181), .C(n171), .Y(n169) );
  OAI21X1 U180 ( .A(n844), .B(n869), .C(n772), .Y(n173) );
  XOR2X1 U185 ( .A(n181), .B(n730), .Y(SUM[36]) );
  AOI21X1 U186 ( .A(n182), .B(n179), .C(n180), .Y(n176) );
  XOR2X1 U193 ( .A(n883), .B(n882), .Y(SUM[35]) );
  OAI21X1 U195 ( .A(n667), .B(n204), .C(n811), .Y(n182) );
  AOI21X1 U197 ( .A(n660), .B(n198), .C(n186), .Y(n184) );
  OAI21X1 U199 ( .A(n903), .B(n644), .C(n753), .Y(n186) );
  XNOR2X1 U204 ( .A(n194), .B(n889), .Y(SUM[34]) );
  AOI21X1 U205 ( .A(n194), .B(n403), .C(n193), .Y(n189) );
  XNOR2X1 U212 ( .A(n201), .B(n713), .Y(SUM[33]) );
  OAI21X1 U213 ( .A(n197), .B(n204), .C(n196), .Y(n194) );
  OAI21X1 U217 ( .A(n848), .B(n868), .C(n771), .Y(n198) );
  XOR2X1 U222 ( .A(n204), .B(n897), .Y(SUM[32]) );
  OAI21X1 U223 ( .A(n912), .B(n204), .C(n847), .Y(n201) );
  XNOR2X1 U228 ( .A(n216), .B(n712), .Y(SUM[31]) );
  OAI21X1 U230 ( .A(n665), .B(n675), .C(n683), .Y(n205) );
  AOI21X1 U232 ( .A(n251), .B(n806), .C(n209), .Y(n207) );
  OAI21X1 U234 ( .A(n816), .B(n795), .C(n681), .Y(n209) );
  AOI21X1 U236 ( .A(n221), .B(n801), .C(n213), .Y(n211) );
  OAI21X1 U238 ( .A(n877), .B(n858), .C(n770), .Y(n213) );
  XOR2X1 U243 ( .A(n825), .B(n729), .Y(SUM[30]) );
  OAI21X1 U244 ( .A(n867), .B(n825), .C(n877), .Y(n216) );
  XNOR2X1 U249 ( .A(n224), .B(n711), .Y(SUM[29]) );
  AOI21X1 U250 ( .A(n227), .B(n798), .C(n221), .Y(n219) );
  OAI21X1 U252 ( .A(n876), .B(n857), .C(n769), .Y(n221) );
  XNOR2X1 U257 ( .A(n227), .B(n710), .Y(SUM[28]) );
  OAI21X1 U258 ( .A(n866), .B(n796), .C(n876), .Y(n224) );
  XNOR2X1 U263 ( .A(n237), .B(n709), .Y(SUM[27]) );
  AOI21X1 U265 ( .A(n248), .B(n231), .C(n794), .Y(n228) );
  AOI21X1 U269 ( .A(n242), .B(n805), .C(n234), .Y(n232) );
  OAI21X1 U271 ( .A(n875), .B(n856), .C(n768), .Y(n234) );
  XOR2X1 U276 ( .A(n824), .B(n728), .Y(SUM[26]) );
  OAI21X1 U277 ( .A(n865), .B(n824), .C(n875), .Y(n237) );
  XNOR2X1 U282 ( .A(n245), .B(n708), .Y(SUM[25]) );
  AOI21X1 U283 ( .A(n248), .B(n745), .C(n242), .Y(n240) );
  OAI21X1 U285 ( .A(n874), .B(n855), .C(n767), .Y(n242) );
  XNOR2X1 U290 ( .A(n248), .B(n707), .Y(SUM[24]) );
  OAI21X1 U291 ( .A(n864), .B(n793), .C(n874), .Y(n245) );
  XNOR2X1 U296 ( .A(n258), .B(n706), .Y(SUM[23]) );
  AOI21X1 U298 ( .A(n292), .B(n810), .C(n251), .Y(n249) );
  OAI21X1 U300 ( .A(n815), .B(n791), .C(n680), .Y(n251) );
  AOI21X1 U302 ( .A(n263), .B(n800), .C(n255), .Y(n253) );
  OAI21X1 U304 ( .A(n873), .B(n854), .C(n766), .Y(n255) );
  XOR2X1 U309 ( .A(n823), .B(n727), .Y(SUM[22]) );
  OAI21X1 U310 ( .A(n863), .B(n823), .C(n873), .Y(n258) );
  XNOR2X1 U315 ( .A(n266), .B(n705), .Y(SUM[21]) );
  AOI21X1 U316 ( .A(n269), .B(n797), .C(n263), .Y(n261) );
  OAI21X1 U318 ( .A(n872), .B(n853), .C(n765), .Y(n263) );
  XNOR2X1 U323 ( .A(n269), .B(n704), .Y(SUM[20]) );
  OAI21X1 U324 ( .A(n862), .B(n792), .C(n872), .Y(n266) );
  XNOR2X1 U329 ( .A(n279), .B(n703), .Y(SUM[19]) );
  AOI21X1 U331 ( .A(n292), .B(n273), .C(n790), .Y(n270) );
  AOI21X1 U335 ( .A(n284), .B(n804), .C(n276), .Y(n274) );
  OAI21X1 U337 ( .A(n871), .B(n906), .C(n764), .Y(n276) );
  XOR2X1 U342 ( .A(n822), .B(n726), .Y(SUM[18]) );
  OAI21X1 U343 ( .A(n915), .B(n822), .C(n871), .Y(n279) );
  XOR2X1 U348 ( .A(n693), .B(n725), .Y(SUM[17]) );
  AOI21X1 U349 ( .A(n292), .B(n809), .C(n284), .Y(n282) );
  OAI21X1 U351 ( .A(n892), .B(n905), .C(n887), .Y(n284) );
  XNOR2X1 U356 ( .A(n292), .B(n702), .Y(SUM[16]) );
  AOI21X1 U357 ( .A(n292), .B(n290), .C(n291), .Y(n287) );
  XOR2X1 U364 ( .A(n692), .B(n724), .Y(SUM[15]) );
  AOI21X1 U366 ( .A(n343), .B(n687), .C(n295), .Y(n293) );
  OAI21X1 U368 ( .A(n663), .B(n788), .C(n679), .Y(n295) );
  AOI21X1 U370 ( .A(n311), .B(n803), .C(n299), .Y(n297) );
  OAI21X1 U372 ( .A(n843), .B(n852), .C(n763), .Y(n299) );
  XNOR2X1 U377 ( .A(n307), .B(n701), .Y(SUM[14]) );
  AOI21X1 U378 ( .A(n307), .B(n305), .C(n306), .Y(n302) );
  XOR2X1 U385 ( .A(n691), .B(n723), .Y(SUM[13]) );
  OAI21X1 U386 ( .A(n310), .B(n319), .C(n309), .Y(n307) );
  OAI21X1 U390 ( .A(n842), .B(n851), .C(n762), .Y(n311) );
  XOR2X1 U395 ( .A(n319), .B(n722), .Y(SUM[12]) );
  AOI21X1 U396 ( .A(n320), .B(n317), .C(n318), .Y(n314) );
  XOR2X1 U403 ( .A(n690), .B(n896), .Y(SUM[11]) );
  OAI21X1 U405 ( .A(n819), .B(n342), .C(n788), .Y(n320) );
  AOI21X1 U407 ( .A(n336), .B(n686), .C(n324), .Y(n322) );
  OAI21X1 U409 ( .A(n841), .B(n920), .C(n752), .Y(n324) );
  XNOR2X1 U414 ( .A(n332), .B(n700), .Y(SUM[10]) );
  AOI21X1 U415 ( .A(n332), .B(n330), .C(n331), .Y(n327) );
  XNOR2X1 U422 ( .A(n339), .B(n881), .Y(SUM[9]) );
  OAI21X1 U423 ( .A(n335), .B(n342), .C(n334), .Y(n332) );
  OAI21X1 U427 ( .A(n907), .B(n893), .C(n888), .Y(n336) );
  XOR2X1 U432 ( .A(n342), .B(n890), .Y(SUM[8]) );
  OAI21X1 U433 ( .A(n913), .B(n342), .C(n907), .Y(n339) );
  XNOR2X1 U438 ( .A(n350), .B(n699), .Y(SUM[7]) );
  OAI21X1 U440 ( .A(n688), .B(n789), .C(n678), .Y(n343) );
  AOI21X1 U442 ( .A(n355), .B(n808), .C(n347), .Y(n345) );
  OAI21X1 U444 ( .A(n870), .B(n850), .C(n761), .Y(n347) );
  XOR2X1 U449 ( .A(n821), .B(n721), .Y(SUM[6]) );
  OAI21X1 U450 ( .A(n861), .B(n821), .C(n870), .Y(n350) );
  XOR2X1 U455 ( .A(n689), .B(n720), .Y(SUM[5]) );
  AOI21X1 U456 ( .A(n363), .B(n802), .C(n355), .Y(n353) );
  OAI21X1 U458 ( .A(n840), .B(n849), .C(n760), .Y(n355) );
  XNOR2X1 U463 ( .A(n363), .B(n698), .Y(SUM[4]) );
  AOI21X1 U464 ( .A(n363), .B(n361), .C(n362), .Y(n358) );
  XNOR2X1 U471 ( .A(n369), .B(n879), .Y(SUM[3]) );
  AOI21X1 U473 ( .A(n373), .B(n685), .C(n366), .Y(n364) );
  OAI21X1 U475 ( .A(n918), .B(n904), .C(n886), .Y(n366) );
  XOR2X1 U480 ( .A(n372), .B(n895), .Y(SUM[2]) );
  OAI21X1 U481 ( .A(n925), .B(n372), .C(n918), .Y(n369) );
  XOR2X1 U486 ( .A(n697), .B(n919), .Y(SUM[1]) );
  OAI21X1 U488 ( .A(n919), .B(n880), .C(n878), .Y(n373) );
  BUFX2 U501 ( .A(B[43]), .Y(n636) );
  AND2X2 U502 ( .A(n775), .B(n131), .Y(n17) );
  INVX2 U503 ( .A(n158), .Y(n820) );
  BUFX2 U504 ( .A(B[31]), .Y(n637) );
  OR2X2 U505 ( .A(n759), .B(n860), .Y(n143) );
  INVX1 U506 ( .A(n145), .Y(n860) );
  OR2X2 U507 ( .A(B[31]), .B(A[31]), .Y(n214) );
  AND2X2 U508 ( .A(n637), .B(A[31]), .Y(n215) );
  AND2X2 U509 ( .A(B[30]), .B(A[30]), .Y(n218) );
  OR2X2 U510 ( .A(B[30]), .B(A[30]), .Y(n217) );
  BUFX2 U511 ( .A(n205), .Y(n638) );
  OR2X1 U512 ( .A(A[16]), .B(B[16]), .Y(n290) );
  OR2X2 U513 ( .A(A[41]), .B(B[41]), .Y(n145) );
  AND2X2 U514 ( .A(B[57]), .B(A[57]), .Y(n72) );
  OR2X2 U515 ( .A(A[57]), .B(B[57]), .Y(n71) );
  AND2X2 U516 ( .A(B[16]), .B(A[16]), .Y(n291) );
  AND2X1 U517 ( .A(n808), .B(n802), .Y(n344) );
  OR2X1 U518 ( .A(A[56]), .B(B[56]), .Y(n929) );
  INVX1 U519 ( .A(n146), .Y(n774) );
  OR2X1 U520 ( .A(B[5]), .B(A[5]), .Y(n356) );
  AND2X1 U521 ( .A(B[45]), .B(A[45]), .Y(n120) );
  AND2X1 U522 ( .A(B[55]), .B(A[55]), .Y(n80) );
  OR2X1 U523 ( .A(A[39]), .B(B[39]), .Y(n162) );
  AND2X1 U524 ( .A(B[39]), .B(A[39]), .Y(n163) );
  OR2X1 U525 ( .A(n858), .B(n867), .Y(n212) );
  OR2X1 U526 ( .A(n856), .B(n865), .Y(n233) );
  OR2X1 U527 ( .A(n815), .B(n676), .Y(n250) );
  AND2X1 U528 ( .A(n746), .B(n803), .Y(n296) );
  AND2X1 U529 ( .A(B[15]), .B(A[15]), .Y(n301) );
  AND2X1 U530 ( .A(n884), .B(n686), .Y(n321) );
  AND2X1 U531 ( .A(B[9]), .B(A[9]), .Y(n338) );
  AND2X1 U532 ( .A(B[53]), .B(A[53]), .Y(n88) );
  AND2X1 U533 ( .A(B[51]), .B(A[51]), .Y(n96) );
  OR2X1 U534 ( .A(A[50]), .B(B[50]), .Y(n931) );
  OR2X1 U535 ( .A(A[48]), .B(B[48]), .Y(n926) );
  AND2X1 U536 ( .A(n636), .B(A[43]), .Y(n132) );
  AND2X1 U537 ( .A(n747), .B(n807), .Y(n183) );
  AND2X1 U538 ( .A(B[27]), .B(A[27]), .Y(n236) );
  OR2X1 U539 ( .A(n855), .B(n864), .Y(n241) );
  AND2X1 U540 ( .A(B[25]), .B(A[25]), .Y(n244) );
  OR2X1 U541 ( .A(n853), .B(n862), .Y(n262) );
  AND2X1 U542 ( .A(B[21]), .B(A[21]), .Y(n265) );
  AND2X1 U543 ( .A(B[20]), .B(A[20]), .Y(n268) );
  OR2X1 U544 ( .A(n756), .B(n905), .Y(n283) );
  AND2X1 U545 ( .A(B[17]), .B(A[17]), .Y(n286) );
  OR2X1 U546 ( .A(B[1]), .B(A[1]), .Y(n374) );
  AND2X1 U547 ( .A(A[1]), .B(B[1]), .Y(n375) );
  AND2X1 U548 ( .A(n743), .B(n930), .Y(n2) );
  AND2X1 U549 ( .A(n899), .B(n929), .Y(n4) );
  AND2X1 U550 ( .A(n901), .B(n933), .Y(n8) );
  AND2X1 U551 ( .A(B[49]), .B(A[49]), .Y(n104) );
  AND2X1 U552 ( .A(n927), .B(n744), .Y(n134) );
  AND2X1 U553 ( .A(n900), .B(n927), .Y(n18) );
  AND2X1 U554 ( .A(n846), .B(n397), .Y(n20) );
  AND2X1 U555 ( .A(B[37]), .B(A[37]), .Y(n175) );
  AND2X1 U556 ( .A(n753), .B(n650), .Y(n25) );
  AND2X1 U557 ( .A(A[32]), .B(B[32]), .Y(n203) );
  OR2X1 U558 ( .A(B[32]), .B(A[32]), .Y(n202) );
  AND2X1 U559 ( .A(B[18]), .B(A[18]), .Y(n281) );
  AND2X1 U560 ( .A(n752), .B(n325), .Y(n49) );
  AND2X1 U561 ( .A(A[5]), .B(B[5]), .Y(n357) );
  AND2X1 U562 ( .A(A[2]), .B(B[2]), .Y(n371) );
  AND2X1 U563 ( .A(B[38]), .B(A[38]), .Y(n168) );
  OR2X1 U564 ( .A(A[38]), .B(B[38]), .Y(n651) );
  OR2X1 U565 ( .A(B[34]), .B(A[34]), .Y(n192) );
  AND2X1 U566 ( .A(n847), .B(n202), .Y(n28) );
  OR2X1 U567 ( .A(n849), .B(n754), .Y(n354) );
  INVX1 U568 ( .A(n377), .Y(n919) );
  OR2X1 U569 ( .A(A[6]), .B(B[6]), .Y(n351) );
  AND2X1 U570 ( .A(B[6]), .B(A[6]), .Y(n352) );
  AND2X1 U571 ( .A(n898), .B(n928), .Y(n14) );
  OAI21X1 U572 ( .A(n846), .B(n860), .C(n774), .Y(n639) );
  BUFX2 U573 ( .A(n144), .Y(n640) );
  OAI21X1 U574 ( .A(n820), .B(n668), .C(n684), .Y(n641) );
  BUFX2 U575 ( .A(n157), .Y(n642) );
  OR2X2 U576 ( .A(A[35]), .B(B[35]), .Y(n643) );
  AND2X2 U577 ( .A(A[36]), .B(B[36]), .Y(n180) );
  OR2X2 U578 ( .A(B[36]), .B(A[36]), .Y(n179) );
  INVX2 U579 ( .A(n187), .Y(n644) );
  BUFX2 U580 ( .A(n812), .Y(n645) );
  BUFX2 U581 ( .A(n834), .Y(n646) );
  INVX1 U582 ( .A(A[41]), .Y(n647) );
  INVX1 U583 ( .A(n647), .Y(n648) );
  BUFX2 U584 ( .A(n831), .Y(n649) );
  INVX1 U585 ( .A(n917), .Y(n650) );
  AND2X2 U586 ( .A(B[42]), .B(A[42]), .Y(n139) );
  OR2X1 U587 ( .A(n851), .B(n757), .Y(n310) );
  AND2X1 U588 ( .A(B[58]), .B(A[58]), .Y(n69) );
  OR2X1 U589 ( .A(A[55]), .B(B[55]), .Y(n79) );
  OR2X1 U590 ( .A(A[45]), .B(B[45]), .Y(n119) );
  AND2X1 U591 ( .A(B[48]), .B(A[48]), .Y(n109) );
  OR2X1 U592 ( .A(A[53]), .B(B[53]), .Y(n87) );
  OR2X1 U593 ( .A(A[25]), .B(B[25]), .Y(n243) );
  AND2X1 U594 ( .A(B[52]), .B(A[52]), .Y(n93) );
  AND2X1 U595 ( .A(B[56]), .B(A[56]), .Y(n77) );
  OR2X1 U596 ( .A(A[20]), .B(B[20]), .Y(n267) );
  OR2X1 U597 ( .A(A[27]), .B(B[27]), .Y(n235) );
  OR2X1 U598 ( .A(A[44]), .B(B[44]), .Y(n124) );
  OR2X1 U599 ( .A(A[51]), .B(B[51]), .Y(n95) );
  OR2X1 U600 ( .A(A[23]), .B(B[23]), .Y(n256) );
  OR2X1 U601 ( .A(A[18]), .B(B[18]), .Y(n280) );
  OR2X1 U602 ( .A(A[49]), .B(B[49]), .Y(n103) );
  INVX1 U603 ( .A(n151), .Y(n846) );
  AND2X1 U604 ( .A(B[40]), .B(A[40]), .Y(n151) );
  OR2X1 U605 ( .A(A[40]), .B(B[40]), .Y(n150) );
  AND2X1 U606 ( .A(B[14]), .B(A[14]), .Y(n306) );
  OR2X1 U607 ( .A(A[21]), .B(B[21]), .Y(n264) );
  OR2X1 U608 ( .A(A[28]), .B(B[28]), .Y(n225) );
  OR2X1 U609 ( .A(A[17]), .B(B[17]), .Y(n285) );
  INVX1 U610 ( .A(n277), .Y(n906) );
  OR2X1 U611 ( .A(A[19]), .B(B[19]), .Y(n277) );
  OR2X1 U612 ( .A(B[2]), .B(A[2]), .Y(n370) );
  OR2X1 U613 ( .A(A[9]), .B(B[9]), .Y(n337) );
  AND2X1 U614 ( .A(B[29]), .B(A[29]), .Y(n223) );
  OR2X1 U615 ( .A(n751), .B(n869), .Y(n172) );
  OR2X2 U616 ( .A(n758), .B(n859), .Y(n160) );
  OR2X1 U617 ( .A(A[37]), .B(B[37]), .Y(n174) );
  BUFX2 U618 ( .A(n836), .Y(n652) );
  XNOR2X1 U619 ( .A(n61), .B(n653), .Y(SUM[63]) );
  XNOR2X1 U620 ( .A(A[63]), .B(B[63]), .Y(n653) );
  INVX1 U621 ( .A(n649), .Y(n654) );
  BUFX2 U622 ( .A(n838), .Y(n655) );
  INVX1 U623 ( .A(n646), .Y(n656) );
  BUFX2 U624 ( .A(n672), .Y(n657) );
  AND2X2 U625 ( .A(B[44]), .B(A[44]), .Y(n125) );
  OAI21X1 U626 ( .A(n671), .B(n839), .C(n783), .Y(n658) );
  OAI21X1 U627 ( .A(n669), .B(n657), .C(n779), .Y(n659) );
  INVX1 U628 ( .A(n185), .Y(n660) );
  AND2X1 U629 ( .A(n127), .B(n124), .Y(n662) );
  OR2X2 U630 ( .A(A[35]), .B(B[35]), .Y(n187) );
  INVX2 U631 ( .A(n643), .Y(n917) );
  OR2X2 U632 ( .A(n917), .B(n885), .Y(n185) );
  BUFX2 U633 ( .A(n814), .Y(n661) );
  AND2X2 U634 ( .A(n797), .B(n800), .Y(n252) );
  OR2X2 U635 ( .A(n857), .B(n866), .Y(n220) );
  AND2X2 U636 ( .A(n809), .B(n804), .Y(n273) );
  OR2X1 U637 ( .A(A[10]), .B(B[10]), .Y(n330) );
  OR2X2 U638 ( .A(A[42]), .B(B[42]), .Y(n927) );
  INVX1 U639 ( .A(n296), .Y(n663) );
  AND2X2 U640 ( .A(n745), .B(n805), .Y(n231) );
  INVX1 U641 ( .A(n231), .Y(n664) );
  AND2X2 U642 ( .A(n810), .B(n806), .Y(n206) );
  INVX1 U643 ( .A(n206), .Y(n665) );
  OR2X2 U644 ( .A(n667), .B(n820), .Y(n156) );
  INVX1 U645 ( .A(n156), .Y(n666) );
  INVX1 U646 ( .A(n183), .Y(n667) );
  BUFX2 U647 ( .A(n184), .Y(n668) );
  INVX1 U648 ( .A(n103), .Y(n669) );
  INVX1 U649 ( .A(n95), .Y(n670) );
  INVX1 U650 ( .A(n71), .Y(n671) );
  BUFX2 U651 ( .A(n105), .Y(n672) );
  BUFX2 U652 ( .A(n73), .Y(n673) );
  OR2X2 U653 ( .A(n817), .B(n916), .Y(n129) );
  AND2X2 U654 ( .A(n648), .B(B[41]), .Y(n146) );
  INVX1 U655 ( .A(n293), .Y(n674) );
  INVX1 U656 ( .A(n674), .Y(n675) );
  INVX1 U657 ( .A(n273), .Y(n676) );
  INVX1 U658 ( .A(n160), .Y(n677) );
  BUFX2 U659 ( .A(n345), .Y(n678) );
  BUFX2 U660 ( .A(n297), .Y(n679) );
  BUFX2 U661 ( .A(n253), .Y(n680) );
  BUFX2 U662 ( .A(n211), .Y(n681) );
  INVX1 U663 ( .A(n207), .Y(n682) );
  INVX1 U664 ( .A(n682), .Y(n683) );
  BUFX2 U665 ( .A(n159), .Y(n684) );
  OR2X1 U666 ( .A(n904), .B(n891), .Y(n365) );
  INVX1 U667 ( .A(n365), .Y(n685) );
  OR2X1 U668 ( .A(n920), .B(n902), .Y(n323) );
  INVX1 U669 ( .A(n323), .Y(n686) );
  OR2X2 U670 ( .A(n663), .B(n819), .Y(n294) );
  INVX1 U671 ( .A(n294), .Y(n687) );
  INVX1 U672 ( .A(n344), .Y(n688) );
  BUFX2 U673 ( .A(n358), .Y(n689) );
  BUFX2 U674 ( .A(n327), .Y(n690) );
  BUFX2 U675 ( .A(n314), .Y(n691) );
  BUFX2 U676 ( .A(n302), .Y(n692) );
  BUFX2 U677 ( .A(n287), .Y(n693) );
  BUFX2 U678 ( .A(n176), .Y(n694) );
  BUFX2 U679 ( .A(n164), .Y(n695) );
  BUFX2 U680 ( .A(n147), .Y(n696) );
  AND2X1 U681 ( .A(n878), .B(n374), .Y(n59) );
  INVX1 U682 ( .A(n59), .Y(n697) );
  AND2X1 U683 ( .A(n840), .B(n361), .Y(n56) );
  INVX1 U684 ( .A(n56), .Y(n698) );
  AND2X1 U685 ( .A(n761), .B(n348), .Y(n53) );
  INVX1 U686 ( .A(n53), .Y(n699) );
  AND2X1 U687 ( .A(n841), .B(n330), .Y(n50) );
  INVX1 U688 ( .A(n50), .Y(n700) );
  AND2X1 U689 ( .A(n843), .B(n305), .Y(n46) );
  INVX1 U690 ( .A(n46), .Y(n701) );
  AND2X1 U691 ( .A(n892), .B(n290), .Y(n44) );
  INVX1 U692 ( .A(n44), .Y(n702) );
  AND2X1 U693 ( .A(n764), .B(n277), .Y(n41) );
  INVX1 U694 ( .A(n41), .Y(n703) );
  AND2X1 U695 ( .A(n872), .B(n267), .Y(n40) );
  INVX1 U696 ( .A(n40), .Y(n704) );
  AND2X1 U697 ( .A(n765), .B(n264), .Y(n39) );
  INVX1 U698 ( .A(n39), .Y(n705) );
  AND2X1 U699 ( .A(n766), .B(n256), .Y(n37) );
  INVX1 U700 ( .A(n37), .Y(n706) );
  AND2X1 U701 ( .A(n874), .B(n246), .Y(n36) );
  INVX1 U702 ( .A(n36), .Y(n707) );
  AND2X1 U703 ( .A(n767), .B(n243), .Y(n35) );
  INVX1 U704 ( .A(n35), .Y(n708) );
  AND2X1 U705 ( .A(n768), .B(n235), .Y(n33) );
  INVX1 U706 ( .A(n33), .Y(n709) );
  AND2X1 U707 ( .A(n876), .B(n225), .Y(n32) );
  INVX1 U708 ( .A(n32), .Y(n710) );
  AND2X1 U709 ( .A(n769), .B(n408), .Y(n31) );
  INVX1 U710 ( .A(n31), .Y(n711) );
  AND2X1 U711 ( .A(n770), .B(n214), .Y(n29) );
  INVX1 U712 ( .A(n29), .Y(n712) );
  AND2X1 U713 ( .A(n771), .B(n199), .Y(n27) );
  INVX1 U714 ( .A(n27), .Y(n713) );
  AND2X1 U715 ( .A(n845), .B(n399), .Y(n22) );
  INVX1 U716 ( .A(n22), .Y(n714) );
  INVX1 U717 ( .A(n17), .Y(n715) );
  AND2X1 U718 ( .A(n776), .B(n124), .Y(n16) );
  INVX1 U719 ( .A(n16), .Y(n716) );
  AND2X1 U720 ( .A(n748), .B(n926), .Y(n12) );
  INVX1 U721 ( .A(n12), .Y(n717) );
  AND2X1 U722 ( .A(n749), .B(n931), .Y(n10) );
  INVX1 U723 ( .A(n10), .Y(n718) );
  AND2X1 U724 ( .A(n750), .B(n934), .Y(n6) );
  INVX1 U725 ( .A(n6), .Y(n719) );
  AND2X1 U726 ( .A(n760), .B(n356), .Y(n55) );
  INVX1 U727 ( .A(n55), .Y(n720) );
  AND2X1 U728 ( .A(n870), .B(n351), .Y(n54) );
  INVX1 U729 ( .A(n54), .Y(n721) );
  AND2X1 U730 ( .A(n842), .B(n317), .Y(n48) );
  INVX1 U731 ( .A(n48), .Y(n722) );
  AND2X1 U732 ( .A(n762), .B(n312), .Y(n47) );
  INVX1 U733 ( .A(n47), .Y(n723) );
  AND2X1 U734 ( .A(n763), .B(n300), .Y(n45) );
  INVX1 U735 ( .A(n45), .Y(n724) );
  AND2X1 U736 ( .A(n887), .B(n285), .Y(n43) );
  INVX1 U737 ( .A(n43), .Y(n725) );
  AND2X1 U738 ( .A(n871), .B(n280), .Y(n42) );
  INVX1 U739 ( .A(n42), .Y(n726) );
  AND2X1 U740 ( .A(n873), .B(n259), .Y(n38) );
  INVX1 U741 ( .A(n38), .Y(n727) );
  AND2X1 U742 ( .A(n875), .B(n238), .Y(n34) );
  INVX1 U743 ( .A(n34), .Y(n728) );
  AND2X1 U744 ( .A(n877), .B(n217), .Y(n30) );
  INVX1 U745 ( .A(n30), .Y(n729) );
  AND2X1 U746 ( .A(n844), .B(n179), .Y(n24) );
  INVX1 U747 ( .A(n24), .Y(n730) );
  AND2X1 U748 ( .A(n772), .B(n400), .Y(n23) );
  INVX1 U749 ( .A(n23), .Y(n731) );
  AND2X1 U750 ( .A(n773), .B(n162), .Y(n21) );
  INVX1 U751 ( .A(n21), .Y(n732) );
  INVX1 U752 ( .A(n20), .Y(n733) );
  AND2X1 U753 ( .A(n774), .B(n396), .Y(n19) );
  INVX1 U754 ( .A(n19), .Y(n734) );
  AND2X1 U755 ( .A(n777), .B(n119), .Y(n15) );
  INVX1 U756 ( .A(n15), .Y(n735) );
  AND2X1 U757 ( .A(n778), .B(n111), .Y(n13) );
  INVX1 U758 ( .A(n13), .Y(n736) );
  AND2X1 U759 ( .A(n779), .B(n103), .Y(n11) );
  INVX1 U760 ( .A(n11), .Y(n737) );
  AND2X1 U761 ( .A(n780), .B(n95), .Y(n9) );
  INVX1 U762 ( .A(n9), .Y(n738) );
  AND2X1 U763 ( .A(n781), .B(n87), .Y(n7) );
  INVX1 U764 ( .A(n7), .Y(n739) );
  AND2X1 U765 ( .A(n782), .B(n79), .Y(n5) );
  INVX1 U766 ( .A(n5), .Y(n740) );
  AND2X1 U767 ( .A(n783), .B(n71), .Y(n3) );
  INVX1 U768 ( .A(n3), .Y(n741) );
  INVX1 U769 ( .A(n172), .Y(n742) );
  INVX1 U770 ( .A(n69), .Y(n743) );
  INVX1 U771 ( .A(n143), .Y(n744) );
  INVX1 U772 ( .A(n241), .Y(n745) );
  INVX1 U773 ( .A(n310), .Y(n746) );
  OR2X1 U774 ( .A(n912), .B(n868), .Y(n197) );
  INVX1 U775 ( .A(n197), .Y(n747) );
  INVX1 U776 ( .A(n109), .Y(n748) );
  AND2X1 U777 ( .A(B[50]), .B(A[50]), .Y(n101) );
  INVX1 U778 ( .A(n101), .Y(n749) );
  AND2X1 U779 ( .A(B[54]), .B(A[54]), .Y(n85) );
  INVX1 U780 ( .A(n85), .Y(n750) );
  INVX1 U781 ( .A(n179), .Y(n751) );
  AND2X1 U782 ( .A(B[11]), .B(A[11]), .Y(n326) );
  INVX1 U783 ( .A(n326), .Y(n752) );
  AND2X1 U784 ( .A(A[35]), .B(B[35]), .Y(n188) );
  INVX1 U785 ( .A(n188), .Y(n753) );
  OR2X1 U786 ( .A(B[4]), .B(A[4]), .Y(n361) );
  INVX1 U787 ( .A(n361), .Y(n754) );
  OR2X1 U788 ( .A(A[14]), .B(B[14]), .Y(n305) );
  INVX1 U789 ( .A(n305), .Y(n755) );
  INVX1 U790 ( .A(n290), .Y(n756) );
  OR2X1 U791 ( .A(A[12]), .B(B[12]), .Y(n317) );
  INVX1 U792 ( .A(n317), .Y(n757) );
  INVX1 U793 ( .A(n651), .Y(n758) );
  INVX1 U794 ( .A(n150), .Y(n759) );
  INVX1 U795 ( .A(n357), .Y(n760) );
  AND2X1 U796 ( .A(B[7]), .B(A[7]), .Y(n349) );
  INVX1 U797 ( .A(n349), .Y(n761) );
  AND2X1 U798 ( .A(B[13]), .B(A[13]), .Y(n313) );
  INVX1 U799 ( .A(n313), .Y(n762) );
  INVX1 U800 ( .A(n301), .Y(n763) );
  AND2X1 U801 ( .A(B[19]), .B(A[19]), .Y(n278) );
  INVX1 U802 ( .A(n278), .Y(n764) );
  INVX1 U803 ( .A(n265), .Y(n765) );
  AND2X1 U804 ( .A(B[23]), .B(A[23]), .Y(n257) );
  INVX1 U805 ( .A(n257), .Y(n766) );
  INVX1 U806 ( .A(n244), .Y(n767) );
  INVX1 U807 ( .A(n236), .Y(n768) );
  INVX1 U808 ( .A(n223), .Y(n769) );
  INVX1 U809 ( .A(n215), .Y(n770) );
  AND2X1 U810 ( .A(A[33]), .B(B[33]), .Y(n200) );
  INVX1 U811 ( .A(n200), .Y(n771) );
  INVX1 U812 ( .A(n175), .Y(n772) );
  INVX1 U813 ( .A(n163), .Y(n773) );
  INVX1 U814 ( .A(n132), .Y(n775) );
  INVX1 U815 ( .A(n125), .Y(n776) );
  INVX1 U816 ( .A(n120), .Y(n777) );
  AND2X1 U817 ( .A(B[47]), .B(A[47]), .Y(n112) );
  INVX1 U818 ( .A(n112), .Y(n778) );
  INVX1 U819 ( .A(n104), .Y(n779) );
  INVX1 U820 ( .A(n96), .Y(n780) );
  INVX1 U821 ( .A(n88), .Y(n781) );
  INVX1 U822 ( .A(n80), .Y(n782) );
  INVX1 U823 ( .A(n72), .Y(n783) );
  INVX1 U824 ( .A(n119), .Y(n784) );
  OR2X1 U825 ( .A(A[47]), .B(B[47]), .Y(n111) );
  INVX1 U826 ( .A(n111), .Y(n785) );
  INVX1 U827 ( .A(n87), .Y(n786) );
  INVX1 U828 ( .A(n79), .Y(n787) );
  BUFX2 U829 ( .A(n322), .Y(n788) );
  BUFX2 U830 ( .A(n364), .Y(n789) );
  INVX1 U831 ( .A(n791), .Y(n790) );
  BUFX2 U832 ( .A(n274), .Y(n791) );
  BUFX2 U833 ( .A(n270), .Y(n792) );
  BUFX2 U834 ( .A(n249), .Y(n793) );
  INVX1 U835 ( .A(n795), .Y(n794) );
  BUFX2 U836 ( .A(n232), .Y(n795) );
  BUFX2 U837 ( .A(n228), .Y(n796) );
  INVX1 U838 ( .A(n262), .Y(n797) );
  INVX1 U839 ( .A(n220), .Y(n798) );
  INVX1 U840 ( .A(n129), .Y(n799) );
  OR2X1 U841 ( .A(n854), .B(n863), .Y(n254) );
  INVX1 U842 ( .A(n254), .Y(n800) );
  INVX1 U843 ( .A(n212), .Y(n801) );
  INVX1 U844 ( .A(n354), .Y(n802) );
  OR2X2 U845 ( .A(n852), .B(n755), .Y(n298) );
  INVX1 U846 ( .A(n298), .Y(n803) );
  OR2X1 U847 ( .A(n906), .B(n915), .Y(n275) );
  INVX1 U848 ( .A(n275), .Y(n804) );
  INVX1 U849 ( .A(n233), .Y(n805) );
  INVX1 U850 ( .A(n208), .Y(n806) );
  OR2X2 U851 ( .A(n664), .B(n816), .Y(n208) );
  INVX1 U852 ( .A(n185), .Y(n807) );
  OR2X1 U853 ( .A(n850), .B(n861), .Y(n346) );
  INVX1 U854 ( .A(n346), .Y(n808) );
  INVX1 U855 ( .A(n283), .Y(n809) );
  INVX1 U856 ( .A(n250), .Y(n810) );
  BUFX2 U857 ( .A(n668), .Y(n811) );
  BUFX2 U858 ( .A(n135), .Y(n812) );
  INVX1 U859 ( .A(n128), .Y(n813) );
  INVX1 U860 ( .A(n813), .Y(n814) );
  INVX1 U861 ( .A(n252), .Y(n815) );
  AND2X2 U862 ( .A(n798), .B(n801), .Y(n210) );
  INVX1 U863 ( .A(n210), .Y(n816) );
  INVX1 U864 ( .A(n134), .Y(n817) );
  AND2X2 U865 ( .A(n666), .B(n799), .Y(n127) );
  INVX1 U866 ( .A(n127), .Y(n818) );
  INVX1 U867 ( .A(n321), .Y(n819) );
  AND2X2 U868 ( .A(n742), .B(n677), .Y(n158) );
  BUFX2 U869 ( .A(n353), .Y(n821) );
  BUFX2 U870 ( .A(n282), .Y(n822) );
  BUFX2 U871 ( .A(n261), .Y(n823) );
  BUFX2 U872 ( .A(n240), .Y(n824) );
  BUFX2 U873 ( .A(n219), .Y(n825) );
  INVX1 U874 ( .A(n121), .Y(n826) );
  INVX1 U875 ( .A(n826), .Y(n827) );
  INVX1 U876 ( .A(n826), .Y(n828) );
  INVX1 U877 ( .A(n113), .Y(n829) );
  INVX1 U878 ( .A(n654), .Y(n830) );
  INVX1 U879 ( .A(n829), .Y(n831) );
  INVX1 U880 ( .A(n97), .Y(n832) );
  INVX1 U881 ( .A(n656), .Y(n833) );
  INVX1 U882 ( .A(n832), .Y(n834) );
  INVX1 U883 ( .A(n89), .Y(n835) );
  INVX1 U884 ( .A(n835), .Y(n836) );
  INVX1 U885 ( .A(n81), .Y(n837) );
  INVX1 U886 ( .A(n837), .Y(n838) );
  BUFX2 U887 ( .A(n673), .Y(n839) );
  INVX1 U888 ( .A(n362), .Y(n840) );
  AND2X1 U889 ( .A(A[4]), .B(B[4]), .Y(n362) );
  INVX1 U890 ( .A(n331), .Y(n841) );
  AND2X1 U891 ( .A(A[10]), .B(B[10]), .Y(n331) );
  INVX1 U892 ( .A(n318), .Y(n842) );
  AND2X1 U893 ( .A(B[12]), .B(A[12]), .Y(n318) );
  INVX1 U894 ( .A(n306), .Y(n843) );
  INVX1 U895 ( .A(n180), .Y(n844) );
  INVX1 U896 ( .A(n168), .Y(n845) );
  INVX1 U897 ( .A(n203), .Y(n847) );
  INVX1 U898 ( .A(n203), .Y(n848) );
  INVX1 U899 ( .A(n356), .Y(n849) );
  INVX1 U900 ( .A(n348), .Y(n850) );
  OR2X1 U901 ( .A(A[7]), .B(B[7]), .Y(n348) );
  INVX1 U902 ( .A(n312), .Y(n851) );
  OR2X1 U903 ( .A(A[13]), .B(B[13]), .Y(n312) );
  INVX1 U904 ( .A(n300), .Y(n852) );
  OR2X1 U905 ( .A(A[15]), .B(B[15]), .Y(n300) );
  INVX1 U906 ( .A(n264), .Y(n853) );
  INVX1 U907 ( .A(n256), .Y(n854) );
  INVX1 U908 ( .A(n243), .Y(n855) );
  INVX1 U909 ( .A(n235), .Y(n856) );
  OR2X1 U910 ( .A(A[29]), .B(B[29]), .Y(n222) );
  INVX1 U911 ( .A(n222), .Y(n857) );
  INVX1 U912 ( .A(n214), .Y(n858) );
  INVX1 U913 ( .A(n162), .Y(n859) );
  INVX1 U914 ( .A(n351), .Y(n861) );
  INVX1 U915 ( .A(n267), .Y(n862) );
  INVX1 U916 ( .A(n259), .Y(n863) );
  OR2X1 U917 ( .A(A[22]), .B(B[22]), .Y(n259) );
  INVX1 U918 ( .A(n246), .Y(n864) );
  OR2X1 U919 ( .A(A[24]), .B(B[24]), .Y(n246) );
  OR2X1 U920 ( .A(A[26]), .B(B[26]), .Y(n238) );
  INVX1 U921 ( .A(n238), .Y(n865) );
  INVX1 U922 ( .A(n225), .Y(n866) );
  INVX1 U923 ( .A(n217), .Y(n867) );
  INVX1 U924 ( .A(n199), .Y(n868) );
  OR2X1 U925 ( .A(B[33]), .B(A[33]), .Y(n199) );
  INVX1 U926 ( .A(n174), .Y(n869) );
  INVX1 U927 ( .A(n352), .Y(n870) );
  INVX1 U928 ( .A(n281), .Y(n871) );
  INVX1 U929 ( .A(n268), .Y(n872) );
  AND2X1 U930 ( .A(B[22]), .B(A[22]), .Y(n260) );
  INVX1 U931 ( .A(n260), .Y(n873) );
  AND2X1 U932 ( .A(B[24]), .B(A[24]), .Y(n247) );
  INVX1 U933 ( .A(n247), .Y(n874) );
  AND2X1 U934 ( .A(B[26]), .B(A[26]), .Y(n239) );
  INVX1 U935 ( .A(n239), .Y(n875) );
  AND2X1 U936 ( .A(B[28]), .B(A[28]), .Y(n226) );
  INVX1 U937 ( .A(n226), .Y(n876) );
  INVX1 U938 ( .A(n218), .Y(n877) );
  OR2X2 U939 ( .A(A[58]), .B(B[58]), .Y(n930) );
  INVX1 U940 ( .A(n375), .Y(n878) );
  AND2X1 U941 ( .A(n919), .B(n932), .Y(SUM[0]) );
  AND2X1 U942 ( .A(n886), .B(n367), .Y(n57) );
  INVX1 U943 ( .A(n57), .Y(n879) );
  INVX1 U944 ( .A(n374), .Y(n880) );
  AND2X1 U945 ( .A(n888), .B(n337), .Y(n51) );
  INVX1 U946 ( .A(n51), .Y(n881) );
  INVX1 U947 ( .A(n25), .Y(n882) );
  BUFX2 U948 ( .A(n189), .Y(n883) );
  OR2X1 U949 ( .A(n893), .B(n913), .Y(n335) );
  INVX1 U950 ( .A(n335), .Y(n884) );
  INVX1 U951 ( .A(n192), .Y(n885) );
  AND2X1 U952 ( .A(A[3]), .B(B[3]), .Y(n368) );
  INVX1 U953 ( .A(n368), .Y(n886) );
  INVX1 U954 ( .A(n286), .Y(n887) );
  INVX1 U955 ( .A(n338), .Y(n888) );
  AND2X1 U956 ( .A(n903), .B(n403), .Y(n26) );
  INVX1 U957 ( .A(n26), .Y(n889) );
  AND2X1 U958 ( .A(n907), .B(n340), .Y(n52) );
  INVX1 U959 ( .A(n52), .Y(n890) );
  INVX1 U960 ( .A(n370), .Y(n891) );
  INVX1 U961 ( .A(n291), .Y(n892) );
  INVX1 U962 ( .A(n337), .Y(n893) );
  INVX1 U963 ( .A(n2), .Y(n894) );
  AND2X1 U964 ( .A(n918), .B(n370), .Y(n58) );
  INVX1 U965 ( .A(n58), .Y(n895) );
  INVX1 U966 ( .A(n49), .Y(n896) );
  INVX1 U967 ( .A(n28), .Y(n897) );
  AND2X1 U968 ( .A(B[46]), .B(A[46]), .Y(n117) );
  INVX1 U969 ( .A(n117), .Y(n898) );
  INVX1 U970 ( .A(n77), .Y(n899) );
  INVX1 U971 ( .A(n139), .Y(n900) );
  INVX1 U972 ( .A(n93), .Y(n901) );
  INVX1 U973 ( .A(n330), .Y(n902) );
  AND2X1 U974 ( .A(A[34]), .B(B[34]), .Y(n193) );
  INVX1 U975 ( .A(n193), .Y(n903) );
  OR2X1 U976 ( .A(B[3]), .B(A[3]), .Y(n367) );
  INVX1 U977 ( .A(n367), .Y(n904) );
  INVX1 U978 ( .A(n285), .Y(n905) );
  AND2X1 U979 ( .A(B[8]), .B(A[8]), .Y(n341) );
  INVX1 U980 ( .A(n341), .Y(n907) );
  INVX1 U981 ( .A(n14), .Y(n908) );
  INVX1 U982 ( .A(n18), .Y(n909) );
  INVX1 U983 ( .A(n8), .Y(n910) );
  INVX1 U984 ( .A(n4), .Y(n911) );
  INVX1 U985 ( .A(n202), .Y(n912) );
  OR2X1 U986 ( .A(A[8]), .B(B[8]), .Y(n340) );
  INVX1 U987 ( .A(n340), .Y(n913) );
  INVX1 U988 ( .A(n124), .Y(n914) );
  INVX1 U989 ( .A(n280), .Y(n915) );
  OR2X1 U990 ( .A(A[43]), .B(B[43]), .Y(n131) );
  INVX1 U991 ( .A(n131), .Y(n916) );
  INVX1 U992 ( .A(n371), .Y(n918) );
  AND2X1 U993 ( .A(A[0]), .B(B[0]), .Y(n377) );
  OR2X1 U994 ( .A(A[11]), .B(B[11]), .Y(n325) );
  INVX1 U995 ( .A(n325), .Y(n920) );
  BUFX2 U996 ( .A(n94), .Y(n921) );
  BUFX2 U997 ( .A(n118), .Y(n922) );
  BUFX2 U998 ( .A(n78), .Y(n923) );
  BUFX2 U999 ( .A(n86), .Y(n924) );
  BUFX2 U1000 ( .A(n891), .Y(n925) );
  INVX1 U1001 ( .A(n182), .Y(n181) );
  INVX1 U1002 ( .A(n792), .Y(n269) );
  INVX1 U1003 ( .A(n153), .Y(n152) );
  INVX1 U1004 ( .A(n320), .Y(n319) );
  INVX1 U1005 ( .A(n793), .Y(n248) );
  INVX1 U1006 ( .A(n796), .Y(n227) );
  INVX1 U1007 ( .A(n373), .Y(n372) );
  INVX1 U1008 ( .A(n789), .Y(n363) );
  INVX1 U1009 ( .A(n640), .Y(n142) );
  INVX1 U1010 ( .A(n885), .Y(n403) );
  INVX1 U1011 ( .A(n311), .Y(n309) );
  INVX1 U1012 ( .A(n173), .Y(n171) );
  INVX1 U1013 ( .A(n742), .Y(n170) );
  INVX1 U1014 ( .A(n198), .Y(n196) );
  INVX1 U1015 ( .A(n642), .Y(n155) );
  INVX1 U1016 ( .A(n343), .Y(n342) );
  INVX1 U1017 ( .A(n860), .Y(n396) );
  INVX1 U1018 ( .A(n758), .Y(n399) );
  INVX1 U1019 ( .A(n759), .Y(n397) );
  OR2X1 U1020 ( .A(A[46]), .B(B[46]), .Y(n928) );
  INVX1 U1021 ( .A(n869), .Y(n400) );
  OR2X1 U1022 ( .A(B[0]), .B(A[0]), .Y(n932) );
  OR2X1 U1023 ( .A(A[52]), .B(B[52]), .Y(n933) );
  OR2X1 U1024 ( .A(A[54]), .B(B[54]), .Y(n934) );
  BUFX2 U1025 ( .A(n110), .Y(n935) );
  INVX1 U1026 ( .A(n857), .Y(n408) );
  INVX1 U1027 ( .A(n65), .Y(n378) );
  INVX1 U1028 ( .A(n675), .Y(n292) );
  INVX1 U1029 ( .A(n638), .Y(n204) );
  INVX1 U1030 ( .A(n336), .Y(n334) );
endmodule


module alu_DW_mult_uns_37 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n2, n8, n12, n14, n18, n20, n24, n26, n30, n32, n36, n38, n42, n44,
         n48, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n115, n116, n120, n121, n122, n123, n124,
         n128, n129, n130, n131, n132, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n148, n149, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n164, n165, n166, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n213, n214, n218, n219, n220, n224, n225, n226, n227,
         n231, n232, n236, n237, n238, n242, n243, n244, n245, n246, n250,
         n251, n252, n253, n254, n258, n259, n260, n261, n262, n263, n277,
         n278, n293, n294, n295, n296, n297, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n576,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n595, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n614, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n633, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n652, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n671, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n690, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n709, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n728, n729, n731, n733, n735, n737, n739, n741,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226;

  XOR2X1 U85 ( .A(n115), .B(n85), .Y(product[31]) );
  XOR2X1 U86 ( .A(n295), .B(n294), .Y(n85) );
  FAX1 U87 ( .A(n296), .B(n299), .C(n263), .YC(n115), .YS(product[30]) );
  XNOR2X1 U89 ( .A(n121), .B(n1073), .Y(product[29]) );
  AOI21X1 U90 ( .A(n121), .B(n1153), .C(n120), .Y(n116) );
  XOR2X1 U97 ( .A(n1038), .B(n1028), .Y(product[28]) );
  OAI21X1 U98 ( .A(n1130), .B(n1039), .C(n1113), .Y(n121) );
  XNOR2X1 U103 ( .A(n129), .B(n1126), .Y(product[27]) );
  AOI21X1 U104 ( .A(n129), .B(n1150), .C(n128), .Y(n124) );
  XOR2X1 U111 ( .A(n1036), .B(n1074), .Y(product[26]) );
  OAI21X1 U112 ( .A(n1006), .B(n1132), .C(n1112), .Y(n129) );
  XNOR2X1 U117 ( .A(n137), .B(n1023), .Y(product[25]) );
  AOI21X1 U118 ( .A(n137), .B(n1151), .C(n136), .Y(n132) );
  XOR2X1 U125 ( .A(n1034), .B(n1027), .Y(product[24]) );
  OAI21X1 U126 ( .A(n1134), .B(n1035), .C(n1116), .Y(n137) );
  XOR2X1 U131 ( .A(n1019), .B(n1026), .Y(product[23]) );
  AOI21X1 U132 ( .A(n177), .B(n1004), .C(n142), .Y(n140) );
  OAI21X1 U134 ( .A(n1032), .B(n1031), .C(n1013), .Y(n142) );
  AOI21X1 U136 ( .A(n1145), .B(n153), .C(n148), .Y(n144) );
  XNOR2X1 U143 ( .A(n154), .B(n1022), .Y(product[22]) );
  AOI21X1 U144 ( .A(n154), .B(n1144), .C(n153), .Y(n149) );
  XOR2X1 U151 ( .A(n1062), .B(n1061), .Y(product[21]) );
  OAI21X1 U152 ( .A(n1003), .B(n176), .C(n1031), .Y(n154) );
  AOI21X1 U154 ( .A(n170), .B(n1002), .C(n158), .Y(n156) );
  OAI21X1 U156 ( .A(n1101), .B(n1136), .C(n1115), .Y(n158) );
  XNOR2X1 U161 ( .A(n166), .B(n1021), .Y(product[20]) );
  AOI21X1 U162 ( .A(n166), .B(n164), .C(n165), .Y(n161) );
  XNOR2X1 U169 ( .A(n173), .B(n1090), .Y(product[19]) );
  OAI21X1 U170 ( .A(n169), .B(n176), .C(n168), .Y(n166) );
  OAI21X1 U174 ( .A(n1137), .B(n1121), .C(n1065), .Y(n170) );
  XOR2X1 U179 ( .A(n176), .B(n1108), .Y(product[18]) );
  OAI21X1 U180 ( .A(n1081), .B(n176), .C(n1137), .Y(n173) );
  XNOR2X1 U185 ( .A(n184), .B(n1050), .Y(product[17]) );
  OAI21X1 U187 ( .A(n1008), .B(n1001), .C(n1012), .Y(n177) );
  AOI21X1 U189 ( .A(n1079), .B(n189), .C(n181), .Y(n179) );
  OAI21X1 U191 ( .A(n1139), .B(n1103), .C(n1057), .Y(n181) );
  XOR2X1 U196 ( .A(n1080), .B(n1092), .Y(product[16]) );
  OAI21X1 U197 ( .A(n1120), .B(n1080), .C(n1139), .Y(n184) );
  XOR2X1 U202 ( .A(n1056), .B(n1055), .Y(product[15]) );
  AOI21X1 U203 ( .A(n197), .B(n1067), .C(n189), .Y(n187) );
  OAI21X1 U205 ( .A(n1135), .B(n1104), .C(n1066), .Y(n189) );
  XNOR2X1 U210 ( .A(n197), .B(n1088), .Y(product[14]) );
  AOI21X1 U211 ( .A(n197), .B(n195), .C(n196), .Y(n192) );
  XNOR2X1 U218 ( .A(n203), .B(n1060), .Y(product[13]) );
  AOI21X1 U220 ( .A(n1014), .B(n207), .C(n200), .Y(n198) );
  OAI21X1 U222 ( .A(n1138), .B(n1102), .C(n1078), .Y(n200) );
  XOR2X1 U227 ( .A(n206), .B(n1091), .Y(product[12]) );
  OAI21X1 U228 ( .A(n1119), .B(n206), .C(n1138), .Y(n203) );
  XOR2X1 U233 ( .A(n1018), .B(n1025), .Y(product[11]) );
  OAI21X1 U235 ( .A(n1005), .B(n1015), .C(n1010), .Y(n207) );
  AOI21X1 U237 ( .A(n1149), .B(n218), .C(n213), .Y(n209) );
  XNOR2X1 U244 ( .A(n219), .B(n1089), .Y(product[10]) );
  AOI21X1 U245 ( .A(n219), .B(n1147), .C(n218), .Y(n214) );
  XNOR2X1 U252 ( .A(n225), .B(n1087), .Y(product[9]) );
  AOI21X1 U254 ( .A(n225), .B(n1152), .C(n224), .Y(n220) );
  XOR2X1 U261 ( .A(n1017), .B(n1024), .Y(product[8]) );
  OAI21X1 U262 ( .A(n1007), .B(n1000), .C(n1009), .Y(n225) );
  AOI21X1 U264 ( .A(n1148), .B(n236), .C(n231), .Y(n227) );
  XNOR2X1 U271 ( .A(n237), .B(n1020), .Y(product[7]) );
  AOI21X1 U272 ( .A(n237), .B(n1146), .C(n236), .Y(n232) );
  XNOR2X1 U279 ( .A(n1070), .B(n243), .Y(product[6]) );
  AOI21X1 U281 ( .A(n243), .B(n1155), .C(n242), .Y(n238) );
  XOR2X1 U288 ( .A(n1072), .B(n1100), .Y(product[5]) );
  OAI21X1 U289 ( .A(n1131), .B(n1100), .C(n1114), .Y(n243) );
  XNOR2X1 U294 ( .A(n1053), .B(n251), .Y(product[4]) );
  AOI21X1 U295 ( .A(n251), .B(n1156), .C(n250), .Y(n246) );
  XOR2X1 U302 ( .A(n1054), .B(n1118), .Y(product[3]) );
  OAI21X1 U303 ( .A(n1133), .B(n1118), .C(n1077), .Y(n251) );
  XNOR2X1 U308 ( .A(n1071), .B(n1099), .Y(product[2]) );
  AOI21X1 U309 ( .A(n1154), .B(n1099), .C(n258), .Y(n254) );
  XOR2X1 U316 ( .A(n260), .B(n1141), .Y(product[1]) );
  XOR2X1 U324 ( .A(n761), .B(n293), .Y(n294) );
  FAX1 U326 ( .A(n297), .B(n762), .C(n301), .YC(n295), .YS(n296) );
  FAX1 U328 ( .A(n763), .B(n302), .C(n305), .YC(n299), .YS(n300) );
  FAX1 U329 ( .A(n779), .B(n1068), .C(n1042), .YC(n301), .YS(n302) );
  FAX1 U330 ( .A(n313), .B(n306), .C(n311), .YC(n303), .YS(n304) );
  FAX1 U331 ( .A(n307), .B(n780), .C(n764), .YC(n305), .YS(n306) );
  FAX1 U333 ( .A(n319), .B(n312), .C(n317), .YC(n309), .YS(n310) );
  FAX1 U334 ( .A(n781), .B(n765), .C(n314), .YC(n311), .YS(n312) );
  FAX1 U335 ( .A(n797), .B(n1105), .C(n1044), .YC(n313), .YS(n314) );
  FAX1 U336 ( .A(n327), .B(n318), .C(n325), .YC(n315), .YS(n316) );
  FAX1 U337 ( .A(n766), .B(n329), .C(n320), .YC(n317), .YS(n318) );
  FAX1 U338 ( .A(n321), .B(n798), .C(n782), .YC(n319), .YS(n320) );
  FAX1 U340 ( .A(n328), .B(n326), .C(n333), .YC(n323), .YS(n324) );
  FAX1 U341 ( .A(n330), .B(n337), .C(n335), .YC(n325), .YS(n326) );
  FAX1 U342 ( .A(n783), .B(n799), .C(n767), .YC(n327), .YS(n328) );
  FAX1 U343 ( .A(n815), .B(n1082), .C(n1043), .YC(n329), .YS(n330) );
  FAX1 U344 ( .A(n345), .B(n334), .C(n343), .YC(n331), .YS(n332) );
  FAX1 U345 ( .A(n338), .B(n347), .C(n336), .YC(n333), .YS(n334) );
  FAX1 U346 ( .A(n800), .B(n768), .C(n349), .YC(n335), .YS(n336) );
  FAX1 U347 ( .A(n339), .B(n816), .C(n784), .YC(n337), .YS(n338) );
  FAX1 U349 ( .A(n355), .B(n344), .C(n353), .YC(n341), .YS(n342) );
  FAX1 U350 ( .A(n357), .B(n348), .C(n346), .YC(n343), .YS(n344) );
  FAX1 U351 ( .A(n785), .B(n350), .C(n359), .YC(n345), .YS(n346) );
  FAX1 U352 ( .A(n817), .B(n801), .C(n769), .YC(n347), .YS(n348) );
  FAX1 U353 ( .A(n833), .B(n1122), .C(n1045), .YC(n349), .YS(n350) );
  FAX1 U354 ( .A(n367), .B(n354), .C(n365), .YC(n351), .YS(n352) );
  FAX1 U355 ( .A(n369), .B(n358), .C(n356), .YC(n353), .YS(n354) );
  FAX1 U356 ( .A(n802), .B(n360), .C(n371), .YC(n355), .YS(n356) );
  FAX1 U357 ( .A(n786), .B(n770), .C(n373), .YC(n357), .YS(n358) );
  FAX1 U358 ( .A(n361), .B(n834), .C(n818), .YC(n359), .YS(n360) );
  FAX1 U360 ( .A(n368), .B(n377), .C(n366), .YC(n363), .YS(n364) );
  FAX1 U361 ( .A(n370), .B(n381), .C(n379), .YC(n365), .YS(n366) );
  FAX1 U362 ( .A(n385), .B(n383), .C(n372), .YC(n367), .YS(n368) );
  FAX1 U363 ( .A(n787), .B(n835), .C(n374), .YC(n369), .YS(n370) );
  FAX1 U364 ( .A(n819), .B(n803), .C(n771), .YC(n371), .YS(n372) );
  FAX1 U365 ( .A(n851), .B(n1140), .C(n1046), .YC(n373), .YS(n374) );
  FAX1 U366 ( .A(n380), .B(n391), .C(n378), .YC(n375), .YS(n376) );
  FAX1 U367 ( .A(n382), .B(n395), .C(n393), .YC(n377), .YS(n378) );
  FAX1 U368 ( .A(n399), .B(n397), .C(n384), .YC(n379), .YS(n380) );
  FAX1 U369 ( .A(n836), .B(n804), .C(n386), .YC(n381), .YS(n382) );
  FAX1 U370 ( .A(n788), .B(n772), .C(n401), .YC(n383), .YS(n384) );
  FAX1 U371 ( .A(n387), .B(n852), .C(n820), .YC(n385), .YS(n386) );
  FAX1 U373 ( .A(n394), .B(n405), .C(n392), .YC(n389), .YS(n390) );
  FAX1 U374 ( .A(n409), .B(n396), .C(n407), .YC(n391), .YS(n392) );
  FAX1 U375 ( .A(n411), .B(n400), .C(n398), .YC(n393), .YS(n394) );
  FAX1 U376 ( .A(n789), .B(n415), .C(n413), .YC(n395), .YS(n396) );
  FAX1 U377 ( .A(n853), .B(n837), .C(n805), .YC(n397), .YS(n398) );
  FAX1 U378 ( .A(n821), .B(n773), .C(n402), .YC(n399), .YS(n400) );
  FAX1 U379 ( .A(n1211), .B(n1143), .C(n1047), .YC(n401), .YS(n402) );
  FAX1 U380 ( .A(n408), .B(n421), .C(n406), .YC(n403), .YS(n404) );
  FAX1 U381 ( .A(n425), .B(n410), .C(n423), .YC(n405), .YS(n406) );
  FAX1 U382 ( .A(n427), .B(n414), .C(n412), .YC(n407), .YS(n408) );
  FAX1 U383 ( .A(n416), .B(n431), .C(n429), .YC(n409), .YS(n410) );
  FAX1 U384 ( .A(n854), .B(n790), .C(n838), .YC(n411), .YS(n412) );
  FAX1 U385 ( .A(n822), .B(n806), .C(n774), .YC(n413), .YS(n414) );
  FAX1 U386 ( .A(n1210), .B(n1117), .C(n870), .YC(n415), .YS(n416) );
  FAX1 U388 ( .A(n424), .B(n436), .C(n422), .YC(n419), .YS(n420) );
  FAX1 U389 ( .A(n440), .B(n426), .C(n438), .YC(n421), .YS(n422) );
  FAX1 U390 ( .A(n444), .B(n430), .C(n428), .YC(n423), .YS(n424) );
  FAX1 U391 ( .A(n446), .B(n432), .C(n442), .YC(n425), .YS(n426) );
  FAX1 U392 ( .A(n855), .B(n791), .C(n839), .YC(n427), .YS(n428) );
  FAX1 U393 ( .A(n823), .B(n807), .C(n775), .YC(n429), .YS(n430) );
  FAX1 U394 ( .A(n1210), .B(n1048), .C(n871), .YC(n431), .YS(n432) );
  FAX1 U396 ( .A(n439), .B(n450), .C(n437), .YC(n434), .YS(n435) );
  FAX1 U397 ( .A(n454), .B(n441), .C(n452), .YC(n436), .YS(n437) );
  FAX1 U398 ( .A(n456), .B(n445), .C(n443), .YC(n438), .YS(n439) );
  FAX1 U399 ( .A(n460), .B(n447), .C(n458), .YC(n440), .YS(n441) );
  FAX1 U400 ( .A(n856), .B(n792), .C(n840), .YC(n442), .YS(n443) );
  FAX1 U401 ( .A(n824), .B(n808), .C(n776), .YC(n444), .YS(n445) );
  FAX1 U402 ( .A(n887), .B(n1051), .C(n872), .YC(n446), .YS(n447) );
  FAX1 U403 ( .A(n453), .B(n464), .C(n451), .YC(n448), .YS(n449) );
  FAX1 U404 ( .A(n468), .B(n455), .C(n466), .YC(n450), .YS(n451) );
  FAX1 U405 ( .A(n470), .B(n459), .C(n457), .YC(n452), .YS(n453) );
  FAX1 U406 ( .A(n793), .B(n461), .C(n472), .YC(n454), .YS(n455) );
  FAX1 U407 ( .A(n857), .B(n841), .C(n809), .YC(n456), .YS(n457) );
  FAX1 U408 ( .A(n825), .B(n777), .C(n474), .YC(n458), .YS(n459) );
  HAX1 U409 ( .A(n888), .B(n873), .YC(n460), .YS(n461) );
  FAX1 U410 ( .A(n467), .B(n478), .C(n465), .YC(n462), .YS(n463) );
  FAX1 U411 ( .A(n482), .B(n469), .C(n480), .YC(n464), .YS(n465) );
  FAX1 U412 ( .A(n484), .B(n471), .C(n473), .YC(n466), .YS(n467) );
  FAX1 U413 ( .A(n826), .B(n858), .C(n486), .YC(n468), .YS(n469) );
  FAX1 U414 ( .A(n874), .B(n794), .C(n475), .YC(n470), .YS(n471) );
  FAX1 U415 ( .A(n778), .B(n810), .C(n842), .YC(n472), .YS(n473) );
  HAX1 U416 ( .A(n889), .B(n743), .YC(n474), .YS(n475) );
  FAX1 U417 ( .A(n481), .B(n490), .C(n479), .YC(n476), .YS(n477) );
  FAX1 U418 ( .A(n485), .B(n483), .C(n492), .YC(n478), .YS(n479) );
  FAX1 U419 ( .A(n487), .B(n496), .C(n494), .YC(n480), .YS(n481) );
  FAX1 U420 ( .A(n859), .B(n795), .C(n843), .YC(n482), .YS(n483) );
  FAX1 U421 ( .A(n827), .B(n811), .C(n498), .YC(n484), .YS(n485) );
  HAX1 U422 ( .A(n890), .B(n875), .YC(n486), .YS(n487) );
  FAX1 U423 ( .A(n493), .B(n502), .C(n491), .YC(n488), .YS(n489) );
  FAX1 U424 ( .A(n497), .B(n495), .C(n504), .YC(n490), .YS(n491) );
  FAX1 U425 ( .A(n828), .B(n508), .C(n506), .YC(n492), .YS(n493) );
  FAX1 U426 ( .A(n876), .B(n860), .C(n499), .YC(n494), .YS(n495) );
  FAX1 U427 ( .A(n796), .B(n844), .C(n812), .YC(n496), .YS(n497) );
  HAX1 U428 ( .A(n891), .B(n744), .YC(n498), .YS(n499) );
  FAX1 U429 ( .A(n505), .B(n512), .C(n503), .YC(n500), .YS(n501) );
  FAX1 U430 ( .A(n516), .B(n514), .C(n507), .YC(n502), .YS(n503) );
  FAX1 U431 ( .A(n861), .B(n845), .C(n509), .YC(n504), .YS(n505) );
  FAX1 U432 ( .A(n829), .B(n813), .C(n518), .YC(n506), .YS(n507) );
  HAX1 U433 ( .A(n892), .B(n877), .YC(n508), .YS(n509) );
  FAX1 U434 ( .A(n515), .B(n522), .C(n513), .YC(n510), .YS(n511) );
  FAX1 U435 ( .A(n526), .B(n524), .C(n517), .YC(n512), .YS(n513) );
  FAX1 U436 ( .A(n878), .B(n830), .C(n519), .YC(n514), .YS(n515) );
  FAX1 U437 ( .A(n814), .B(n862), .C(n846), .YC(n516), .YS(n517) );
  HAX1 U438 ( .A(n893), .B(n745), .YC(n518), .YS(n519) );
  FAX1 U439 ( .A(n525), .B(n530), .C(n523), .YC(n520), .YS(n521) );
  FAX1 U440 ( .A(n863), .B(n527), .C(n532), .YC(n522), .YS(n523) );
  FAX1 U441 ( .A(n831), .B(n847), .C(n534), .YC(n524), .YS(n525) );
  HAX1 U442 ( .A(n894), .B(n879), .YC(n526), .YS(n527) );
  FAX1 U443 ( .A(n538), .B(n533), .C(n531), .YC(n528), .YS(n529) );
  FAX1 U444 ( .A(n880), .B(n535), .C(n540), .YC(n530), .YS(n531) );
  FAX1 U445 ( .A(n832), .B(n864), .C(n848), .YC(n532), .YS(n533) );
  HAX1 U446 ( .A(n895), .B(n746), .YC(n534), .YS(n535) );
  FAX1 U447 ( .A(n541), .B(n544), .C(n539), .YC(n536), .YS(n537) );
  FAX1 U448 ( .A(n865), .B(n849), .C(n546), .YC(n538), .YS(n539) );
  HAX1 U449 ( .A(n896), .B(n881), .YC(n540), .YS(n541) );
  FAX1 U450 ( .A(n547), .B(n550), .C(n545), .YC(n542), .YS(n543) );
  FAX1 U451 ( .A(n850), .B(n882), .C(n866), .YC(n544), .YS(n545) );
  HAX1 U452 ( .A(n897), .B(n747), .YC(n546), .YS(n547) );
  FAX1 U453 ( .A(n867), .B(n554), .C(n551), .YC(n548), .YS(n549) );
  HAX1 U454 ( .A(n898), .B(n883), .YC(n550), .YS(n551) );
  FAX1 U455 ( .A(n868), .B(n884), .C(n555), .YC(n552), .YS(n553) );
  HAX1 U456 ( .A(n899), .B(n748), .YC(n554), .YS(n555) );
  HAX1 U457 ( .A(n900), .B(n885), .YC(n556), .YS(n557) );
  HAX1 U458 ( .A(n901), .B(n749), .YC(n558), .YS(n559) );
  MUX2X1 U460 ( .B(n1206), .A(n1203), .S(n999), .Y(n560) );
  MUX2X1 U462 ( .B(n1203), .A(n1200), .S(n999), .Y(n561) );
  MUX2X1 U464 ( .B(n1200), .A(b[12]), .S(n999), .Y(n562) );
  MUX2X1 U466 ( .B(b[12]), .A(n1198), .S(n999), .Y(n563) );
  MUX2X1 U468 ( .B(n1198), .A(b[10]), .S(n999), .Y(n564) );
  MUX2X1 U470 ( .B(b[10]), .A(b[9]), .S(n999), .Y(n565) );
  MUX2X1 U472 ( .B(b[9]), .A(b[8]), .S(n1219), .Y(n566) );
  MUX2X1 U474 ( .B(b[8]), .A(b[7]), .S(n1219), .Y(n567) );
  MUX2X1 U476 ( .B(b[7]), .A(n1195), .S(n1219), .Y(n568) );
  MUX2X1 U478 ( .B(n1195), .A(b[5]), .S(n1219), .Y(n569) );
  MUX2X1 U480 ( .B(b[5]), .A(b[4]), .S(n1219), .Y(n570) );
  MUX2X1 U482 ( .B(b[4]), .A(b[3]), .S(n1219), .Y(n571) );
  MUX2X1 U484 ( .B(b[3]), .A(n1192), .S(n1219), .Y(n572) );
  MUX2X1 U486 ( .B(n1192), .A(n1190), .S(n1219), .Y(n573) );
  MUX2X1 U488 ( .B(n1190), .A(n1188), .S(n1219), .Y(n574) );
  MUX2X1 U495 ( .B(n1187), .A(n761), .S(n1016), .Y(n762) );
  MUX2X1 U497 ( .B(n1187), .A(n761), .S(n579), .Y(n763) );
  MUX2X1 U498 ( .B(n1206), .A(n1203), .S(n1185), .Y(n579) );
  MUX2X1 U499 ( .B(n1187), .A(n761), .S(n580), .Y(n764) );
  MUX2X1 U500 ( .B(n1203), .A(n1200), .S(n1185), .Y(n580) );
  MUX2X1 U501 ( .B(n1187), .A(n761), .S(n581), .Y(n765) );
  MUX2X1 U502 ( .B(n1200), .A(b[12]), .S(n1185), .Y(n581) );
  MUX2X1 U503 ( .B(n1187), .A(n761), .S(n582), .Y(n766) );
  MUX2X1 U504 ( .B(b[12]), .A(n1198), .S(n1185), .Y(n582) );
  MUX2X1 U505 ( .B(n1187), .A(n761), .S(n583), .Y(n767) );
  MUX2X1 U506 ( .B(n1198), .A(b[10]), .S(n1185), .Y(n583) );
  MUX2X1 U507 ( .B(n1187), .A(n761), .S(n584), .Y(n768) );
  MUX2X1 U508 ( .B(b[10]), .A(b[9]), .S(n1185), .Y(n584) );
  MUX2X1 U509 ( .B(n1187), .A(n761), .S(n585), .Y(n769) );
  MUX2X1 U510 ( .B(b[9]), .A(b[8]), .S(n1185), .Y(n585) );
  MUX2X1 U511 ( .B(n1186), .A(n761), .S(n586), .Y(n770) );
  MUX2X1 U512 ( .B(b[8]), .A(b[7]), .S(n1184), .Y(n586) );
  MUX2X1 U513 ( .B(n1186), .A(n761), .S(n587), .Y(n771) );
  MUX2X1 U514 ( .B(b[7]), .A(n1195), .S(n1184), .Y(n587) );
  MUX2X1 U515 ( .B(n1186), .A(n761), .S(n588), .Y(n772) );
  MUX2X1 U516 ( .B(n1195), .A(b[5]), .S(n1184), .Y(n588) );
  MUX2X1 U517 ( .B(n1186), .A(n761), .S(n589), .Y(n773) );
  MUX2X1 U518 ( .B(b[5]), .A(b[4]), .S(n1184), .Y(n589) );
  MUX2X1 U519 ( .B(n1186), .A(n761), .S(n590), .Y(n774) );
  MUX2X1 U520 ( .B(b[4]), .A(b[3]), .S(n1184), .Y(n590) );
  MUX2X1 U521 ( .B(n1186), .A(n761), .S(n591), .Y(n775) );
  MUX2X1 U522 ( .B(b[3]), .A(n1192), .S(n1184), .Y(n591) );
  MUX2X1 U523 ( .B(n1186), .A(n761), .S(n592), .Y(n776) );
  MUX2X1 U524 ( .B(n1192), .A(n1190), .S(n1184), .Y(n592) );
  MUX2X1 U525 ( .B(n1186), .A(n761), .S(n593), .Y(n777) );
  MUX2X1 U526 ( .B(n1190), .A(n1188), .S(n1184), .Y(n593) );
  MUX2X1 U527 ( .B(n1186), .A(n761), .S(n595), .Y(n778) );
  AND2X1 U530 ( .A(n1183), .B(n731), .Y(n744) );
  MUX2X1 U533 ( .B(n1183), .A(n779), .S(n1085), .Y(n780) );
  MUX2X1 U535 ( .B(n1183), .A(n779), .S(n598), .Y(n781) );
  MUX2X1 U536 ( .B(n1206), .A(n1203), .S(n1181), .Y(n598) );
  MUX2X1 U537 ( .B(n1183), .A(n779), .S(n599), .Y(n782) );
  MUX2X1 U538 ( .B(n1204), .A(n1200), .S(n1181), .Y(n599) );
  MUX2X1 U539 ( .B(n1183), .A(n779), .S(n600), .Y(n783) );
  MUX2X1 U540 ( .B(n1201), .A(b[12]), .S(n1181), .Y(n600) );
  MUX2X1 U541 ( .B(n1183), .A(n779), .S(n601), .Y(n784) );
  MUX2X1 U542 ( .B(b[12]), .A(n1198), .S(n1181), .Y(n601) );
  MUX2X1 U543 ( .B(n1183), .A(n779), .S(n602), .Y(n785) );
  MUX2X1 U544 ( .B(b[11]), .A(b[10]), .S(n1181), .Y(n602) );
  MUX2X1 U545 ( .B(n1183), .A(n779), .S(n603), .Y(n786) );
  MUX2X1 U546 ( .B(b[10]), .A(b[9]), .S(n1181), .Y(n603) );
  MUX2X1 U547 ( .B(n1183), .A(n779), .S(n604), .Y(n787) );
  MUX2X1 U548 ( .B(b[9]), .A(b[8]), .S(n1181), .Y(n604) );
  MUX2X1 U549 ( .B(n1182), .A(n779), .S(n605), .Y(n788) );
  MUX2X1 U550 ( .B(b[8]), .A(b[7]), .S(n1180), .Y(n605) );
  MUX2X1 U551 ( .B(n1182), .A(n779), .S(n606), .Y(n789) );
  MUX2X1 U552 ( .B(b[7]), .A(n1195), .S(n1180), .Y(n606) );
  MUX2X1 U553 ( .B(n1182), .A(n779), .S(n607), .Y(n790) );
  MUX2X1 U554 ( .B(n1196), .A(b[5]), .S(n1180), .Y(n607) );
  MUX2X1 U555 ( .B(n1182), .A(n779), .S(n608), .Y(n791) );
  MUX2X1 U556 ( .B(b[5]), .A(b[4]), .S(n1180), .Y(n608) );
  MUX2X1 U557 ( .B(n1182), .A(n779), .S(n609), .Y(n792) );
  MUX2X1 U558 ( .B(b[4]), .A(b[3]), .S(n1180), .Y(n609) );
  MUX2X1 U559 ( .B(n1182), .A(n779), .S(n610), .Y(n793) );
  MUX2X1 U560 ( .B(b[3]), .A(n1192), .S(n1180), .Y(n610) );
  MUX2X1 U561 ( .B(n1182), .A(n779), .S(n611), .Y(n794) );
  MUX2X1 U562 ( .B(n1193), .A(n1190), .S(n1180), .Y(n611) );
  MUX2X1 U563 ( .B(n1182), .A(n779), .S(n612), .Y(n795) );
  MUX2X1 U564 ( .B(b[1]), .A(n1188), .S(n1180), .Y(n612) );
  MUX2X1 U565 ( .B(n1182), .A(n779), .S(n614), .Y(n796) );
  OR2X1 U566 ( .A(n1181), .B(n1189), .Y(n614) );
  AND2X1 U568 ( .A(n1179), .B(n733), .Y(n745) );
  MUX2X1 U571 ( .B(n1179), .A(n797), .S(n1106), .Y(n798) );
  MUX2X1 U573 ( .B(n1179), .A(n797), .S(n617), .Y(n799) );
  MUX2X1 U574 ( .B(n1206), .A(n1203), .S(n1177), .Y(n617) );
  MUX2X1 U575 ( .B(n1179), .A(n797), .S(n618), .Y(n800) );
  MUX2X1 U576 ( .B(n1204), .A(n1200), .S(n1177), .Y(n618) );
  MUX2X1 U577 ( .B(n1179), .A(n797), .S(n619), .Y(n801) );
  MUX2X1 U578 ( .B(n1201), .A(b[12]), .S(n1177), .Y(n619) );
  MUX2X1 U579 ( .B(n1179), .A(n797), .S(n620), .Y(n802) );
  MUX2X1 U580 ( .B(b[12]), .A(n1198), .S(n1177), .Y(n620) );
  MUX2X1 U581 ( .B(n1179), .A(n797), .S(n621), .Y(n803) );
  MUX2X1 U582 ( .B(b[11]), .A(b[10]), .S(n1177), .Y(n621) );
  MUX2X1 U583 ( .B(n1179), .A(n797), .S(n622), .Y(n804) );
  MUX2X1 U584 ( .B(b[10]), .A(b[9]), .S(n1177), .Y(n622) );
  MUX2X1 U585 ( .B(n1179), .A(n797), .S(n623), .Y(n805) );
  MUX2X1 U586 ( .B(b[9]), .A(b[8]), .S(n1177), .Y(n623) );
  MUX2X1 U587 ( .B(n1178), .A(n797), .S(n624), .Y(n806) );
  MUX2X1 U588 ( .B(b[8]), .A(b[7]), .S(n1176), .Y(n624) );
  MUX2X1 U589 ( .B(n1178), .A(n797), .S(n625), .Y(n807) );
  MUX2X1 U590 ( .B(b[7]), .A(n1195), .S(n1176), .Y(n625) );
  MUX2X1 U591 ( .B(n1178), .A(n797), .S(n626), .Y(n808) );
  MUX2X1 U592 ( .B(n1196), .A(b[5]), .S(n1176), .Y(n626) );
  MUX2X1 U593 ( .B(n1178), .A(n797), .S(n627), .Y(n809) );
  MUX2X1 U594 ( .B(b[5]), .A(b[4]), .S(n1176), .Y(n627) );
  MUX2X1 U595 ( .B(n1178), .A(n797), .S(n628), .Y(n810) );
  MUX2X1 U596 ( .B(b[4]), .A(b[3]), .S(n1176), .Y(n628) );
  MUX2X1 U597 ( .B(n1178), .A(n797), .S(n629), .Y(n811) );
  MUX2X1 U598 ( .B(b[3]), .A(n1192), .S(n1176), .Y(n629) );
  MUX2X1 U599 ( .B(n1178), .A(n797), .S(n630), .Y(n812) );
  MUX2X1 U600 ( .B(n1193), .A(n1190), .S(n1176), .Y(n630) );
  MUX2X1 U601 ( .B(n1178), .A(n797), .S(n631), .Y(n813) );
  MUX2X1 U602 ( .B(b[1]), .A(n1188), .S(n1176), .Y(n631) );
  MUX2X1 U603 ( .B(n1178), .A(n797), .S(n633), .Y(n814) );
  OR2X1 U604 ( .A(n1177), .B(n1189), .Y(n633) );
  AND2X1 U606 ( .A(n1175), .B(n735), .Y(n746) );
  MUX2X1 U609 ( .B(n1175), .A(n815), .S(n1059), .Y(n816) );
  MUX2X1 U611 ( .B(n1175), .A(n815), .S(n636), .Y(n817) );
  MUX2X1 U612 ( .B(n1206), .A(n1203), .S(n1173), .Y(n636) );
  MUX2X1 U613 ( .B(n1175), .A(n815), .S(n637), .Y(n818) );
  MUX2X1 U614 ( .B(n1203), .A(n1200), .S(n1173), .Y(n637) );
  MUX2X1 U615 ( .B(n1175), .A(n815), .S(n638), .Y(n819) );
  MUX2X1 U616 ( .B(n1200), .A(b[12]), .S(n1173), .Y(n638) );
  MUX2X1 U617 ( .B(n1175), .A(n815), .S(n639), .Y(n820) );
  MUX2X1 U618 ( .B(b[12]), .A(n1198), .S(n1173), .Y(n639) );
  MUX2X1 U619 ( .B(n1175), .A(n815), .S(n640), .Y(n821) );
  MUX2X1 U620 ( .B(n1198), .A(b[10]), .S(n1173), .Y(n640) );
  MUX2X1 U621 ( .B(n1175), .A(n815), .S(n641), .Y(n822) );
  MUX2X1 U622 ( .B(b[10]), .A(b[9]), .S(n1173), .Y(n641) );
  MUX2X1 U623 ( .B(n1175), .A(n815), .S(n642), .Y(n823) );
  MUX2X1 U624 ( .B(b[9]), .A(b[8]), .S(n1173), .Y(n642) );
  MUX2X1 U625 ( .B(n1174), .A(n815), .S(n643), .Y(n824) );
  MUX2X1 U626 ( .B(b[8]), .A(b[7]), .S(n1172), .Y(n643) );
  MUX2X1 U627 ( .B(n1174), .A(n815), .S(n644), .Y(n825) );
  MUX2X1 U628 ( .B(b[7]), .A(n1195), .S(n1172), .Y(n644) );
  MUX2X1 U629 ( .B(n1174), .A(n815), .S(n645), .Y(n826) );
  MUX2X1 U630 ( .B(n1195), .A(b[5]), .S(n1172), .Y(n645) );
  MUX2X1 U631 ( .B(n1174), .A(n815), .S(n646), .Y(n827) );
  MUX2X1 U632 ( .B(b[5]), .A(b[4]), .S(n1172), .Y(n646) );
  MUX2X1 U633 ( .B(n1174), .A(n815), .S(n647), .Y(n828) );
  MUX2X1 U634 ( .B(b[4]), .A(b[3]), .S(n1172), .Y(n647) );
  MUX2X1 U635 ( .B(n1174), .A(n815), .S(n648), .Y(n829) );
  MUX2X1 U636 ( .B(b[3]), .A(n1192), .S(n1172), .Y(n648) );
  MUX2X1 U637 ( .B(n1174), .A(n815), .S(n649), .Y(n830) );
  MUX2X1 U638 ( .B(n1192), .A(n1190), .S(n1172), .Y(n649) );
  MUX2X1 U639 ( .B(n1174), .A(n815), .S(n650), .Y(n831) );
  MUX2X1 U640 ( .B(n1190), .A(n1188), .S(n1172), .Y(n650) );
  MUX2X1 U641 ( .B(n1174), .A(n815), .S(n652), .Y(n832) );
  MUX2X1 U647 ( .B(n1171), .A(n833), .S(n1125), .Y(n834) );
  MUX2X1 U649 ( .B(n1171), .A(n833), .S(n655), .Y(n835) );
  MUX2X1 U650 ( .B(n1206), .A(n1203), .S(n1169), .Y(n655) );
  MUX2X1 U651 ( .B(n1171), .A(n833), .S(n656), .Y(n836) );
  MUX2X1 U652 ( .B(n1203), .A(n1200), .S(n1169), .Y(n656) );
  MUX2X1 U653 ( .B(n1171), .A(n833), .S(n657), .Y(n837) );
  MUX2X1 U654 ( .B(n1200), .A(b[12]), .S(n1169), .Y(n657) );
  MUX2X1 U655 ( .B(n1171), .A(n833), .S(n658), .Y(n838) );
  MUX2X1 U656 ( .B(b[12]), .A(n1198), .S(n1169), .Y(n658) );
  MUX2X1 U657 ( .B(n1171), .A(n833), .S(n659), .Y(n839) );
  MUX2X1 U658 ( .B(n1198), .A(b[10]), .S(n1169), .Y(n659) );
  MUX2X1 U659 ( .B(n1171), .A(n833), .S(n660), .Y(n840) );
  MUX2X1 U660 ( .B(b[10]), .A(b[9]), .S(n1169), .Y(n660) );
  MUX2X1 U661 ( .B(n1171), .A(n833), .S(n661), .Y(n841) );
  MUX2X1 U662 ( .B(b[9]), .A(b[8]), .S(n1169), .Y(n661) );
  MUX2X1 U663 ( .B(n1170), .A(n833), .S(n662), .Y(n842) );
  MUX2X1 U664 ( .B(b[8]), .A(b[7]), .S(n1168), .Y(n662) );
  MUX2X1 U665 ( .B(n1170), .A(n833), .S(n663), .Y(n843) );
  MUX2X1 U666 ( .B(b[7]), .A(n1195), .S(n1168), .Y(n663) );
  MUX2X1 U667 ( .B(n1170), .A(n833), .S(n664), .Y(n844) );
  MUX2X1 U668 ( .B(n1195), .A(b[5]), .S(n1168), .Y(n664) );
  MUX2X1 U669 ( .B(n1170), .A(n833), .S(n665), .Y(n845) );
  MUX2X1 U670 ( .B(b[5]), .A(b[4]), .S(n1168), .Y(n665) );
  MUX2X1 U671 ( .B(n1170), .A(n833), .S(n666), .Y(n846) );
  MUX2X1 U672 ( .B(b[4]), .A(b[3]), .S(n1168), .Y(n666) );
  MUX2X1 U673 ( .B(n1170), .A(n833), .S(n667), .Y(n847) );
  MUX2X1 U674 ( .B(b[3]), .A(n1192), .S(n1168), .Y(n667) );
  MUX2X1 U675 ( .B(n1170), .A(n833), .S(n668), .Y(n848) );
  MUX2X1 U676 ( .B(n1192), .A(n1190), .S(n1168), .Y(n668) );
  MUX2X1 U677 ( .B(n1170), .A(n833), .S(n669), .Y(n849) );
  MUX2X1 U678 ( .B(n1190), .A(n1188), .S(n1168), .Y(n669) );
  MUX2X1 U679 ( .B(n1170), .A(n833), .S(n671), .Y(n850) );
  OR2X1 U680 ( .A(n1169), .B(n1189), .Y(n671) );
  AND2X1 U682 ( .A(n1167), .B(n739), .Y(n748) );
  MUX2X1 U685 ( .B(n1167), .A(n851), .S(n1107), .Y(n852) );
  MUX2X1 U687 ( .B(n1167), .A(n851), .S(n674), .Y(n853) );
  MUX2X1 U688 ( .B(n1206), .A(n1203), .S(n1165), .Y(n674) );
  MUX2X1 U689 ( .B(n1167), .A(n851), .S(n675), .Y(n854) );
  MUX2X1 U690 ( .B(n1204), .A(n1200), .S(n1165), .Y(n675) );
  MUX2X1 U691 ( .B(n1167), .A(n851), .S(n676), .Y(n855) );
  MUX2X1 U692 ( .B(n1201), .A(b[12]), .S(n1165), .Y(n676) );
  MUX2X1 U693 ( .B(n1167), .A(n851), .S(n677), .Y(n856) );
  MUX2X1 U694 ( .B(b[12]), .A(n1198), .S(n1165), .Y(n677) );
  MUX2X1 U695 ( .B(n1167), .A(n851), .S(n678), .Y(n857) );
  MUX2X1 U696 ( .B(n1198), .A(b[10]), .S(n1165), .Y(n678) );
  MUX2X1 U697 ( .B(n1167), .A(n851), .S(n679), .Y(n858) );
  MUX2X1 U698 ( .B(b[10]), .A(b[9]), .S(n1165), .Y(n679) );
  MUX2X1 U699 ( .B(n1167), .A(n851), .S(n680), .Y(n859) );
  MUX2X1 U700 ( .B(b[9]), .A(b[8]), .S(n1165), .Y(n680) );
  MUX2X1 U701 ( .B(n1166), .A(n851), .S(n681), .Y(n860) );
  MUX2X1 U702 ( .B(b[8]), .A(b[7]), .S(n1164), .Y(n681) );
  MUX2X1 U703 ( .B(n1166), .A(n851), .S(n682), .Y(n861) );
  MUX2X1 U704 ( .B(b[7]), .A(n1195), .S(n1164), .Y(n682) );
  MUX2X1 U705 ( .B(n1166), .A(n851), .S(n683), .Y(n862) );
  MUX2X1 U706 ( .B(n1196), .A(b[5]), .S(n1164), .Y(n683) );
  MUX2X1 U707 ( .B(n1166), .A(n851), .S(n684), .Y(n863) );
  MUX2X1 U708 ( .B(b[5]), .A(b[4]), .S(n1164), .Y(n684) );
  MUX2X1 U709 ( .B(n1166), .A(n851), .S(n685), .Y(n864) );
  MUX2X1 U710 ( .B(b[4]), .A(b[3]), .S(n1164), .Y(n685) );
  MUX2X1 U711 ( .B(n1166), .A(n851), .S(n686), .Y(n865) );
  MUX2X1 U712 ( .B(b[3]), .A(n1192), .S(n1164), .Y(n686) );
  MUX2X1 U713 ( .B(n1166), .A(n851), .S(n687), .Y(n866) );
  MUX2X1 U714 ( .B(n1193), .A(n1190), .S(n1164), .Y(n687) );
  MUX2X1 U715 ( .B(n1166), .A(n851), .S(n688), .Y(n867) );
  MUX2X1 U716 ( .B(b[1]), .A(n1188), .S(n1164), .Y(n688) );
  MUX2X1 U717 ( .B(n1166), .A(n851), .S(n690), .Y(n868) );
  OR2X1 U718 ( .A(n1165), .B(n1189), .Y(n690) );
  AND2X1 U720 ( .A(n1163), .B(n741), .Y(n749) );
  MUX2X1 U723 ( .B(n1163), .A(n1143), .S(n1086), .Y(n870) );
  MUX2X1 U725 ( .B(n1163), .A(n1143), .S(n693), .Y(n871) );
  MUX2X1 U726 ( .B(n1206), .A(n1203), .S(n1161), .Y(n693) );
  MUX2X1 U727 ( .B(n1163), .A(n1143), .S(n694), .Y(n872) );
  MUX2X1 U728 ( .B(n1204), .A(n1200), .S(n1161), .Y(n694) );
  MUX2X1 U729 ( .B(n1163), .A(n1143), .S(n695), .Y(n873) );
  MUX2X1 U730 ( .B(n1201), .A(b[12]), .S(n1161), .Y(n695) );
  MUX2X1 U731 ( .B(n1163), .A(n1143), .S(n696), .Y(n874) );
  MUX2X1 U732 ( .B(b[12]), .A(n1198), .S(n1161), .Y(n696) );
  MUX2X1 U733 ( .B(n1163), .A(n1143), .S(n697), .Y(n875) );
  MUX2X1 U734 ( .B(b[11]), .A(b[10]), .S(n1161), .Y(n697) );
  MUX2X1 U735 ( .B(n1163), .A(n1143), .S(n698), .Y(n876) );
  MUX2X1 U736 ( .B(b[10]), .A(b[9]), .S(n1161), .Y(n698) );
  MUX2X1 U737 ( .B(n1163), .A(n1143), .S(n699), .Y(n877) );
  MUX2X1 U738 ( .B(b[9]), .A(b[8]), .S(n1161), .Y(n699) );
  MUX2X1 U739 ( .B(n1162), .A(n1143), .S(n700), .Y(n878) );
  MUX2X1 U740 ( .B(b[8]), .A(b[7]), .S(n1160), .Y(n700) );
  MUX2X1 U741 ( .B(n1162), .A(n1143), .S(n701), .Y(n879) );
  MUX2X1 U742 ( .B(b[7]), .A(n1195), .S(n1160), .Y(n701) );
  MUX2X1 U743 ( .B(n1162), .A(n1143), .S(n702), .Y(n880) );
  MUX2X1 U744 ( .B(n1196), .A(b[5]), .S(n1160), .Y(n702) );
  MUX2X1 U745 ( .B(n1162), .A(n1143), .S(n703), .Y(n881) );
  MUX2X1 U746 ( .B(b[5]), .A(b[4]), .S(n1160), .Y(n703) );
  MUX2X1 U747 ( .B(n1162), .A(n1143), .S(n704), .Y(n882) );
  MUX2X1 U748 ( .B(b[4]), .A(b[3]), .S(n1160), .Y(n704) );
  MUX2X1 U749 ( .B(n1162), .A(n1143), .S(n705), .Y(n883) );
  MUX2X1 U750 ( .B(b[3]), .A(n1192), .S(n1160), .Y(n705) );
  MUX2X1 U751 ( .B(n1162), .A(n1143), .S(n706), .Y(n884) );
  MUX2X1 U752 ( .B(n1193), .A(n1190), .S(n1160), .Y(n706) );
  MUX2X1 U753 ( .B(n1162), .A(n1143), .S(n707), .Y(n885) );
  MUX2X1 U754 ( .B(n1190), .A(n1188), .S(n1160), .Y(n707) );
  MUX2X1 U755 ( .B(n1162), .A(n1143), .S(n709), .Y(n886) );
  OR2X1 U756 ( .A(n1161), .B(n1189), .Y(n709) );
  AND2X1 U758 ( .A(n1158), .B(a[1]), .Y(n750) );
  MUX2X1 U761 ( .B(n1159), .A(n1211), .S(n1124), .Y(n887) );
  MUX2X1 U763 ( .B(n1159), .A(n1211), .S(n712), .Y(n888) );
  MUX2X1 U764 ( .B(n1206), .A(n1203), .S(n1208), .Y(n712) );
  MUX2X1 U765 ( .B(n1159), .A(n1211), .S(n713), .Y(n889) );
  MUX2X1 U766 ( .B(n1204), .A(n1200), .S(n1208), .Y(n713) );
  MUX2X1 U767 ( .B(n1159), .A(n1211), .S(n714), .Y(n890) );
  MUX2X1 U768 ( .B(n1201), .A(b[12]), .S(n1208), .Y(n714) );
  MUX2X1 U769 ( .B(n1159), .A(n1211), .S(n715), .Y(n891) );
  MUX2X1 U770 ( .B(b[12]), .A(n1198), .S(n1208), .Y(n715) );
  MUX2X1 U771 ( .B(n1159), .A(n1211), .S(n716), .Y(n892) );
  MUX2X1 U772 ( .B(n1198), .A(b[10]), .S(n1208), .Y(n716) );
  MUX2X1 U773 ( .B(n1159), .A(n1211), .S(n717), .Y(n893) );
  MUX2X1 U774 ( .B(b[10]), .A(b[9]), .S(n1208), .Y(n717) );
  MUX2X1 U775 ( .B(n1159), .A(n1211), .S(n718), .Y(n894) );
  MUX2X1 U776 ( .B(b[9]), .A(b[8]), .S(n1208), .Y(n718) );
  MUX2X1 U777 ( .B(n1159), .A(n1211), .S(n719), .Y(n895) );
  MUX2X1 U778 ( .B(b[8]), .A(b[7]), .S(n1208), .Y(n719) );
  MUX2X1 U779 ( .B(n1159), .A(n1211), .S(n720), .Y(n896) );
  MUX2X1 U780 ( .B(b[7]), .A(n1195), .S(n1208), .Y(n720) );
  MUX2X1 U781 ( .B(n1159), .A(n1211), .S(n721), .Y(n897) );
  MUX2X1 U782 ( .B(n1196), .A(b[5]), .S(n1209), .Y(n721) );
  MUX2X1 U783 ( .B(n1159), .A(n1211), .S(n722), .Y(n898) );
  MUX2X1 U784 ( .B(b[5]), .A(b[4]), .S(n1209), .Y(n722) );
  MUX2X1 U785 ( .B(n1159), .A(n1211), .S(n723), .Y(n899) );
  MUX2X1 U786 ( .B(b[4]), .A(b[3]), .S(n1209), .Y(n723) );
  MUX2X1 U787 ( .B(n1159), .A(n1211), .S(n724), .Y(n900) );
  MUX2X1 U788 ( .B(b[3]), .A(n1192), .S(n1208), .Y(n724) );
  MUX2X1 U789 ( .B(n1158), .A(n1211), .S(n725), .Y(n901) );
  MUX2X1 U790 ( .B(n1193), .A(n1190), .S(n1208), .Y(n725) );
  MUX2X1 U791 ( .B(n1158), .A(n1211), .S(n726), .Y(n902) );
  MUX2X1 U792 ( .B(n1190), .A(n1188), .S(n1208), .Y(n726) );
  MUX2X1 U793 ( .B(n1158), .A(n1211), .S(n728), .Y(n903) );
  OR2X1 U794 ( .A(n1209), .B(n1189), .Y(n728) );
  OAI21X1 U798 ( .A(a[13]), .B(a[14]), .C(n1219), .Y(n44) );
  XNOR2X1 U801 ( .A(a[14]), .B(a[13]), .Y(n48) );
  OAI21X1 U803 ( .A(a[12]), .B(a[11]), .C(n1218), .Y(n38) );
  XNOR2X1 U806 ( .A(a[11]), .B(a[12]), .Y(n42) );
  OAI21X1 U808 ( .A(a[10]), .B(n1215), .C(n1217), .Y(n32) );
  XNOR2X1 U811 ( .A(n1215), .B(a[10]), .Y(n36) );
  OAI21X1 U813 ( .A(a[8]), .B(a[7]), .C(n1216), .Y(n26) );
  XNOR2X1 U816 ( .A(a[7]), .B(a[8]), .Y(n30) );
  OAI21X1 U818 ( .A(a[5]), .B(a[6]), .C(n1214), .Y(n20) );
  XNOR2X1 U821 ( .A(a[6]), .B(a[5]), .Y(n24) );
  OAI21X1 U823 ( .A(a[4]), .B(a[3]), .C(n1213), .Y(n14) );
  XNOR2X1 U826 ( .A(a[3]), .B(a[4]), .Y(n18) );
  OAI21X1 U828 ( .A(a[2]), .B(n1210), .C(n1212), .Y(n8) );
  XNOR2X1 U831 ( .A(n1210), .B(a[2]), .Y(n12) );
  INVX2 U838 ( .A(n1207), .Y(n1206) );
  BUFX2 U839 ( .A(a[15]), .Y(n998) );
  INVX1 U840 ( .A(a[15]), .Y(n999) );
  AND2X2 U841 ( .A(b[15]), .B(n1169), .Y(n654) );
  AND2X2 U842 ( .A(b[15]), .B(n1165), .Y(n673) );
  AND2X2 U843 ( .A(b[15]), .B(n1181), .Y(n597) );
  AND2X2 U844 ( .A(b[15]), .B(n1185), .Y(n578) );
  INVX2 U845 ( .A(b[0]), .Y(n1189) );
  INVX1 U846 ( .A(b[1]), .Y(n1191) );
  INVX2 U847 ( .A(n733), .Y(n797) );
  AND2X1 U848 ( .A(n1206), .B(n1173), .Y(n635) );
  OR2X1 U849 ( .A(n576), .B(n1219), .Y(n760) );
  OR2X1 U850 ( .A(n1219), .B(n1189), .Y(n576) );
  AND2X1 U851 ( .A(n1206), .B(n1161), .Y(n692) );
  AND2X1 U852 ( .A(n1187), .B(n729), .Y(n743) );
  OR2X1 U853 ( .A(n1185), .B(n1189), .Y(n595) );
  OR2X1 U854 ( .A(n568), .B(n1219), .Y(n755) );
  OR2X1 U855 ( .A(n570), .B(n1219), .Y(n756) );
  BUFX2 U856 ( .A(n48), .Y(n1184) );
  INVX1 U857 ( .A(n757), .Y(n1047) );
  OR2X1 U858 ( .A(n574), .B(n1219), .Y(n759) );
  BUFX2 U859 ( .A(n42), .Y(n1180) );
  OR2X1 U860 ( .A(n1173), .B(n1189), .Y(n652) );
  OR2X1 U861 ( .A(n566), .B(n999), .Y(n754) );
  OR2X1 U862 ( .A(n1103), .B(n1120), .Y(n180) );
  INVX1 U863 ( .A(n190), .Y(n1104) );
  OR2X1 U864 ( .A(n1076), .B(n1136), .Y(n157) );
  OR2X1 U865 ( .A(n364), .B(n375), .Y(n159) );
  AND2X1 U866 ( .A(n434), .B(n420), .Y(n183) );
  AND2X1 U867 ( .A(a[5]), .B(n1212), .Y(n1221) );
  OR2X1 U868 ( .A(n564), .B(n999), .Y(n753) );
  AND2X1 U869 ( .A(n1145), .B(n1144), .Y(n143) );
  AND2X1 U870 ( .A(n1065), .B(n171), .Y(n96) );
  AND2X1 U871 ( .A(n1146), .B(n1148), .Y(n226) );
  OR2X1 U872 ( .A(n529), .B(n536), .Y(n1148) );
  AND2X1 U873 ( .A(n1171), .B(n737), .Y(n747) );
  INVX1 U874 ( .A(n1189), .Y(n1188) );
  INVX2 U875 ( .A(n1191), .Y(n1190) );
  BUFX2 U876 ( .A(n12), .Y(n1160) );
  AND2X1 U877 ( .A(n1093), .B(n1150), .Y(n88) );
  OR2X1 U878 ( .A(n553), .B(n556), .Y(n1156) );
  AND2X1 U879 ( .A(n1063), .B(n1154), .Y(n113) );
  AND2X1 U880 ( .A(n750), .B(n903), .Y(n262) );
  OR2X1 U881 ( .A(n562), .B(n999), .Y(n752) );
  BUFX2 U882 ( .A(n48), .Y(n1185) );
  OR2X1 U883 ( .A(n560), .B(n999), .Y(n751) );
  INVX1 U884 ( .A(a[11]), .Y(n1217) );
  INVX1 U885 ( .A(b[15]), .Y(n1207) );
  OR2X1 U886 ( .A(n561), .B(n999), .Y(n297) );
  INVX1 U887 ( .A(a[7]), .Y(n1214) );
  AND2X1 U888 ( .A(n886), .B(n559), .Y(n258) );
  INVX2 U889 ( .A(n739), .Y(n851) );
  INVX2 U890 ( .A(n731), .Y(n779) );
  OR2X1 U891 ( .A(n903), .B(n750), .Y(n261) );
  INVX2 U892 ( .A(n729), .Y(n761) );
  INVX1 U893 ( .A(a[5]), .Y(n1213) );
  INVX2 U894 ( .A(n737), .Y(n833) );
  OR2X2 U895 ( .A(n1104), .B(n1111), .Y(n188) );
  OR2X2 U896 ( .A(n559), .B(n886), .Y(n1154) );
  AND2X2 U897 ( .A(a[3]), .B(n1211), .Y(n1220) );
  OR2X2 U898 ( .A(n1141), .B(n260), .Y(n259) );
  INVX2 U899 ( .A(n1199), .Y(n1198) );
  INVX2 U900 ( .A(n1202), .Y(n1200) );
  INVX2 U901 ( .A(a[0]), .Y(n1208) );
  AND2X2 U902 ( .A(a[0]), .B(n1211), .Y(n2) );
  INVX8 U903 ( .A(a[15]), .Y(n1219) );
  INVX4 U904 ( .A(n1142), .Y(n1210) );
  INVX8 U905 ( .A(n1210), .Y(n1211) );
  INVX1 U906 ( .A(n226), .Y(n1000) );
  AND2X2 U907 ( .A(n1067), .B(n1079), .Y(n178) );
  INVX1 U908 ( .A(n178), .Y(n1001) );
  INVX1 U909 ( .A(n157), .Y(n1002) );
  AND2X2 U910 ( .A(n1002), .B(n1029), .Y(n155) );
  INVX1 U911 ( .A(n155), .Y(n1003) );
  OR2X2 U912 ( .A(n1003), .B(n1032), .Y(n141) );
  INVX1 U913 ( .A(n141), .Y(n1004) );
  BUFX2 U914 ( .A(n220), .Y(n1005) );
  BUFX2 U915 ( .A(n132), .Y(n1006) );
  BUFX2 U916 ( .A(n238), .Y(n1007) );
  BUFX2 U917 ( .A(n198), .Y(n1008) );
  BUFX2 U918 ( .A(n227), .Y(n1009) );
  BUFX2 U919 ( .A(n209), .Y(n1010) );
  INVX1 U920 ( .A(n179), .Y(n1011) );
  INVX1 U921 ( .A(n1011), .Y(n1012) );
  BUFX2 U922 ( .A(n144), .Y(n1013) );
  OR2X1 U923 ( .A(n1102), .B(n1119), .Y(n199) );
  INVX1 U924 ( .A(n199), .Y(n1014) );
  AND2X1 U925 ( .A(n1147), .B(n1149), .Y(n208) );
  INVX1 U926 ( .A(n208), .Y(n1015) );
  INVX1 U927 ( .A(n578), .Y(n1016) );
  BUFX2 U928 ( .A(n232), .Y(n1017) );
  BUFX2 U929 ( .A(n214), .Y(n1018) );
  BUFX2 U930 ( .A(n149), .Y(n1019) );
  AND2X1 U931 ( .A(n1129), .B(n1146), .Y(n108) );
  INVX1 U932 ( .A(n108), .Y(n1020) );
  AND2X1 U933 ( .A(n1101), .B(n164), .Y(n95) );
  INVX1 U934 ( .A(n95), .Y(n1021) );
  AND2X1 U935 ( .A(n1098), .B(n1144), .Y(n93) );
  INVX1 U936 ( .A(n93), .Y(n1022) );
  AND2X1 U937 ( .A(n1095), .B(n1151), .Y(n90) );
  INVX1 U938 ( .A(n90), .Y(n1023) );
  AND2X1 U939 ( .A(n1109), .B(n1148), .Y(n107) );
  INVX1 U940 ( .A(n107), .Y(n1024) );
  AND2X1 U941 ( .A(n1094), .B(n1149), .Y(n104) );
  INVX1 U942 ( .A(n104), .Y(n1025) );
  AND2X1 U943 ( .A(n1075), .B(n1145), .Y(n92) );
  INVX1 U944 ( .A(n92), .Y(n1026) );
  AND2X1 U945 ( .A(n1116), .B(n138), .Y(n91) );
  INVX1 U946 ( .A(n91), .Y(n1027) );
  AND2X1 U947 ( .A(n1113), .B(n122), .Y(n87) );
  INVX1 U948 ( .A(n87), .Y(n1028) );
  OR2X1 U949 ( .A(n1081), .B(n1121), .Y(n169) );
  INVX1 U950 ( .A(n169), .Y(n1029) );
  INVX1 U951 ( .A(n156), .Y(n1030) );
  INVX1 U952 ( .A(n1030), .Y(n1031) );
  INVX1 U953 ( .A(n143), .Y(n1032) );
  INVX1 U954 ( .A(n140), .Y(n1033) );
  INVX1 U955 ( .A(n1033), .Y(n1034) );
  INVX1 U956 ( .A(n1033), .Y(n1035) );
  BUFX2 U957 ( .A(n1006), .Y(n1036) );
  INVX1 U958 ( .A(n124), .Y(n1037) );
  INVX1 U959 ( .A(n1037), .Y(n1038) );
  INVX1 U960 ( .A(n1037), .Y(n1039) );
  AND2X1 U961 ( .A(n998), .B(n1218), .Y(n1226) );
  INVX1 U962 ( .A(n1226), .Y(n1040) );
  INVX1 U963 ( .A(n751), .Y(n1041) );
  INVX1 U964 ( .A(n752), .Y(n1042) );
  INVX1 U965 ( .A(n754), .Y(n1043) );
  INVX1 U966 ( .A(n753), .Y(n1044) );
  INVX1 U967 ( .A(n755), .Y(n1045) );
  INVX1 U968 ( .A(n756), .Y(n1046) );
  OR2X1 U969 ( .A(n572), .B(n1219), .Y(n757) );
  INVX1 U970 ( .A(n759), .Y(n1048) );
  INVX1 U971 ( .A(n1221), .Y(n1049) );
  AND2X1 U972 ( .A(n1057), .B(n182), .Y(n98) );
  INVX1 U973 ( .A(n98), .Y(n1050) );
  INVX1 U974 ( .A(n760), .Y(n1051) );
  AND2X1 U975 ( .A(a[13]), .B(n1217), .Y(n1225) );
  INVX1 U976 ( .A(n1225), .Y(n1052) );
  AND2X1 U977 ( .A(n1064), .B(n1156), .Y(n111) );
  INVX1 U978 ( .A(n111), .Y(n1053) );
  AND2X1 U979 ( .A(n1077), .B(n252), .Y(n112) );
  INVX1 U980 ( .A(n112), .Y(n1054) );
  AND2X1 U981 ( .A(n1066), .B(n278), .Y(n100) );
  INVX1 U982 ( .A(n100), .Y(n1055) );
  BUFX2 U983 ( .A(n192), .Y(n1056) );
  INVX1 U984 ( .A(n183), .Y(n1057) );
  INVX1 U985 ( .A(n297), .Y(n1058) );
  INVX1 U986 ( .A(n635), .Y(n1059) );
  AND2X1 U987 ( .A(n1078), .B(n201), .Y(n102) );
  INVX1 U988 ( .A(n102), .Y(n1060) );
  AND2X1 U989 ( .A(n1115), .B(n159), .Y(n94) );
  INVX1 U990 ( .A(n94), .Y(n1061) );
  BUFX2 U991 ( .A(n161), .Y(n1062) );
  INVX1 U992 ( .A(n258), .Y(n1063) );
  AND2X1 U993 ( .A(n556), .B(n553), .Y(n250) );
  INVX1 U994 ( .A(n250), .Y(n1064) );
  AND2X1 U995 ( .A(n403), .B(n390), .Y(n172) );
  INVX1 U996 ( .A(n172), .Y(n1065) );
  AND2X1 U997 ( .A(n462), .B(n449), .Y(n191) );
  INVX1 U998 ( .A(n191), .Y(n1066) );
  INVX1 U999 ( .A(n188), .Y(n1067) );
  OR2X1 U1000 ( .A(n563), .B(n999), .Y(n307) );
  INVX1 U1001 ( .A(n307), .Y(n1068) );
  AND2X1 U1002 ( .A(a[11]), .B(n1216), .Y(n1224) );
  INVX1 U1003 ( .A(n1224), .Y(n1069) );
  AND2X1 U1004 ( .A(n1097), .B(n1155), .Y(n109) );
  INVX1 U1005 ( .A(n109), .Y(n1070) );
  INVX1 U1006 ( .A(n113), .Y(n1071) );
  AND2X1 U1007 ( .A(n1114), .B(n244), .Y(n110) );
  INVX1 U1008 ( .A(n110), .Y(n1072) );
  AND2X1 U1009 ( .A(n1096), .B(n1153), .Y(n86) );
  INVX1 U1010 ( .A(n86), .Y(n1073) );
  AND2X1 U1011 ( .A(n1112), .B(n130), .Y(n89) );
  INVX1 U1012 ( .A(n89), .Y(n1074) );
  AND2X1 U1013 ( .A(n342), .B(n351), .Y(n148) );
  INVX1 U1014 ( .A(n148), .Y(n1075) );
  OR2X1 U1015 ( .A(n376), .B(n389), .Y(n164) );
  INVX1 U1016 ( .A(n164), .Y(n1076) );
  AND2X1 U1017 ( .A(n558), .B(n557), .Y(n253) );
  INVX1 U1018 ( .A(n253), .Y(n1077) );
  AND2X1 U1019 ( .A(n488), .B(n477), .Y(n202) );
  INVX1 U1020 ( .A(n202), .Y(n1078) );
  INVX1 U1021 ( .A(n180), .Y(n1079) );
  BUFX2 U1022 ( .A(n187), .Y(n1080) );
  OR2X1 U1023 ( .A(n404), .B(n419), .Y(n174) );
  INVX1 U1024 ( .A(n174), .Y(n1081) );
  OR2X1 U1025 ( .A(n567), .B(n1219), .Y(n339) );
  INVX1 U1026 ( .A(n339), .Y(n1082) );
  AND2X2 U1027 ( .A(a[7]), .B(n1213), .Y(n1222) );
  INVX1 U1028 ( .A(n1222), .Y(n1083) );
  INVX1 U1029 ( .A(n1220), .Y(n1084) );
  INVX1 U1030 ( .A(n597), .Y(n1085) );
  INVX1 U1031 ( .A(n692), .Y(n1086) );
  AND2X1 U1032 ( .A(n1128), .B(n1152), .Y(n106) );
  INVX1 U1033 ( .A(n106), .Y(n1087) );
  AND2X1 U1034 ( .A(n1135), .B(n195), .Y(n101) );
  INVX1 U1035 ( .A(n101), .Y(n1088) );
  AND2X1 U1036 ( .A(n1110), .B(n1147), .Y(n105) );
  INVX1 U1037 ( .A(n105), .Y(n1089) );
  INVX1 U1038 ( .A(n96), .Y(n1090) );
  AND2X1 U1039 ( .A(n1138), .B(n204), .Y(n103) );
  INVX1 U1040 ( .A(n103), .Y(n1091) );
  AND2X1 U1041 ( .A(n1139), .B(n277), .Y(n99) );
  INVX1 U1042 ( .A(n99), .Y(n1092) );
  AND2X1 U1043 ( .A(n310), .B(n315), .Y(n128) );
  INVX1 U1044 ( .A(n128), .Y(n1093) );
  AND2X1 U1045 ( .A(n510), .B(n501), .Y(n213) );
  INVX1 U1046 ( .A(n213), .Y(n1094) );
  AND2X1 U1047 ( .A(n324), .B(n331), .Y(n136) );
  INVX1 U1048 ( .A(n136), .Y(n1095) );
  AND2X1 U1049 ( .A(n300), .B(n303), .Y(n120) );
  INVX1 U1050 ( .A(n120), .Y(n1096) );
  AND2X1 U1051 ( .A(n548), .B(n543), .Y(n242) );
  INVX1 U1052 ( .A(n242), .Y(n1097) );
  AND2X1 U1053 ( .A(n363), .B(n352), .Y(n153) );
  INVX1 U1054 ( .A(n153), .Y(n1098) );
  INVX1 U1055 ( .A(n259), .Y(n1099) );
  BUFX2 U1056 ( .A(n246), .Y(n1100) );
  AND2X1 U1057 ( .A(n389), .B(n376), .Y(n165) );
  INVX1 U1058 ( .A(n165), .Y(n1101) );
  OR2X1 U1059 ( .A(n477), .B(n488), .Y(n201) );
  INVX1 U1060 ( .A(n201), .Y(n1102) );
  OR2X1 U1061 ( .A(n420), .B(n434), .Y(n182) );
  INVX1 U1062 ( .A(n182), .Y(n1103) );
  OR2X1 U1063 ( .A(n449), .B(n462), .Y(n190) );
  OR2X1 U1064 ( .A(n565), .B(n999), .Y(n321) );
  INVX1 U1065 ( .A(n321), .Y(n1105) );
  AND2X1 U1066 ( .A(n1206), .B(n1177), .Y(n616) );
  INVX1 U1067 ( .A(n616), .Y(n1106) );
  INVX1 U1068 ( .A(n673), .Y(n1107) );
  AND2X1 U1069 ( .A(n1137), .B(n174), .Y(n97) );
  INVX1 U1070 ( .A(n97), .Y(n1108) );
  AND2X1 U1071 ( .A(n536), .B(n529), .Y(n231) );
  INVX1 U1072 ( .A(n231), .Y(n1109) );
  AND2X1 U1073 ( .A(n520), .B(n511), .Y(n218) );
  INVX1 U1074 ( .A(n218), .Y(n1110) );
  OR2X1 U1075 ( .A(n463), .B(n476), .Y(n195) );
  INVX1 U1076 ( .A(n195), .Y(n1111) );
  AND2X1 U1077 ( .A(n316), .B(n323), .Y(n131) );
  INVX1 U1078 ( .A(n131), .Y(n1112) );
  AND2X1 U1079 ( .A(n304), .B(n309), .Y(n123) );
  INVX1 U1080 ( .A(n123), .Y(n1113) );
  AND2X1 U1081 ( .A(n552), .B(n549), .Y(n245) );
  INVX1 U1082 ( .A(n245), .Y(n1114) );
  AND2X1 U1083 ( .A(n375), .B(n364), .Y(n160) );
  INVX1 U1084 ( .A(n160), .Y(n1115) );
  AND2X1 U1085 ( .A(n332), .B(n341), .Y(n139) );
  INVX1 U1086 ( .A(n139), .Y(n1116) );
  OR2X1 U1087 ( .A(n573), .B(n1219), .Y(n758) );
  INVX1 U1088 ( .A(n758), .Y(n1117) );
  BUFX2 U1089 ( .A(n254), .Y(n1118) );
  OR2X1 U1090 ( .A(n489), .B(n500), .Y(n204) );
  INVX1 U1091 ( .A(n204), .Y(n1119) );
  OR2X1 U1092 ( .A(n435), .B(n448), .Y(n185) );
  INVX1 U1093 ( .A(n185), .Y(n1120) );
  OR2X1 U1094 ( .A(n390), .B(n403), .Y(n171) );
  INVX1 U1095 ( .A(n171), .Y(n1121) );
  OR2X1 U1096 ( .A(n569), .B(n1219), .Y(n361) );
  INVX1 U1097 ( .A(n361), .Y(n1122) );
  AND2X1 U1098 ( .A(n1215), .B(n1214), .Y(n1223) );
  INVX1 U1099 ( .A(n1223), .Y(n1123) );
  AND2X1 U1100 ( .A(n1206), .B(n1209), .Y(n711) );
  INVX1 U1101 ( .A(n711), .Y(n1124) );
  INVX1 U1102 ( .A(n654), .Y(n1125) );
  INVX1 U1103 ( .A(n88), .Y(n1126) );
  INVX1 U1104 ( .A(n2), .Y(n1127) );
  AND2X1 U1105 ( .A(n528), .B(n521), .Y(n224) );
  INVX1 U1106 ( .A(n224), .Y(n1128) );
  AND2X1 U1107 ( .A(n542), .B(n537), .Y(n236) );
  INVX1 U1108 ( .A(n236), .Y(n1129) );
  OR2X1 U1109 ( .A(n309), .B(n304), .Y(n122) );
  INVX1 U1110 ( .A(n122), .Y(n1130) );
  OR2X1 U1111 ( .A(n549), .B(n552), .Y(n244) );
  INVX1 U1112 ( .A(n244), .Y(n1131) );
  OR2X1 U1113 ( .A(n323), .B(n316), .Y(n130) );
  INVX1 U1114 ( .A(n130), .Y(n1132) );
  OR2X1 U1115 ( .A(n557), .B(n558), .Y(n252) );
  INVX1 U1116 ( .A(n252), .Y(n1133) );
  OR2X1 U1117 ( .A(n341), .B(n332), .Y(n138) );
  INVX1 U1118 ( .A(n138), .Y(n1134) );
  AND2X1 U1119 ( .A(n476), .B(n463), .Y(n196) );
  INVX1 U1120 ( .A(n196), .Y(n1135) );
  INVX1 U1121 ( .A(n159), .Y(n1136) );
  AND2X1 U1122 ( .A(n419), .B(n404), .Y(n175) );
  INVX1 U1123 ( .A(n175), .Y(n1137) );
  AND2X1 U1124 ( .A(n500), .B(n489), .Y(n205) );
  INVX1 U1125 ( .A(n205), .Y(n1138) );
  AND2X1 U1126 ( .A(n448), .B(n435), .Y(n186) );
  INVX1 U1127 ( .A(n186), .Y(n1139) );
  OR2X1 U1128 ( .A(n571), .B(n1219), .Y(n387) );
  INVX1 U1129 ( .A(n387), .Y(n1140) );
  INVX1 U1130 ( .A(n262), .Y(n1141) );
  INVX2 U1131 ( .A(n735), .Y(n815) );
  AND2X2 U1132 ( .A(n1141), .B(n261), .Y(product[0]) );
  INVX1 U1133 ( .A(a[1]), .Y(n1142) );
  INVX2 U1134 ( .A(b[2]), .Y(n1194) );
  INVX2 U1135 ( .A(n741), .Y(n1143) );
  INVX1 U1136 ( .A(n170), .Y(n168) );
  INVX1 U1137 ( .A(n177), .Y(n176) );
  INVX1 U1138 ( .A(n1104), .Y(n278) );
  INVX1 U1139 ( .A(n1120), .Y(n277) );
  INVX1 U1140 ( .A(n207), .Y(n206) );
  INVX1 U1141 ( .A(n1008), .Y(n197) );
  INVX1 U1142 ( .A(n1005), .Y(n219) );
  INVX1 U1143 ( .A(n1007), .Y(n237) );
  OR2X1 U1144 ( .A(n352), .B(n363), .Y(n1144) );
  OR2X1 U1145 ( .A(n351), .B(n342), .Y(n1145) );
  OR2X1 U1146 ( .A(n537), .B(n542), .Y(n1146) );
  OR2X1 U1147 ( .A(n511), .B(n520), .Y(n1147) );
  OR2X1 U1148 ( .A(n501), .B(n510), .Y(n1149) );
  OR2X1 U1149 ( .A(n315), .B(n310), .Y(n1150) );
  OR2X1 U1150 ( .A(n331), .B(n324), .Y(n1151) );
  OR2X1 U1151 ( .A(n521), .B(n528), .Y(n1152) );
  BUFX2 U1152 ( .A(n44), .Y(n1186) );
  BUFX2 U1153 ( .A(n44), .Y(n1187) );
  INVX1 U1154 ( .A(n116), .Y(n263) );
  OR2X1 U1155 ( .A(n303), .B(n300), .Y(n1153) );
  OR2X1 U1156 ( .A(n543), .B(n548), .Y(n1155) );
  BUFX2 U1157 ( .A(n24), .Y(n1169) );
  BUFX2 U1158 ( .A(n18), .Y(n1165) );
  BUFX2 U1159 ( .A(n42), .Y(n1181) );
  BUFX2 U1160 ( .A(n36), .Y(n1177) );
  BUFX2 U1161 ( .A(n12), .Y(n1161) );
  BUFX2 U1162 ( .A(n30), .Y(n1173) );
  BUFX2 U1163 ( .A(n24), .Y(n1168) );
  BUFX2 U1164 ( .A(n18), .Y(n1164) );
  BUFX2 U1165 ( .A(n36), .Y(n1176) );
  BUFX2 U1166 ( .A(n30), .Y(n1172) );
  BUFX2 U1167 ( .A(n20), .Y(n1170) );
  BUFX2 U1168 ( .A(n14), .Y(n1166) );
  BUFX2 U1169 ( .A(n38), .Y(n1182) );
  BUFX2 U1170 ( .A(n8), .Y(n1162) );
  BUFX2 U1171 ( .A(n32), .Y(n1178) );
  BUFX2 U1172 ( .A(n26), .Y(n1174) );
  BUFX2 U1173 ( .A(n1127), .Y(n1158) );
  BUFX2 U1174 ( .A(n20), .Y(n1171) );
  BUFX2 U1175 ( .A(n14), .Y(n1167) );
  BUFX2 U1176 ( .A(n38), .Y(n1183) );
  BUFX2 U1177 ( .A(n8), .Y(n1163) );
  BUFX2 U1178 ( .A(n32), .Y(n1179) );
  BUFX2 U1179 ( .A(n26), .Y(n1175) );
  BUFX2 U1180 ( .A(n1127), .Y(n1159) );
  INVX1 U1181 ( .A(n1194), .Y(n1192) );
  INVX1 U1182 ( .A(n902), .Y(n260) );
  INVX1 U1183 ( .A(n1194), .Y(n1193) );
  INVX1 U1184 ( .A(n1216), .Y(n1215) );
  INVX1 U1185 ( .A(a[13]), .Y(n1218) );
  INVX1 U1186 ( .A(n1205), .Y(n1203) );
  INVX1 U1187 ( .A(n1197), .Y(n1195) );
  INVX1 U1188 ( .A(a[3]), .Y(n1212) );
  INVX1 U1189 ( .A(a[9]), .Y(n1216) );
  INVX1 U1190 ( .A(n1205), .Y(n1204) );
  INVX1 U1191 ( .A(n1202), .Y(n1201) );
  INVX1 U1192 ( .A(n1197), .Y(n1196) );
  INVX1 U1193 ( .A(b[14]), .Y(n1205) );
  INVX1 U1194 ( .A(b[13]), .Y(n1202) );
  INVX1 U1195 ( .A(b[11]), .Y(n1199) );
  INVX1 U1196 ( .A(b[6]), .Y(n1197) );
  INVX1 U1197 ( .A(a[0]), .Y(n1209) );
  OAI21X1 U1198 ( .A(a[2]), .B(n1212), .C(n1084), .Y(n741) );
  OAI21X1 U1199 ( .A(a[4]), .B(n1213), .C(n1049), .Y(n739) );
  OAI21X1 U1200 ( .A(a[6]), .B(n1214), .C(n1083), .Y(n737) );
  OAI21X1 U1201 ( .A(a[8]), .B(n1216), .C(n1123), .Y(n735) );
  OAI21X1 U1202 ( .A(a[10]), .B(n1217), .C(n1069), .Y(n733) );
  OAI21X1 U1203 ( .A(a[12]), .B(n1218), .C(n1052), .Y(n731) );
  OAI21X1 U1204 ( .A(a[14]), .B(n1219), .C(n1040), .Y(n729) );
  XOR2X1 U1205 ( .A(n1041), .B(n1058), .Y(n293) );
endmodule


module alu_DW_mult_uns_36 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n2, n8, n9, n12, n14, n18, n20, n24, n26, n30, n32, n36, n38, n42,
         n44, n48, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n115, n116, n120, n121, n122, n123, n124,
         n128, n129, n130, n131, n132, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n148, n149, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n163, n164, n165, n166, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n189, n190, n191, n192, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n213, n214, n218, n219, n220, n224, n225, n226, n227,
         n231, n232, n236, n237, n238, n242, n243, n244, n245, n246, n250,
         n251, n252, n253, n254, n258, n259, n260, n261, n262, n263, n273,
         n275, n276, n277, n293, n294, n295, n296, n297, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n576, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n595, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n614, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n633, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n652, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n671, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n690, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n709,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n728, n729, n731, n733, n735, n737,
         n739, n741, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247;

  FAX1 U87 ( .A(n296), .B(n299), .C(n263), .YC(n115), .YS(product[30]) );
  XNOR2X1 U89 ( .A(n1007), .B(n1146), .Y(product[29]) );
  AOI21X1 U90 ( .A(n121), .B(n1176), .C(n120), .Y(n116) );
  XOR2X1 U97 ( .A(n1064), .B(n1051), .Y(product[28]) );
  OAI21X1 U98 ( .A(n1149), .B(n1025), .C(n1130), .Y(n121) );
  XNOR2X1 U103 ( .A(n1004), .B(n1095), .Y(product[27]) );
  AOI21X1 U104 ( .A(n129), .B(n1170), .C(n128), .Y(n124) );
  XOR2X1 U111 ( .A(n1062), .B(n1096), .Y(product[26]) );
  OAI21X1 U112 ( .A(n1150), .B(n1063), .C(n1129), .Y(n129) );
  XNOR2X1 U117 ( .A(n1165), .B(n1145), .Y(product[25]) );
  AOI21X1 U118 ( .A(n137), .B(n1169), .C(n136), .Y(n132) );
  XOR2X1 U125 ( .A(n1059), .B(n1050), .Y(product[24]) );
  OAI21X1 U126 ( .A(n1151), .B(n1060), .C(n1131), .Y(n137) );
  XOR2X1 U131 ( .A(n1038), .B(n1049), .Y(product[23]) );
  AOI21X1 U132 ( .A(n177), .B(n1020), .C(n142), .Y(n140) );
  OAI21X1 U134 ( .A(n1056), .B(n1022), .C(n1032), .Y(n142) );
  AOI21X1 U136 ( .A(n1167), .B(n153), .C(n148), .Y(n144) );
  XNOR2X1 U143 ( .A(n154), .B(n1045), .Y(product[22]) );
  AOI21X1 U144 ( .A(n154), .B(n1168), .C(n153), .Y(n149) );
  XOR2X1 U151 ( .A(n1081), .B(n1080), .Y(product[21]) );
  OAI21X1 U152 ( .A(n1055), .B(n176), .C(n1022), .Y(n154) );
  AOI21X1 U154 ( .A(n170), .B(n1054), .C(n158), .Y(n156) );
  OAI21X1 U156 ( .A(n1135), .B(n1159), .C(n1115), .Y(n158) );
  XNOR2X1 U161 ( .A(n166), .B(n1044), .Y(product[20]) );
  AOI21X1 U162 ( .A(n166), .B(n273), .C(n163), .Y(n161) );
  XNOR2X1 U169 ( .A(n173), .B(n1084), .Y(product[19]) );
  OAI21X1 U170 ( .A(n169), .B(n176), .C(n168), .Y(n166) );
  OAI21X1 U174 ( .A(n1139), .B(n1160), .C(n1099), .Y(n170) );
  XOR2X1 U179 ( .A(n176), .B(n1097), .Y(product[18]) );
  OAI21X1 U180 ( .A(n1118), .B(n176), .C(n1139), .Y(n173) );
  XNOR2X1 U185 ( .A(n184), .B(n1043), .Y(product[17]) );
  OAI21X1 U187 ( .A(n1021), .B(n1024), .C(n1019), .Y(n177) );
  AOI21X1 U189 ( .A(n1028), .B(n189), .C(n181), .Y(n179) );
  OAI21X1 U191 ( .A(n1067), .B(n1157), .C(n1098), .Y(n181) );
  XOR2X1 U196 ( .A(n1057), .B(n1048), .Y(product[16]) );
  OAI21X1 U197 ( .A(n1138), .B(n1057), .C(n1067), .Y(n184) );
  XOR2X1 U202 ( .A(n1086), .B(n1085), .Y(product[15]) );
  AOI21X1 U203 ( .A(n197), .B(n1053), .C(n189), .Y(n187) );
  OAI21X1 U205 ( .A(n1100), .B(n1155), .C(n1114), .Y(n189) );
  XNOR2X1 U210 ( .A(n197), .B(n1042), .Y(product[14]) );
  AOI21X1 U211 ( .A(n197), .B(n195), .C(n196), .Y(n192) );
  XNOR2X1 U218 ( .A(n203), .B(n1094), .Y(product[13]) );
  AOI21X1 U220 ( .A(n207), .B(n1033), .C(n200), .Y(n198) );
  OAI21X1 U222 ( .A(n1162), .B(n1119), .C(n1089), .Y(n200) );
  XOR2X1 U227 ( .A(n206), .B(n1105), .Y(product[12]) );
  OAI21X1 U228 ( .A(n1136), .B(n206), .C(n1162), .Y(n203) );
  XOR2X1 U233 ( .A(n1037), .B(n1047), .Y(product[11]) );
  OAI21X1 U235 ( .A(n1017), .B(n1026), .C(n1031), .Y(n207) );
  AOI21X1 U237 ( .A(n1175), .B(n218), .C(n213), .Y(n209) );
  XNOR2X1 U244 ( .A(n219), .B(n1123), .Y(product[10]) );
  AOI21X1 U245 ( .A(n219), .B(n1173), .C(n218), .Y(n214) );
  XNOR2X1 U252 ( .A(n225), .B(n1041), .Y(product[9]) );
  AOI21X1 U254 ( .A(n999), .B(n1177), .C(n224), .Y(n220) );
  XOR2X1 U261 ( .A(n1036), .B(n1046), .Y(product[8]) );
  OAI21X1 U262 ( .A(n1016), .B(n1023), .C(n1030), .Y(n225) );
  AOI21X1 U264 ( .A(n236), .B(n1174), .C(n231), .Y(n227) );
  XNOR2X1 U271 ( .A(n237), .B(n1040), .Y(product[7]) );
  AOI21X1 U272 ( .A(n237), .B(n1172), .C(n236), .Y(n232) );
  XNOR2X1 U279 ( .A(n1144), .B(n1166), .Y(product[6]) );
  AOI21X1 U281 ( .A(n243), .B(n1179), .C(n242), .Y(n238) );
  XOR2X1 U288 ( .A(n1039), .B(n1015), .Y(product[5]) );
  OAI21X1 U289 ( .A(n1152), .B(n1066), .C(n1132), .Y(n243) );
  XNOR2X1 U294 ( .A(n1035), .B(n1008), .Y(product[4]) );
  AOI21X1 U295 ( .A(n251), .B(n1180), .C(n250), .Y(n246) );
  XOR2X1 U302 ( .A(n1093), .B(n1116), .Y(product[3]) );
  OAI21X1 U303 ( .A(n1153), .B(n1116), .C(n1133), .Y(n251) );
  XNOR2X1 U308 ( .A(n1092), .B(n1134), .Y(product[2]) );
  AOI21X1 U309 ( .A(n1171), .B(n1012), .C(n258), .Y(n254) );
  XOR2X1 U316 ( .A(n260), .B(n1164), .Y(product[1]) );
  XOR2X1 U324 ( .A(n761), .B(n293), .Y(n294) );
  FAX1 U326 ( .A(n297), .B(n762), .C(n301), .YC(n295), .YS(n296) );
  FAX1 U328 ( .A(n763), .B(n302), .C(n305), .YC(n299), .YS(n300) );
  FAX1 U329 ( .A(n779), .B(n1090), .C(n1070), .YC(n301), .YS(n302) );
  FAX1 U330 ( .A(n313), .B(n306), .C(n311), .YC(n303), .YS(n304) );
  FAX1 U331 ( .A(n307), .B(n780), .C(n764), .YC(n305), .YS(n306) );
  FAX1 U333 ( .A(n319), .B(n312), .C(n317), .YC(n309), .YS(n310) );
  FAX1 U334 ( .A(n781), .B(n765), .C(n314), .YC(n311), .YS(n312) );
  FAX1 U335 ( .A(n797), .B(n1101), .C(n1072), .YC(n313), .YS(n314) );
  FAX1 U336 ( .A(n327), .B(n318), .C(n325), .YC(n315), .YS(n316) );
  FAX1 U337 ( .A(n766), .B(n329), .C(n320), .YC(n317), .YS(n318) );
  FAX1 U338 ( .A(n321), .B(n798), .C(n782), .YC(n319), .YS(n320) );
  FAX1 U340 ( .A(n328), .B(n326), .C(n333), .YC(n323), .YS(n324) );
  FAX1 U341 ( .A(n330), .B(n337), .C(n335), .YC(n325), .YS(n326) );
  FAX1 U342 ( .A(n783), .B(n799), .C(n767), .YC(n327), .YS(n328) );
  FAX1 U343 ( .A(n815), .B(n1120), .C(n1071), .YC(n329), .YS(n330) );
  FAX1 U344 ( .A(n345), .B(n334), .C(n343), .YC(n331), .YS(n332) );
  FAX1 U345 ( .A(n338), .B(n347), .C(n336), .YC(n333), .YS(n334) );
  FAX1 U346 ( .A(n800), .B(n768), .C(n349), .YC(n335), .YS(n336) );
  FAX1 U347 ( .A(n339), .B(n816), .C(n784), .YC(n337), .YS(n338) );
  FAX1 U349 ( .A(n355), .B(n344), .C(n353), .YC(n341), .YS(n342) );
  FAX1 U350 ( .A(n357), .B(n348), .C(n346), .YC(n343), .YS(n344) );
  FAX1 U351 ( .A(n785), .B(n350), .C(n359), .YC(n345), .YS(n346) );
  FAX1 U352 ( .A(n817), .B(n801), .C(n769), .YC(n347), .YS(n348) );
  FAX1 U353 ( .A(n833), .B(n1163), .C(n1074), .YC(n349), .YS(n350) );
  FAX1 U354 ( .A(n367), .B(n354), .C(n365), .YC(n351), .YS(n352) );
  FAX1 U355 ( .A(n358), .B(n369), .C(n356), .YC(n353), .YS(n354) );
  FAX1 U356 ( .A(n373), .B(n360), .C(n371), .YC(n355), .YS(n356) );
  FAX1 U357 ( .A(n786), .B(n802), .C(n770), .YC(n357), .YS(n358) );
  FAX1 U358 ( .A(n361), .B(n834), .C(n818), .YC(n359), .YS(n360) );
  FAX1 U360 ( .A(n368), .B(n377), .C(n366), .YC(n363), .YS(n364) );
  FAX1 U361 ( .A(n370), .B(n381), .C(n379), .YC(n365), .YS(n366) );
  FAX1 U362 ( .A(n385), .B(n383), .C(n372), .YC(n367), .YS(n368) );
  FAX1 U363 ( .A(n787), .B(n835), .C(n374), .YC(n369), .YS(n370) );
  FAX1 U364 ( .A(n819), .B(n803), .C(n771), .YC(n371), .YS(n372) );
  FAX1 U365 ( .A(n851), .B(n1140), .C(n1076), .YC(n373), .YS(n374) );
  FAX1 U366 ( .A(n380), .B(n391), .C(n378), .YC(n375), .YS(n376) );
  FAX1 U367 ( .A(n382), .B(n395), .C(n393), .YC(n377), .YS(n378) );
  FAX1 U368 ( .A(n397), .B(n399), .C(n384), .YC(n379), .YS(n380) );
  FAX1 U369 ( .A(n836), .B(n804), .C(n386), .YC(n381), .YS(n382) );
  FAX1 U370 ( .A(n401), .B(n772), .C(n788), .YC(n383), .YS(n384) );
  FAX1 U371 ( .A(n387), .B(n852), .C(n820), .YC(n385), .YS(n386) );
  FAX1 U373 ( .A(n394), .B(n405), .C(n392), .YC(n389), .YS(n390) );
  FAX1 U374 ( .A(n409), .B(n396), .C(n407), .YC(n391), .YS(n392) );
  FAX1 U375 ( .A(n411), .B(n400), .C(n398), .YC(n393), .YS(n394) );
  FAX1 U376 ( .A(n789), .B(n415), .C(n413), .YC(n395), .YS(n396) );
  FAX1 U377 ( .A(n853), .B(n837), .C(n805), .YC(n397), .YS(n398) );
  FAX1 U378 ( .A(n821), .B(n402), .C(n773), .YC(n399), .YS(n400) );
  FAX1 U379 ( .A(n1228), .B(n9), .C(n1075), .YC(n401), .YS(n402) );
  FAX1 U380 ( .A(n408), .B(n421), .C(n406), .YC(n403), .YS(n404) );
  FAX1 U381 ( .A(n425), .B(n410), .C(n423), .YC(n405), .YS(n406) );
  FAX1 U382 ( .A(n427), .B(n414), .C(n412), .YC(n407), .YS(n408) );
  FAX1 U383 ( .A(n416), .B(n431), .C(n429), .YC(n409), .YS(n410) );
  FAX1 U384 ( .A(n854), .B(n838), .C(n790), .YC(n411), .YS(n412) );
  FAX1 U385 ( .A(n822), .B(n806), .C(n774), .YC(n413), .YS(n414) );
  FAX1 U386 ( .A(a[1]), .B(n1154), .C(n870), .YC(n415), .YS(n416) );
  FAX1 U388 ( .A(n424), .B(n436), .C(n422), .YC(n419), .YS(n420) );
  FAX1 U389 ( .A(n440), .B(n426), .C(n438), .YC(n421), .YS(n422) );
  FAX1 U390 ( .A(n444), .B(n430), .C(n428), .YC(n423), .YS(n424) );
  FAX1 U391 ( .A(n446), .B(n432), .C(n442), .YC(n425), .YS(n426) );
  FAX1 U392 ( .A(n855), .B(n839), .C(n791), .YC(n427), .YS(n428) );
  FAX1 U393 ( .A(n823), .B(n807), .C(n775), .YC(n429), .YS(n430) );
  FAX1 U394 ( .A(a[1]), .B(n1077), .C(n871), .YC(n431), .YS(n432) );
  FAX1 U396 ( .A(n439), .B(n450), .C(n437), .YC(n434), .YS(n435) );
  FAX1 U397 ( .A(n454), .B(n441), .C(n452), .YC(n436), .YS(n437) );
  FAX1 U398 ( .A(n456), .B(n445), .C(n443), .YC(n438), .YS(n439) );
  FAX1 U399 ( .A(n460), .B(n447), .C(n458), .YC(n440), .YS(n441) );
  FAX1 U400 ( .A(n856), .B(n840), .C(n792), .YC(n442), .YS(n443) );
  FAX1 U401 ( .A(n824), .B(n808), .C(n776), .YC(n444), .YS(n445) );
  FAX1 U402 ( .A(n887), .B(n1078), .C(n872), .YC(n446), .YS(n447) );
  FAX1 U403 ( .A(n453), .B(n464), .C(n451), .YC(n448), .YS(n449) );
  FAX1 U404 ( .A(n468), .B(n455), .C(n466), .YC(n450), .YS(n451) );
  FAX1 U405 ( .A(n470), .B(n459), .C(n457), .YC(n452), .YS(n453) );
  FAX1 U406 ( .A(n793), .B(n461), .C(n472), .YC(n454), .YS(n455) );
  FAX1 U407 ( .A(n857), .B(n841), .C(n809), .YC(n456), .YS(n457) );
  FAX1 U408 ( .A(n825), .B(n777), .C(n474), .YC(n458), .YS(n459) );
  HAX1 U409 ( .A(n888), .B(n873), .YC(n460), .YS(n461) );
  FAX1 U410 ( .A(n467), .B(n478), .C(n465), .YC(n462), .YS(n463) );
  FAX1 U411 ( .A(n482), .B(n469), .C(n480), .YC(n464), .YS(n465) );
  FAX1 U412 ( .A(n484), .B(n473), .C(n471), .YC(n466), .YS(n467) );
  FAX1 U413 ( .A(n826), .B(n858), .C(n486), .YC(n468), .YS(n469) );
  FAX1 U414 ( .A(n874), .B(n794), .C(n475), .YC(n470), .YS(n471) );
  FAX1 U415 ( .A(n778), .B(n842), .C(n810), .YC(n472), .YS(n473) );
  HAX1 U416 ( .A(n889), .B(n743), .YC(n474), .YS(n475) );
  FAX1 U417 ( .A(n481), .B(n490), .C(n479), .YC(n476), .YS(n477) );
  FAX1 U418 ( .A(n485), .B(n483), .C(n492), .YC(n478), .YS(n479) );
  FAX1 U419 ( .A(n487), .B(n496), .C(n494), .YC(n480), .YS(n481) );
  FAX1 U420 ( .A(n859), .B(n795), .C(n843), .YC(n482), .YS(n483) );
  FAX1 U421 ( .A(n827), .B(n811), .C(n498), .YC(n484), .YS(n485) );
  HAX1 U422 ( .A(n890), .B(n875), .YC(n486), .YS(n487) );
  FAX1 U423 ( .A(n493), .B(n502), .C(n491), .YC(n488), .YS(n489) );
  FAX1 U424 ( .A(n497), .B(n495), .C(n504), .YC(n490), .YS(n491) );
  FAX1 U425 ( .A(n828), .B(n508), .C(n506), .YC(n492), .YS(n493) );
  FAX1 U426 ( .A(n876), .B(n860), .C(n499), .YC(n494), .YS(n495) );
  FAX1 U427 ( .A(n796), .B(n844), .C(n812), .YC(n496), .YS(n497) );
  HAX1 U428 ( .A(n744), .B(n891), .YC(n498), .YS(n499) );
  FAX1 U429 ( .A(n505), .B(n512), .C(n503), .YC(n500), .YS(n501) );
  FAX1 U430 ( .A(n516), .B(n514), .C(n507), .YC(n502), .YS(n503) );
  FAX1 U431 ( .A(n861), .B(n845), .C(n509), .YC(n504), .YS(n505) );
  FAX1 U432 ( .A(n829), .B(n813), .C(n518), .YC(n506), .YS(n507) );
  HAX1 U433 ( .A(n892), .B(n877), .YC(n508), .YS(n509) );
  FAX1 U434 ( .A(n515), .B(n522), .C(n513), .YC(n510), .YS(n511) );
  FAX1 U435 ( .A(n526), .B(n524), .C(n517), .YC(n512), .YS(n513) );
  FAX1 U436 ( .A(n878), .B(n830), .C(n519), .YC(n514), .YS(n515) );
  FAX1 U437 ( .A(n814), .B(n862), .C(n846), .YC(n516), .YS(n517) );
  HAX1 U438 ( .A(n893), .B(n745), .YC(n518), .YS(n519) );
  FAX1 U439 ( .A(n525), .B(n530), .C(n523), .YC(n520), .YS(n521) );
  FAX1 U440 ( .A(n863), .B(n527), .C(n532), .YC(n522), .YS(n523) );
  FAX1 U441 ( .A(n831), .B(n847), .C(n534), .YC(n524), .YS(n525) );
  HAX1 U442 ( .A(n894), .B(n879), .YC(n526), .YS(n527) );
  FAX1 U443 ( .A(n538), .B(n533), .C(n531), .YC(n528), .YS(n529) );
  FAX1 U444 ( .A(n880), .B(n535), .C(n540), .YC(n530), .YS(n531) );
  FAX1 U445 ( .A(n832), .B(n864), .C(n848), .YC(n532), .YS(n533) );
  HAX1 U446 ( .A(n895), .B(n746), .YC(n534), .YS(n535) );
  FAX1 U447 ( .A(n541), .B(n544), .C(n539), .YC(n536), .YS(n537) );
  FAX1 U448 ( .A(n546), .B(n849), .C(n865), .YC(n538), .YS(n539) );
  HAX1 U449 ( .A(n896), .B(n881), .YC(n540), .YS(n541) );
  FAX1 U450 ( .A(n547), .B(n550), .C(n545), .YC(n542), .YS(n543) );
  FAX1 U451 ( .A(n866), .B(n882), .C(n850), .YC(n544), .YS(n545) );
  HAX1 U452 ( .A(n897), .B(n747), .YC(n546), .YS(n547) );
  FAX1 U453 ( .A(n867), .B(n554), .C(n551), .YC(n548), .YS(n549) );
  HAX1 U454 ( .A(n898), .B(n883), .YC(n550), .YS(n551) );
  FAX1 U455 ( .A(n868), .B(n884), .C(n555), .YC(n552), .YS(n553) );
  HAX1 U456 ( .A(n899), .B(n748), .YC(n554), .YS(n555) );
  HAX1 U457 ( .A(n900), .B(n885), .YC(n556), .YS(n557) );
  HAX1 U458 ( .A(n901), .B(n749), .YC(n558), .YS(n559) );
  MUX2X1 U460 ( .B(b[15]), .A(b[14]), .S(n1238), .Y(n560) );
  MUX2X1 U462 ( .B(b[14]), .A(b[13]), .S(n1238), .Y(n561) );
  MUX2X1 U464 ( .B(b[13]), .A(n1223), .S(n1238), .Y(n562) );
  MUX2X1 U466 ( .B(n1223), .A(b[11]), .S(n1238), .Y(n563) );
  MUX2X1 U468 ( .B(b[11]), .A(n1220), .S(n1238), .Y(n564) );
  MUX2X1 U470 ( .B(n1220), .A(n1217), .S(n1238), .Y(n565) );
  MUX2X1 U472 ( .B(n1217), .A(b[8]), .S(n1238), .Y(n566) );
  MUX2X1 U474 ( .B(b[8]), .A(b[7]), .S(n1238), .Y(n567) );
  MUX2X1 U476 ( .B(b[7]), .A(b[6]), .S(n1239), .Y(n568) );
  MUX2X1 U478 ( .B(b[6]), .A(b[5]), .S(n1239), .Y(n569) );
  MUX2X1 U480 ( .B(b[5]), .A(b[4]), .S(n1239), .Y(n570) );
  MUX2X1 U482 ( .B(b[4]), .A(b[3]), .S(n1238), .Y(n571) );
  MUX2X1 U484 ( .B(b[3]), .A(n1215), .S(n1238), .Y(n572) );
  MUX2X1 U486 ( .B(n1215), .A(n1212), .S(n1238), .Y(n573) );
  MUX2X1 U488 ( .B(n1212), .A(n1210), .S(n1238), .Y(n574) );
  AND2X1 U492 ( .A(n1209), .B(n729), .Y(n743) );
  MUX2X1 U495 ( .B(n1209), .A(n761), .S(n1034), .Y(n762) );
  MUX2X1 U497 ( .B(n1209), .A(n761), .S(n579), .Y(n763) );
  MUX2X1 U498 ( .B(b[15]), .A(b[14]), .S(n1207), .Y(n579) );
  MUX2X1 U499 ( .B(n1209), .A(n761), .S(n580), .Y(n764) );
  MUX2X1 U500 ( .B(b[14]), .A(b[13]), .S(n1207), .Y(n580) );
  MUX2X1 U501 ( .B(n1209), .A(n761), .S(n581), .Y(n765) );
  MUX2X1 U502 ( .B(b[13]), .A(n1223), .S(n1207), .Y(n581) );
  MUX2X1 U503 ( .B(n1209), .A(n761), .S(n582), .Y(n766) );
  MUX2X1 U504 ( .B(n1223), .A(b[11]), .S(n1207), .Y(n582) );
  MUX2X1 U505 ( .B(n1209), .A(n761), .S(n583), .Y(n767) );
  MUX2X1 U506 ( .B(b[11]), .A(n1220), .S(n1207), .Y(n583) );
  MUX2X1 U507 ( .B(n1209), .A(n761), .S(n584), .Y(n768) );
  MUX2X1 U508 ( .B(n1220), .A(n1217), .S(n1207), .Y(n584) );
  MUX2X1 U509 ( .B(n1209), .A(n761), .S(n585), .Y(n769) );
  MUX2X1 U510 ( .B(n1217), .A(b[8]), .S(n1207), .Y(n585) );
  MUX2X1 U511 ( .B(n1208), .A(n761), .S(n586), .Y(n770) );
  MUX2X1 U512 ( .B(b[8]), .A(b[7]), .S(n1206), .Y(n586) );
  MUX2X1 U513 ( .B(n1208), .A(n761), .S(n587), .Y(n771) );
  MUX2X1 U514 ( .B(b[7]), .A(b[6]), .S(n1206), .Y(n587) );
  MUX2X1 U515 ( .B(n1208), .A(n761), .S(n588), .Y(n772) );
  MUX2X1 U516 ( .B(b[6]), .A(b[5]), .S(n1206), .Y(n588) );
  MUX2X1 U517 ( .B(n1208), .A(n761), .S(n589), .Y(n773) );
  MUX2X1 U518 ( .B(b[5]), .A(b[4]), .S(n1206), .Y(n589) );
  MUX2X1 U519 ( .B(n1208), .A(n761), .S(n590), .Y(n774) );
  MUX2X1 U520 ( .B(b[4]), .A(b[3]), .S(n1206), .Y(n590) );
  MUX2X1 U521 ( .B(n1208), .A(n761), .S(n591), .Y(n775) );
  MUX2X1 U522 ( .B(b[3]), .A(n1215), .S(n1206), .Y(n591) );
  MUX2X1 U523 ( .B(n1208), .A(n761), .S(n592), .Y(n776) );
  MUX2X1 U524 ( .B(n1215), .A(n1212), .S(n1206), .Y(n592) );
  MUX2X1 U525 ( .B(n1208), .A(n761), .S(n593), .Y(n777) );
  MUX2X1 U526 ( .B(n1212), .A(n1210), .S(n1206), .Y(n593) );
  MUX2X1 U527 ( .B(n1208), .A(n761), .S(n595), .Y(n778) );
  AND2X1 U530 ( .A(n1205), .B(n731), .Y(n744) );
  MUX2X1 U533 ( .B(n1205), .A(n779), .S(n1103), .Y(n780) );
  MUX2X1 U535 ( .B(n1205), .A(n779), .S(n598), .Y(n781) );
  MUX2X1 U536 ( .B(b[15]), .A(b[14]), .S(n1203), .Y(n598) );
  MUX2X1 U537 ( .B(n1205), .A(n779), .S(n599), .Y(n782) );
  MUX2X1 U538 ( .B(b[14]), .A(b[13]), .S(n1203), .Y(n599) );
  MUX2X1 U539 ( .B(n1205), .A(n779), .S(n600), .Y(n783) );
  MUX2X1 U540 ( .B(b[13]), .A(n1223), .S(n1203), .Y(n600) );
  MUX2X1 U541 ( .B(n1205), .A(n779), .S(n601), .Y(n784) );
  MUX2X1 U542 ( .B(n1224), .A(b[11]), .S(n1203), .Y(n601) );
  MUX2X1 U543 ( .B(n1205), .A(n779), .S(n602), .Y(n785) );
  MUX2X1 U544 ( .B(b[11]), .A(n1220), .S(n1203), .Y(n602) );
  MUX2X1 U545 ( .B(n1205), .A(n779), .S(n603), .Y(n786) );
  MUX2X1 U546 ( .B(n1221), .A(n1217), .S(n1203), .Y(n603) );
  MUX2X1 U547 ( .B(n1205), .A(n779), .S(n604), .Y(n787) );
  MUX2X1 U548 ( .B(n1218), .A(b[8]), .S(n1203), .Y(n604) );
  MUX2X1 U549 ( .B(n1204), .A(n779), .S(n605), .Y(n788) );
  MUX2X1 U550 ( .B(b[8]), .A(b[7]), .S(n1202), .Y(n605) );
  MUX2X1 U551 ( .B(n1204), .A(n779), .S(n606), .Y(n789) );
  MUX2X1 U552 ( .B(b[7]), .A(b[6]), .S(n1202), .Y(n606) );
  MUX2X1 U553 ( .B(n1204), .A(n779), .S(n607), .Y(n790) );
  MUX2X1 U554 ( .B(b[6]), .A(b[5]), .S(n1202), .Y(n607) );
  MUX2X1 U555 ( .B(n1204), .A(n779), .S(n608), .Y(n791) );
  MUX2X1 U556 ( .B(b[5]), .A(b[4]), .S(n1202), .Y(n608) );
  MUX2X1 U557 ( .B(n1204), .A(n779), .S(n609), .Y(n792) );
  MUX2X1 U558 ( .B(b[4]), .A(b[3]), .S(n1202), .Y(n609) );
  MUX2X1 U559 ( .B(n1204), .A(n779), .S(n610), .Y(n793) );
  MUX2X1 U560 ( .B(n998), .A(n1215), .S(n1202), .Y(n610) );
  MUX2X1 U561 ( .B(n1204), .A(n779), .S(n611), .Y(n794) );
  MUX2X1 U562 ( .B(n1215), .A(n1212), .S(n1202), .Y(n611) );
  MUX2X1 U563 ( .B(n1204), .A(n779), .S(n612), .Y(n795) );
  MUX2X1 U564 ( .B(n1213), .A(n1210), .S(n1202), .Y(n612) );
  MUX2X1 U565 ( .B(n1204), .A(n779), .S(n614), .Y(n796) );
  MUX2X1 U571 ( .B(n1201), .A(n797), .S(n1104), .Y(n798) );
  MUX2X1 U573 ( .B(n1201), .A(n797), .S(n617), .Y(n799) );
  MUX2X1 U574 ( .B(b[15]), .A(b[14]), .S(n1003), .Y(n617) );
  MUX2X1 U575 ( .B(n1201), .A(n797), .S(n618), .Y(n800) );
  MUX2X1 U576 ( .B(b[14]), .A(b[13]), .S(n1003), .Y(n618) );
  MUX2X1 U577 ( .B(n1201), .A(n797), .S(n619), .Y(n801) );
  MUX2X1 U578 ( .B(b[13]), .A(n1223), .S(n1003), .Y(n619) );
  MUX2X1 U579 ( .B(n1201), .A(n797), .S(n620), .Y(n802) );
  MUX2X1 U580 ( .B(n1224), .A(b[11]), .S(n1003), .Y(n620) );
  MUX2X1 U581 ( .B(n1201), .A(n797), .S(n621), .Y(n803) );
  MUX2X1 U582 ( .B(b[11]), .A(n1220), .S(n1003), .Y(n621) );
  MUX2X1 U583 ( .B(n1201), .A(n797), .S(n622), .Y(n804) );
  MUX2X1 U584 ( .B(n1221), .A(n1217), .S(n1003), .Y(n622) );
  MUX2X1 U585 ( .B(n1201), .A(n797), .S(n623), .Y(n805) );
  MUX2X1 U586 ( .B(n1218), .A(b[8]), .S(n1002), .Y(n623) );
  MUX2X1 U587 ( .B(n1200), .A(n797), .S(n624), .Y(n806) );
  MUX2X1 U588 ( .B(b[8]), .A(b[7]), .S(n1198), .Y(n624) );
  MUX2X1 U589 ( .B(n1200), .A(n797), .S(n625), .Y(n807) );
  MUX2X1 U590 ( .B(b[7]), .A(b[6]), .S(n1198), .Y(n625) );
  MUX2X1 U591 ( .B(n1200), .A(n797), .S(n626), .Y(n808) );
  MUX2X1 U592 ( .B(b[6]), .A(b[5]), .S(n1198), .Y(n626) );
  MUX2X1 U593 ( .B(n1200), .A(n797), .S(n627), .Y(n809) );
  MUX2X1 U594 ( .B(b[5]), .A(b[4]), .S(n1198), .Y(n627) );
  MUX2X1 U595 ( .B(n1200), .A(n797), .S(n628), .Y(n810) );
  MUX2X1 U596 ( .B(b[4]), .A(b[3]), .S(n1198), .Y(n628) );
  MUX2X1 U597 ( .B(n1200), .A(n797), .S(n629), .Y(n811) );
  MUX2X1 U598 ( .B(b[3]), .A(n1215), .S(n1198), .Y(n629) );
  MUX2X1 U599 ( .B(n1200), .A(n797), .S(n630), .Y(n812) );
  MUX2X1 U600 ( .B(n1215), .A(n1212), .S(n1198), .Y(n630) );
  MUX2X1 U601 ( .B(n1200), .A(n797), .S(n631), .Y(n813) );
  MUX2X1 U602 ( .B(n1213), .A(n1210), .S(n1198), .Y(n631) );
  MUX2X1 U603 ( .B(n1200), .A(n797), .S(n633), .Y(n814) );
  AND2X1 U606 ( .A(n1197), .B(n735), .Y(n746) );
  MUX2X1 U609 ( .B(n1197), .A(n815), .S(n1142), .Y(n816) );
  MUX2X1 U611 ( .B(n1197), .A(n815), .S(n636), .Y(n817) );
  MUX2X1 U612 ( .B(b[15]), .A(b[14]), .S(n1194), .Y(n636) );
  MUX2X1 U613 ( .B(n1197), .A(n815), .S(n637), .Y(n818) );
  MUX2X1 U614 ( .B(b[14]), .A(b[13]), .S(n1194), .Y(n637) );
  MUX2X1 U615 ( .B(n1197), .A(n815), .S(n638), .Y(n819) );
  MUX2X1 U616 ( .B(b[13]), .A(n1223), .S(n1194), .Y(n638) );
  MUX2X1 U617 ( .B(n1197), .A(n815), .S(n639), .Y(n820) );
  MUX2X1 U618 ( .B(n1223), .A(b[11]), .S(n1195), .Y(n639) );
  MUX2X1 U619 ( .B(n1197), .A(n815), .S(n640), .Y(n821) );
  MUX2X1 U620 ( .B(b[11]), .A(n1220), .S(n1195), .Y(n640) );
  MUX2X1 U621 ( .B(n1197), .A(n815), .S(n641), .Y(n822) );
  MUX2X1 U622 ( .B(n1220), .A(n1217), .S(n1195), .Y(n641) );
  MUX2X1 U623 ( .B(n1197), .A(n815), .S(n642), .Y(n823) );
  MUX2X1 U624 ( .B(n1217), .A(b[8]), .S(n1195), .Y(n642) );
  MUX2X1 U625 ( .B(n1196), .A(n815), .S(n643), .Y(n824) );
  MUX2X1 U626 ( .B(b[8]), .A(b[7]), .S(n1195), .Y(n643) );
  MUX2X1 U627 ( .B(n1196), .A(n815), .S(n644), .Y(n825) );
  MUX2X1 U628 ( .B(b[7]), .A(b[6]), .S(n1195), .Y(n644) );
  MUX2X1 U629 ( .B(n1196), .A(n815), .S(n645), .Y(n826) );
  MUX2X1 U630 ( .B(b[6]), .A(b[5]), .S(n1194), .Y(n645) );
  MUX2X1 U631 ( .B(n1196), .A(n815), .S(n646), .Y(n827) );
  MUX2X1 U632 ( .B(b[5]), .A(b[4]), .S(n1194), .Y(n646) );
  MUX2X1 U633 ( .B(n1196), .A(n815), .S(n647), .Y(n828) );
  MUX2X1 U634 ( .B(b[4]), .A(n998), .S(n1194), .Y(n647) );
  MUX2X1 U635 ( .B(n1196), .A(n815), .S(n648), .Y(n829) );
  MUX2X1 U636 ( .B(b[3]), .A(n1215), .S(n1194), .Y(n648) );
  MUX2X1 U637 ( .B(n1196), .A(n815), .S(n649), .Y(n830) );
  MUX2X1 U638 ( .B(n1215), .A(n1212), .S(n1194), .Y(n649) );
  MUX2X1 U639 ( .B(n1196), .A(n815), .S(n650), .Y(n831) );
  MUX2X1 U640 ( .B(n1212), .A(n1210), .S(n1194), .Y(n650) );
  MUX2X1 U641 ( .B(n1196), .A(n815), .S(n652), .Y(n832) );
  MUX2X1 U647 ( .B(n1193), .A(n833), .S(n1122), .Y(n834) );
  MUX2X1 U649 ( .B(n1193), .A(n833), .S(n655), .Y(n835) );
  MUX2X1 U650 ( .B(b[15]), .A(b[14]), .S(n1191), .Y(n655) );
  MUX2X1 U651 ( .B(n1193), .A(n833), .S(n656), .Y(n836) );
  MUX2X1 U652 ( .B(b[14]), .A(b[13]), .S(n1191), .Y(n656) );
  MUX2X1 U653 ( .B(n1193), .A(n833), .S(n657), .Y(n837) );
  MUX2X1 U654 ( .B(b[13]), .A(n1223), .S(n1190), .Y(n657) );
  MUX2X1 U655 ( .B(n1193), .A(n833), .S(n658), .Y(n838) );
  MUX2X1 U656 ( .B(n1223), .A(b[11]), .S(n1190), .Y(n658) );
  MUX2X1 U657 ( .B(n1193), .A(n833), .S(n659), .Y(n839) );
  MUX2X1 U658 ( .B(b[11]), .A(n1220), .S(n1190), .Y(n659) );
  MUX2X1 U659 ( .B(n1193), .A(n833), .S(n660), .Y(n840) );
  MUX2X1 U660 ( .B(n1220), .A(n1217), .S(n1191), .Y(n660) );
  MUX2X1 U661 ( .B(n1193), .A(n833), .S(n661), .Y(n841) );
  MUX2X1 U662 ( .B(n1217), .A(b[8]), .S(n1190), .Y(n661) );
  MUX2X1 U663 ( .B(n1192), .A(n833), .S(n662), .Y(n842) );
  MUX2X1 U664 ( .B(b[8]), .A(b[7]), .S(n1190), .Y(n662) );
  MUX2X1 U665 ( .B(n1192), .A(n833), .S(n663), .Y(n843) );
  MUX2X1 U666 ( .B(b[7]), .A(b[6]), .S(n1191), .Y(n663) );
  MUX2X1 U667 ( .B(n1192), .A(n833), .S(n664), .Y(n844) );
  MUX2X1 U668 ( .B(b[6]), .A(b[5]), .S(n1191), .Y(n664) );
  MUX2X1 U669 ( .B(n1192), .A(n833), .S(n665), .Y(n845) );
  MUX2X1 U670 ( .B(b[5]), .A(b[4]), .S(n1191), .Y(n665) );
  MUX2X1 U671 ( .B(n1192), .A(n833), .S(n666), .Y(n846) );
  MUX2X1 U672 ( .B(b[4]), .A(n998), .S(n1191), .Y(n666) );
  MUX2X1 U673 ( .B(n1192), .A(n833), .S(n667), .Y(n847) );
  MUX2X1 U674 ( .B(n998), .A(n1215), .S(n1191), .Y(n667) );
  MUX2X1 U675 ( .B(n1192), .A(n833), .S(n668), .Y(n848) );
  MUX2X1 U676 ( .B(n1215), .A(n1212), .S(n1191), .Y(n668) );
  MUX2X1 U677 ( .B(n1192), .A(n833), .S(n669), .Y(n849) );
  MUX2X1 U678 ( .B(n1212), .A(n1210), .S(n1190), .Y(n669) );
  MUX2X1 U679 ( .B(n1192), .A(n833), .S(n671), .Y(n850) );
  AND2X1 U682 ( .A(n1189), .B(n739), .Y(n748) );
  MUX2X1 U685 ( .B(n1189), .A(n851), .S(n1143), .Y(n852) );
  MUX2X1 U687 ( .B(n1189), .A(n851), .S(n674), .Y(n853) );
  MUX2X1 U688 ( .B(b[15]), .A(b[14]), .S(n1187), .Y(n674) );
  MUX2X1 U689 ( .B(n1189), .A(n851), .S(n675), .Y(n854) );
  MUX2X1 U690 ( .B(b[14]), .A(b[13]), .S(n1187), .Y(n675) );
  MUX2X1 U691 ( .B(n1189), .A(n851), .S(n676), .Y(n855) );
  MUX2X1 U692 ( .B(b[13]), .A(n1223), .S(n1187), .Y(n676) );
  MUX2X1 U693 ( .B(n1189), .A(n851), .S(n677), .Y(n856) );
  MUX2X1 U694 ( .B(n1224), .A(b[11]), .S(n1187), .Y(n677) );
  MUX2X1 U695 ( .B(n1189), .A(n851), .S(n678), .Y(n857) );
  MUX2X1 U696 ( .B(b[11]), .A(n1220), .S(n1187), .Y(n678) );
  MUX2X1 U697 ( .B(n1189), .A(n851), .S(n679), .Y(n858) );
  MUX2X1 U698 ( .B(n1221), .A(n1217), .S(n1187), .Y(n679) );
  MUX2X1 U699 ( .B(n1189), .A(n851), .S(n680), .Y(n859) );
  MUX2X1 U700 ( .B(n1218), .A(b[8]), .S(n1187), .Y(n680) );
  MUX2X1 U701 ( .B(n1188), .A(n851), .S(n681), .Y(n860) );
  MUX2X1 U702 ( .B(b[8]), .A(b[7]), .S(n1186), .Y(n681) );
  MUX2X1 U703 ( .B(n1188), .A(n851), .S(n682), .Y(n861) );
  MUX2X1 U704 ( .B(b[7]), .A(b[6]), .S(n1186), .Y(n682) );
  MUX2X1 U705 ( .B(n1188), .A(n851), .S(n683), .Y(n862) );
  MUX2X1 U706 ( .B(b[6]), .A(b[5]), .S(n1186), .Y(n683) );
  MUX2X1 U707 ( .B(n1188), .A(n851), .S(n684), .Y(n863) );
  MUX2X1 U708 ( .B(b[5]), .A(b[4]), .S(n1186), .Y(n684) );
  MUX2X1 U709 ( .B(n1188), .A(n851), .S(n685), .Y(n864) );
  MUX2X1 U710 ( .B(b[4]), .A(b[3]), .S(n1186), .Y(n685) );
  MUX2X1 U711 ( .B(n1188), .A(n851), .S(n686), .Y(n865) );
  MUX2X1 U712 ( .B(b[3]), .A(n1215), .S(n1186), .Y(n686) );
  MUX2X1 U713 ( .B(n1188), .A(n851), .S(n687), .Y(n866) );
  MUX2X1 U714 ( .B(n1215), .A(n1212), .S(n1186), .Y(n687) );
  MUX2X1 U715 ( .B(n1188), .A(n851), .S(n688), .Y(n867) );
  MUX2X1 U716 ( .B(n1213), .A(n1210), .S(n1186), .Y(n688) );
  MUX2X1 U717 ( .B(n1188), .A(n851), .S(n690), .Y(n868) );
  MUX2X1 U723 ( .B(n1185), .A(n9), .S(n1121), .Y(n870) );
  MUX2X1 U725 ( .B(n1185), .A(n9), .S(n693), .Y(n871) );
  MUX2X1 U726 ( .B(b[15]), .A(b[14]), .S(n1183), .Y(n693) );
  MUX2X1 U727 ( .B(n1185), .A(n9), .S(n694), .Y(n872) );
  MUX2X1 U728 ( .B(b[14]), .A(b[13]), .S(n1183), .Y(n694) );
  MUX2X1 U729 ( .B(n1185), .A(n9), .S(n695), .Y(n873) );
  MUX2X1 U730 ( .B(b[13]), .A(n1223), .S(n1183), .Y(n695) );
  MUX2X1 U731 ( .B(n1185), .A(n9), .S(n696), .Y(n874) );
  MUX2X1 U732 ( .B(n1224), .A(b[11]), .S(n1183), .Y(n696) );
  MUX2X1 U733 ( .B(n1185), .A(n9), .S(n697), .Y(n875) );
  MUX2X1 U734 ( .B(b[11]), .A(n1220), .S(n1183), .Y(n697) );
  MUX2X1 U735 ( .B(n1185), .A(n9), .S(n698), .Y(n876) );
  MUX2X1 U736 ( .B(n1221), .A(n1217), .S(n1183), .Y(n698) );
  MUX2X1 U737 ( .B(n1185), .A(n9), .S(n699), .Y(n877) );
  MUX2X1 U738 ( .B(n1218), .A(b[8]), .S(n1183), .Y(n699) );
  MUX2X1 U739 ( .B(n1184), .A(n9), .S(n700), .Y(n878) );
  MUX2X1 U740 ( .B(b[8]), .A(b[7]), .S(n1182), .Y(n700) );
  MUX2X1 U741 ( .B(n1184), .A(n9), .S(n701), .Y(n879) );
  MUX2X1 U742 ( .B(b[7]), .A(b[6]), .S(n1182), .Y(n701) );
  MUX2X1 U743 ( .B(n1184), .A(n9), .S(n702), .Y(n880) );
  MUX2X1 U744 ( .B(b[6]), .A(b[5]), .S(n1182), .Y(n702) );
  MUX2X1 U745 ( .B(n1184), .A(n9), .S(n703), .Y(n881) );
  MUX2X1 U746 ( .B(b[5]), .A(b[4]), .S(n1182), .Y(n703) );
  MUX2X1 U747 ( .B(n1184), .A(n9), .S(n704), .Y(n882) );
  MUX2X1 U748 ( .B(b[4]), .A(n998), .S(n1182), .Y(n704) );
  MUX2X1 U749 ( .B(n1184), .A(n9), .S(n705), .Y(n883) );
  MUX2X1 U750 ( .B(b[3]), .A(n1215), .S(n1182), .Y(n705) );
  MUX2X1 U751 ( .B(n1184), .A(n9), .S(n706), .Y(n884) );
  MUX2X1 U752 ( .B(n1215), .A(n1212), .S(n1182), .Y(n706) );
  MUX2X1 U753 ( .B(n1184), .A(n9), .S(n707), .Y(n885) );
  MUX2X1 U754 ( .B(n1213), .A(n1210), .S(n1182), .Y(n707) );
  MUX2X1 U755 ( .B(n1184), .A(n9), .S(n709), .Y(n886) );
  AND2X1 U758 ( .A(n1124), .B(a[1]), .Y(n750) );
  MUX2X1 U763 ( .B(n1124), .A(n1228), .S(n712), .Y(n888) );
  MUX2X1 U764 ( .B(b[15]), .A(b[14]), .S(n1226), .Y(n712) );
  MUX2X1 U765 ( .B(n1124), .A(n1228), .S(n713), .Y(n889) );
  MUX2X1 U766 ( .B(b[14]), .A(b[13]), .S(n1226), .Y(n713) );
  MUX2X1 U767 ( .B(n1181), .A(n1228), .S(n714), .Y(n890) );
  MUX2X1 U768 ( .B(b[13]), .A(n1223), .S(n1226), .Y(n714) );
  MUX2X1 U769 ( .B(n1124), .A(n1228), .S(n715), .Y(n891) );
  MUX2X1 U770 ( .B(n1224), .A(b[11]), .S(n1226), .Y(n715) );
  MUX2X1 U771 ( .B(n1124), .A(n1228), .S(n716), .Y(n892) );
  MUX2X1 U772 ( .B(b[11]), .A(n1220), .S(n1226), .Y(n716) );
  MUX2X1 U773 ( .B(n1124), .A(n1228), .S(n717), .Y(n893) );
  MUX2X1 U774 ( .B(n1221), .A(n1217), .S(n1226), .Y(n717) );
  MUX2X1 U775 ( .B(n1181), .A(n1228), .S(n718), .Y(n894) );
  MUX2X1 U776 ( .B(n1218), .A(b[8]), .S(n1226), .Y(n718) );
  MUX2X1 U777 ( .B(n1181), .A(n1228), .S(n719), .Y(n895) );
  MUX2X1 U778 ( .B(b[8]), .A(b[7]), .S(n1226), .Y(n719) );
  MUX2X1 U779 ( .B(n1181), .A(n1228), .S(n720), .Y(n896) );
  MUX2X1 U780 ( .B(b[7]), .A(b[6]), .S(n1226), .Y(n720) );
  MUX2X1 U781 ( .B(n1181), .A(n1228), .S(n721), .Y(n897) );
  MUX2X1 U782 ( .B(b[6]), .A(b[5]), .S(n1227), .Y(n721) );
  MUX2X1 U783 ( .B(n1181), .A(n1228), .S(n722), .Y(n898) );
  MUX2X1 U784 ( .B(b[5]), .A(b[4]), .S(n1227), .Y(n722) );
  MUX2X1 U785 ( .B(n1181), .A(n1228), .S(n723), .Y(n899) );
  MUX2X1 U786 ( .B(b[4]), .A(b[3]), .S(n1227), .Y(n723) );
  MUX2X1 U787 ( .B(n1181), .A(n1228), .S(n724), .Y(n900) );
  MUX2X1 U788 ( .B(b[3]), .A(n1215), .S(n1226), .Y(n724) );
  MUX2X1 U789 ( .B(n1181), .A(n1228), .S(n725), .Y(n901) );
  MUX2X1 U790 ( .B(n1215), .A(n1212), .S(n1226), .Y(n725) );
  MUX2X1 U791 ( .B(n1181), .A(n1228), .S(n726), .Y(n902) );
  MUX2X1 U792 ( .B(n1213), .A(n1210), .S(n1226), .Y(n726) );
  MUX2X1 U793 ( .B(n1181), .A(n1228), .S(n728), .Y(n903) );
  OAI21X1 U798 ( .A(a[13]), .B(a[14]), .C(n1240), .Y(n44) );
  XNOR2X1 U801 ( .A(a[14]), .B(a[13]), .Y(n48) );
  OAI21X1 U803 ( .A(a[12]), .B(a[11]), .C(n1014), .Y(n38) );
  XNOR2X1 U806 ( .A(a[11]), .B(a[12]), .Y(n42) );
  OAI21X1 U808 ( .A(n1011), .B(a[9]), .C(n1233), .Y(n32) );
  OAI21X1 U813 ( .A(a[8]), .B(a[7]), .C(n1232), .Y(n26) );
  XNOR2X1 U816 ( .A(a[7]), .B(a[8]), .Y(n30) );
  OAI21X1 U818 ( .A(a[5]), .B(a[6]), .C(n1231), .Y(n20) );
  XNOR2X1 U821 ( .A(a[6]), .B(a[5]), .Y(n24) );
  OAI21X1 U823 ( .A(a[4]), .B(a[3]), .C(n1230), .Y(n14) );
  XNOR2X1 U826 ( .A(a[3]), .B(a[4]), .Y(n18) );
  OAI21X1 U828 ( .A(a[2]), .B(a[1]), .C(n1229), .Y(n8) );
  XNOR2X1 U831 ( .A(a[1]), .B(a[2]), .Y(n12) );
  BUFX4 U838 ( .A(n24), .Y(n1190) );
  INVX2 U839 ( .A(n1237), .Y(n1236) );
  BUFX2 U840 ( .A(b[3]), .Y(n998) );
  INVX2 U841 ( .A(n1225), .Y(n1224) );
  MUX2X1 U842 ( .B(n1228), .A(n1124), .S(n711), .Y(n887) );
  INVX4 U843 ( .A(n741), .Y(n9) );
  OAI21X1 U844 ( .A(n1016), .B(n1023), .C(n1030), .Y(n999) );
  INVX2 U845 ( .A(n226), .Y(n1016) );
  INVX4 U846 ( .A(n1225), .Y(n1223) );
  BUFX2 U847 ( .A(n177), .Y(n1000) );
  INVX4 U848 ( .A(n1214), .Y(n1212) );
  BUFX4 U849 ( .A(n24), .Y(n1191) );
  INVX8 U850 ( .A(n737), .Y(n833) );
  INVX4 U851 ( .A(n729), .Y(n761) );
  BUFX4 U852 ( .A(n18), .Y(n1187) );
  INVX4 U853 ( .A(n739), .Y(n851) );
  INVX4 U854 ( .A(n1199), .Y(n1001) );
  INVX1 U855 ( .A(n1001), .Y(n1002) );
  INVX8 U856 ( .A(n1001), .Y(n1003) );
  BUFX4 U857 ( .A(n42), .Y(n1203) );
  BUFX4 U858 ( .A(n36), .Y(n1198) );
  OR2X1 U859 ( .A(n1227), .B(n1211), .Y(n728) );
  INVX1 U860 ( .A(a[11]), .Y(n1233) );
  INVX1 U861 ( .A(b[10]), .Y(n1222) );
  INVX2 U862 ( .A(n1222), .Y(n1220) );
  INVX2 U863 ( .A(n731), .Y(n779) );
  INVX2 U864 ( .A(n1235), .Y(n1239) );
  INVX1 U865 ( .A(b[2]), .Y(n1216) );
  INVX1 U866 ( .A(a[0]), .Y(n1226) );
  INVX1 U867 ( .A(n205), .Y(n1162) );
  OR2X1 U868 ( .A(n1183), .B(n1211), .Y(n709) );
  OR2X1 U869 ( .A(n559), .B(n886), .Y(n1171) );
  AND2X1 U870 ( .A(n886), .B(n559), .Y(n258) );
  AND2X1 U871 ( .A(n1164), .B(n261), .Y(product[0]) );
  AND2X1 U872 ( .A(b[15]), .B(n1194), .Y(n635) );
  AND2X1 U873 ( .A(b[15]), .B(n1227), .Y(n711) );
  OR2X1 U874 ( .A(n576), .B(n1239), .Y(n760) );
  OR2X1 U875 ( .A(n1239), .B(n1211), .Y(n576) );
  OR2X1 U876 ( .A(n568), .B(n1239), .Y(n755) );
  OR2X1 U877 ( .A(n570), .B(n1239), .Y(n756) );
  AND2X1 U878 ( .A(b[15]), .B(n1187), .Y(n673) );
  INVX1 U879 ( .A(n759), .Y(n1077) );
  OR2X1 U880 ( .A(n574), .B(n1239), .Y(n759) );
  INVX1 U881 ( .A(n758), .Y(n1154) );
  OR2X1 U882 ( .A(n573), .B(n1240), .Y(n758) );
  BUFX2 U883 ( .A(n36), .Y(n1199) );
  BUFX2 U884 ( .A(n30), .Y(n1195) );
  OR2X1 U885 ( .A(n572), .B(n1240), .Y(n757) );
  OR2X1 U886 ( .A(n1003), .B(n1211), .Y(n633) );
  AND2X1 U887 ( .A(n1201), .B(n733), .Y(n745) );
  OR2X1 U888 ( .A(n566), .B(n1239), .Y(n754) );
  OR2X1 U889 ( .A(n1207), .B(n1211), .Y(n595) );
  OR2X1 U890 ( .A(n1203), .B(n1211), .Y(n614) );
  BUFX2 U891 ( .A(n30), .Y(n1194) );
  OR2X1 U892 ( .A(n1194), .B(n1211), .Y(n652) );
  INVX2 U893 ( .A(n735), .Y(n815) );
  AND2X1 U894 ( .A(n1236), .B(n1234), .Y(n1247) );
  OR2X1 U895 ( .A(n564), .B(n1239), .Y(n753) );
  OR2X1 U896 ( .A(n1088), .B(n1158), .Y(n157) );
  OR2X1 U897 ( .A(n364), .B(n375), .Y(n159) );
  AND2X1 U898 ( .A(n375), .B(n1006), .Y(n160) );
  OR2X1 U899 ( .A(n420), .B(n434), .Y(n182) );
  AND2X1 U900 ( .A(n434), .B(n420), .Y(n183) );
  OR2X1 U901 ( .A(n435), .B(n448), .Y(n185) );
  AND2X1 U902 ( .A(n462), .B(n449), .Y(n191) );
  AND2X1 U903 ( .A(n1172), .B(n1174), .Y(n226) );
  AND2X1 U904 ( .A(a[5]), .B(n1229), .Y(n1242) );
  OR2X1 U905 ( .A(n1191), .B(n1211), .Y(n671) );
  AND2X1 U906 ( .A(a[0]), .B(n1228), .Y(n2) );
  OR2X1 U907 ( .A(n562), .B(n1239), .Y(n752) );
  OR2X1 U908 ( .A(n560), .B(n1239), .Y(n751) );
  AND2X1 U909 ( .A(n1107), .B(n1169), .Y(n90) );
  OR2X1 U910 ( .A(n1055), .B(n1056), .Y(n141) );
  AND2X1 U911 ( .A(n1115), .B(n159), .Y(n94) );
  OR2X1 U912 ( .A(n1117), .B(n1161), .Y(n169) );
  AND2X1 U913 ( .A(n1099), .B(n171), .Y(n96) );
  INVX1 U914 ( .A(n175), .Y(n1139) );
  AND2X1 U915 ( .A(n419), .B(n404), .Y(n175) );
  OR2X1 U916 ( .A(n1156), .B(n1128), .Y(n1029) );
  AND2X1 U917 ( .A(n448), .B(n435), .Y(n186) );
  AND2X1 U918 ( .A(n1114), .B(n190), .Y(n100) );
  AND2X1 U919 ( .A(n1173), .B(n1175), .Y(n208) );
  OR2X1 U920 ( .A(n1187), .B(n1211), .Y(n690) );
  BUFX2 U921 ( .A(n18), .Y(n1186) );
  AND2X1 U922 ( .A(n1193), .B(n737), .Y(n747) );
  INVX2 U923 ( .A(n1211), .Y(n1210) );
  AND2X1 U924 ( .A(n389), .B(n376), .Y(n165) );
  AND2X1 U925 ( .A(n476), .B(n463), .Y(n196) );
  AND2X1 U926 ( .A(n488), .B(n477), .Y(n202) );
  AND2X1 U927 ( .A(n1162), .B(n204), .Y(n103) );
  OR2X1 U928 ( .A(n553), .B(n556), .Y(n1180) );
  AND2X1 U929 ( .A(n1185), .B(n741), .Y(n749) );
  AND2X1 U930 ( .A(n750), .B(n903), .Y(n262) );
  AND2X1 U931 ( .A(n1106), .B(n1176), .Y(n86) );
  OR2X1 U932 ( .A(n463), .B(n476), .Y(n195) );
  AND2X1 U933 ( .A(n1110), .B(n1174), .Y(n107) );
  AND2X1 U934 ( .A(n1147), .B(n1172), .Y(n108) );
  OR2X1 U935 ( .A(n1164), .B(n260), .Y(n259) );
  AND2X1 U936 ( .A(n1108), .B(n1179), .Y(n109) );
  AND2X1 U937 ( .A(n1087), .B(n1171), .Y(n113) );
  BUFX2 U938 ( .A(n129), .Y(n1004) );
  INVX1 U939 ( .A(n364), .Y(n1005) );
  INVX1 U940 ( .A(n1005), .Y(n1006) );
  INVX4 U941 ( .A(n733), .Y(n797) );
  INVX1 U942 ( .A(a[7]), .Y(n1231) );
  INVX1 U943 ( .A(a[3]), .Y(n1229) );
  AND2X1 U944 ( .A(n542), .B(n537), .Y(n236) );
  AND2X1 U945 ( .A(n520), .B(n511), .Y(n218) );
  OR2X1 U946 ( .A(n561), .B(n1239), .Y(n297) );
  OR2X1 U947 ( .A(n376), .B(n389), .Y(n164) );
  INVX1 U948 ( .A(a[9]), .Y(n1232) );
  AND2X1 U949 ( .A(n556), .B(n553), .Y(n250) );
  AND2X1 U950 ( .A(n548), .B(n543), .Y(n242) );
  AND2X1 U951 ( .A(n510), .B(n501), .Y(n213) );
  OR2X1 U952 ( .A(n477), .B(n488), .Y(n201) );
  OR2X1 U953 ( .A(n489), .B(n500), .Y(n204) );
  AND2X1 U954 ( .A(n536), .B(n529), .Y(n231) );
  OR2X1 U955 ( .A(n903), .B(n750), .Y(n261) );
  INVX1 U956 ( .A(a[5]), .Y(n1230) );
  INVX1 U957 ( .A(b[1]), .Y(n1214) );
  INVX1 U958 ( .A(a[0]), .Y(n1227) );
  INVX1 U959 ( .A(b[0]), .Y(n1211) );
  OAI21X1 U960 ( .A(n1149), .B(n1025), .C(n1130), .Y(n1007) );
  INVX4 U961 ( .A(b[12]), .Y(n1225) );
  INVX1 U962 ( .A(b[9]), .Y(n1219) );
  OAI21X1 U963 ( .A(n1153), .B(n1116), .C(n1133), .Y(n1008) );
  BUFX2 U964 ( .A(n259), .Y(n1009) );
  BUFX4 U965 ( .A(n48), .Y(n1207) );
  INVX1 U966 ( .A(a[10]), .Y(n1010) );
  INVX1 U967 ( .A(n1010), .Y(n1011) );
  INVX1 U968 ( .A(n259), .Y(n1012) );
  XNOR2X1 U969 ( .A(n115), .B(n1013), .Y(product[31]) );
  XNOR2X1 U970 ( .A(n295), .B(n294), .Y(n1013) );
  INVX1 U971 ( .A(a[13]), .Y(n1014) );
  INVX1 U972 ( .A(n262), .Y(n1164) );
  OR2X2 U973 ( .A(n543), .B(n548), .Y(n1179) );
  BUFX4 U974 ( .A(n42), .Y(n1202) );
  BUFX2 U975 ( .A(n1066), .Y(n1015) );
  INVX1 U976 ( .A(n1065), .Y(n1066) );
  INVX8 U977 ( .A(n1219), .Y(n1217) );
  BUFX4 U978 ( .A(n48), .Y(n1206) );
  OR2X2 U979 ( .A(n537), .B(n542), .Y(n1172) );
  OR2X2 U980 ( .A(n529), .B(n536), .Y(n1174) );
  INVX8 U981 ( .A(n1236), .Y(n1238) );
  INVX8 U982 ( .A(n1216), .Y(n1215) );
  INVX8 U983 ( .A(a[1]), .Y(n1228) );
  INVX1 U984 ( .A(n208), .Y(n1017) );
  INVX1 U985 ( .A(n169), .Y(n1018) );
  AND2X2 U986 ( .A(n1054), .B(n1018), .Y(n155) );
  BUFX2 U987 ( .A(n179), .Y(n1019) );
  INVX1 U988 ( .A(n141), .Y(n1020) );
  AND2X2 U989 ( .A(n1052), .B(n1027), .Y(n178) );
  INVX1 U990 ( .A(n178), .Y(n1021) );
  BUFX2 U991 ( .A(n156), .Y(n1022) );
  BUFX2 U992 ( .A(n238), .Y(n1023) );
  BUFX2 U993 ( .A(n198), .Y(n1024) );
  BUFX2 U994 ( .A(n124), .Y(n1025) );
  BUFX2 U995 ( .A(n220), .Y(n1026) );
  BUFX4 U996 ( .A(n12), .Y(n1182) );
  OR2X2 U997 ( .A(n1157), .B(n1137), .Y(n180) );
  INVX1 U998 ( .A(n180), .Y(n1027) );
  INVX1 U999 ( .A(n180), .Y(n1028) );
  BUFX2 U1000 ( .A(n227), .Y(n1030) );
  BUFX2 U1001 ( .A(n209), .Y(n1031) );
  BUFX2 U1002 ( .A(n144), .Y(n1032) );
  OR2X1 U1003 ( .A(n1119), .B(n1136), .Y(n199) );
  INVX1 U1004 ( .A(n199), .Y(n1033) );
  AND2X1 U1005 ( .A(b[15]), .B(n1207), .Y(n578) );
  INVX1 U1006 ( .A(n578), .Y(n1034) );
  AND2X1 U1007 ( .A(n1113), .B(n1180), .Y(n111) );
  INVX1 U1008 ( .A(n111), .Y(n1035) );
  BUFX2 U1009 ( .A(n232), .Y(n1036) );
  BUFX2 U1010 ( .A(n214), .Y(n1037) );
  BUFX2 U1011 ( .A(n149), .Y(n1038) );
  AND2X1 U1012 ( .A(n1132), .B(n244), .Y(n110) );
  INVX1 U1013 ( .A(n110), .Y(n1039) );
  INVX1 U1014 ( .A(n108), .Y(n1040) );
  AND2X1 U1015 ( .A(n1126), .B(n1177), .Y(n106) );
  INVX1 U1016 ( .A(n106), .Y(n1041) );
  AND2X1 U1017 ( .A(n1100), .B(n195), .Y(n101) );
  INVX1 U1018 ( .A(n101), .Y(n1042) );
  AND2X1 U1019 ( .A(n1098), .B(n276), .Y(n98) );
  INVX1 U1020 ( .A(n98), .Y(n1043) );
  AND2X1 U1021 ( .A(n1135), .B(n273), .Y(n95) );
  INVX1 U1022 ( .A(n95), .Y(n1044) );
  AND2X1 U1023 ( .A(n1127), .B(n1168), .Y(n93) );
  INVX1 U1024 ( .A(n93), .Y(n1045) );
  INVX1 U1025 ( .A(n107), .Y(n1046) );
  AND2X1 U1026 ( .A(n1111), .B(n1175), .Y(n104) );
  INVX1 U1027 ( .A(n104), .Y(n1047) );
  AND2X1 U1028 ( .A(n1067), .B(n277), .Y(n99) );
  INVX1 U1029 ( .A(n99), .Y(n1048) );
  AND2X1 U1030 ( .A(n1112), .B(n1167), .Y(n92) );
  INVX1 U1031 ( .A(n92), .Y(n1049) );
  AND2X1 U1032 ( .A(n1131), .B(n138), .Y(n91) );
  INVX1 U1033 ( .A(n91), .Y(n1050) );
  AND2X1 U1034 ( .A(n1130), .B(n122), .Y(n87) );
  INVX1 U1035 ( .A(n87), .Y(n1051) );
  INVX1 U1036 ( .A(n1029), .Y(n1052) );
  INVX1 U1037 ( .A(n1029), .Y(n1053) );
  INVX1 U1038 ( .A(n157), .Y(n1054) );
  INVX1 U1039 ( .A(n155), .Y(n1055) );
  AND2X1 U1040 ( .A(n1167), .B(n1168), .Y(n143) );
  INVX1 U1041 ( .A(n143), .Y(n1056) );
  BUFX2 U1042 ( .A(n187), .Y(n1057) );
  INVX1 U1043 ( .A(n140), .Y(n1058) );
  INVX1 U1044 ( .A(n1058), .Y(n1059) );
  INVX1 U1045 ( .A(n1058), .Y(n1060) );
  INVX1 U1046 ( .A(n132), .Y(n1061) );
  INVX1 U1047 ( .A(n1061), .Y(n1062) );
  INVX1 U1048 ( .A(n1061), .Y(n1063) );
  BUFX2 U1049 ( .A(n1025), .Y(n1064) );
  INVX1 U1050 ( .A(n246), .Y(n1065) );
  INVX1 U1051 ( .A(n186), .Y(n1067) );
  INVX1 U1052 ( .A(n1247), .Y(n1068) );
  INVX1 U1053 ( .A(n751), .Y(n1069) );
  INVX1 U1054 ( .A(n752), .Y(n1070) );
  INVX1 U1055 ( .A(n754), .Y(n1071) );
  INVX1 U1056 ( .A(n753), .Y(n1072) );
  AND2X2 U1057 ( .A(a[3]), .B(n1228), .Y(n1241) );
  INVX1 U1058 ( .A(n1241), .Y(n1073) );
  INVX1 U1059 ( .A(n755), .Y(n1074) );
  INVX1 U1060 ( .A(n757), .Y(n1075) );
  INVX1 U1061 ( .A(n756), .Y(n1076) );
  INVX1 U1062 ( .A(n760), .Y(n1078) );
  AND2X2 U1063 ( .A(a[13]), .B(n1233), .Y(n1246) );
  INVX1 U1064 ( .A(n1246), .Y(n1079) );
  INVX1 U1065 ( .A(n94), .Y(n1080) );
  BUFX2 U1066 ( .A(n161), .Y(n1081) );
  INVX1 U1067 ( .A(n297), .Y(n1082) );
  AND2X1 U1068 ( .A(a[11]), .B(n1232), .Y(n1245) );
  INVX1 U1069 ( .A(n1245), .Y(n1083) );
  INVX1 U1070 ( .A(n96), .Y(n1084) );
  INVX1 U1071 ( .A(n100), .Y(n1085) );
  BUFX2 U1072 ( .A(n192), .Y(n1086) );
  INVX1 U1073 ( .A(n258), .Y(n1087) );
  INVX1 U1074 ( .A(n164), .Y(n1088) );
  INVX1 U1075 ( .A(n202), .Y(n1089) );
  OR2X1 U1076 ( .A(n563), .B(n1239), .Y(n307) );
  INVX1 U1077 ( .A(n307), .Y(n1090) );
  INVX1 U1078 ( .A(n1242), .Y(n1091) );
  INVX1 U1079 ( .A(n113), .Y(n1092) );
  AND2X1 U1080 ( .A(n1133), .B(n252), .Y(n112) );
  INVX1 U1081 ( .A(n112), .Y(n1093) );
  AND2X2 U1082 ( .A(n1089), .B(n201), .Y(n102) );
  INVX1 U1083 ( .A(n102), .Y(n1094) );
  AND2X1 U1084 ( .A(n1109), .B(n1170), .Y(n88) );
  INVX1 U1085 ( .A(n88), .Y(n1095) );
  AND2X1 U1086 ( .A(n1129), .B(n130), .Y(n89) );
  INVX1 U1087 ( .A(n89), .Y(n1096) );
  AND2X1 U1088 ( .A(n1139), .B(n275), .Y(n97) );
  INVX1 U1089 ( .A(n97), .Y(n1097) );
  INVX1 U1090 ( .A(n183), .Y(n1098) );
  AND2X2 U1091 ( .A(n403), .B(n390), .Y(n172) );
  INVX1 U1092 ( .A(n172), .Y(n1099) );
  INVX1 U1093 ( .A(n196), .Y(n1100) );
  OR2X1 U1094 ( .A(n565), .B(n1239), .Y(n321) );
  INVX1 U1095 ( .A(n321), .Y(n1101) );
  AND2X2 U1096 ( .A(a[7]), .B(n1230), .Y(n1243) );
  INVX1 U1097 ( .A(n1243), .Y(n1102) );
  AND2X1 U1098 ( .A(b[15]), .B(n1203), .Y(n597) );
  INVX1 U1099 ( .A(n597), .Y(n1103) );
  AND2X1 U1100 ( .A(b[15]), .B(n1003), .Y(n616) );
  INVX1 U1101 ( .A(n616), .Y(n1104) );
  INVX1 U1102 ( .A(n103), .Y(n1105) );
  AND2X1 U1103 ( .A(n300), .B(n303), .Y(n120) );
  INVX1 U1104 ( .A(n120), .Y(n1106) );
  AND2X1 U1105 ( .A(n324), .B(n331), .Y(n136) );
  INVX1 U1106 ( .A(n136), .Y(n1107) );
  INVX1 U1107 ( .A(n242), .Y(n1108) );
  AND2X1 U1108 ( .A(n310), .B(n315), .Y(n128) );
  INVX1 U1109 ( .A(n128), .Y(n1109) );
  INVX1 U1110 ( .A(n231), .Y(n1110) );
  INVX1 U1111 ( .A(n213), .Y(n1111) );
  AND2X1 U1112 ( .A(n342), .B(n351), .Y(n148) );
  INVX1 U1113 ( .A(n148), .Y(n1112) );
  INVX1 U1114 ( .A(n250), .Y(n1113) );
  INVX1 U1115 ( .A(n191), .Y(n1114) );
  INVX1 U1116 ( .A(n160), .Y(n1115) );
  BUFX2 U1117 ( .A(n254), .Y(n1116) );
  OR2X2 U1118 ( .A(n404), .B(n419), .Y(n174) );
  INVX1 U1119 ( .A(n174), .Y(n1117) );
  INVX1 U1120 ( .A(n174), .Y(n1118) );
  INVX1 U1121 ( .A(n201), .Y(n1119) );
  OR2X1 U1122 ( .A(n567), .B(n1239), .Y(n339) );
  INVX1 U1123 ( .A(n339), .Y(n1120) );
  AND2X2 U1124 ( .A(b[15]), .B(n1183), .Y(n692) );
  INVX1 U1125 ( .A(n692), .Y(n1121) );
  BUFX4 U1126 ( .A(n12), .Y(n1183) );
  AND2X1 U1127 ( .A(b[15]), .B(n1190), .Y(n654) );
  INVX1 U1128 ( .A(n654), .Y(n1122) );
  AND2X1 U1129 ( .A(n1148), .B(n1173), .Y(n105) );
  INVX1 U1130 ( .A(n105), .Y(n1123) );
  INVX1 U1131 ( .A(n2), .Y(n1124) );
  INVX1 U1132 ( .A(n2), .Y(n1125) );
  AND2X1 U1133 ( .A(n528), .B(n521), .Y(n224) );
  INVX1 U1134 ( .A(n224), .Y(n1126) );
  AND2X1 U1135 ( .A(n363), .B(n352), .Y(n153) );
  INVX1 U1136 ( .A(n153), .Y(n1127) );
  INVX1 U1137 ( .A(n195), .Y(n1128) );
  AND2X1 U1138 ( .A(n316), .B(n323), .Y(n131) );
  INVX1 U1139 ( .A(n131), .Y(n1129) );
  AND2X1 U1140 ( .A(n304), .B(n309), .Y(n123) );
  INVX1 U1141 ( .A(n123), .Y(n1130) );
  AND2X1 U1142 ( .A(n332), .B(n341), .Y(n139) );
  INVX1 U1143 ( .A(n139), .Y(n1131) );
  AND2X1 U1144 ( .A(n552), .B(n549), .Y(n245) );
  INVX1 U1145 ( .A(n245), .Y(n1132) );
  AND2X1 U1146 ( .A(n558), .B(n557), .Y(n253) );
  INVX1 U1147 ( .A(n253), .Y(n1133) );
  INVX1 U1148 ( .A(n1009), .Y(n1134) );
  INVX1 U1149 ( .A(n165), .Y(n1135) );
  INVX1 U1150 ( .A(n204), .Y(n1136) );
  INVX1 U1151 ( .A(n185), .Y(n1137) );
  INVX1 U1152 ( .A(n185), .Y(n1138) );
  OR2X1 U1153 ( .A(n571), .B(n1239), .Y(n387) );
  INVX1 U1154 ( .A(n387), .Y(n1140) );
  AND2X1 U1155 ( .A(a[9]), .B(n1231), .Y(n1244) );
  INVX1 U1156 ( .A(n1244), .Y(n1141) );
  INVX1 U1157 ( .A(n635), .Y(n1142) );
  INVX1 U1158 ( .A(n673), .Y(n1143) );
  INVX1 U1159 ( .A(n109), .Y(n1144) );
  INVX1 U1160 ( .A(n90), .Y(n1145) );
  INVX1 U1161 ( .A(n86), .Y(n1146) );
  INVX1 U1162 ( .A(n236), .Y(n1147) );
  INVX1 U1163 ( .A(n218), .Y(n1148) );
  OR2X1 U1164 ( .A(n309), .B(n304), .Y(n122) );
  INVX1 U1165 ( .A(n122), .Y(n1149) );
  OR2X1 U1166 ( .A(n323), .B(n316), .Y(n130) );
  INVX1 U1167 ( .A(n130), .Y(n1150) );
  OR2X1 U1168 ( .A(n341), .B(n332), .Y(n138) );
  INVX1 U1169 ( .A(n138), .Y(n1151) );
  OR2X1 U1170 ( .A(n549), .B(n552), .Y(n244) );
  INVX1 U1171 ( .A(n244), .Y(n1152) );
  OR2X1 U1172 ( .A(n557), .B(n558), .Y(n252) );
  INVX1 U1173 ( .A(n252), .Y(n1153) );
  OR2X2 U1174 ( .A(n449), .B(n462), .Y(n190) );
  INVX1 U1175 ( .A(n190), .Y(n1155) );
  INVX1 U1176 ( .A(n190), .Y(n1156) );
  INVX1 U1177 ( .A(n182), .Y(n1157) );
  INVX1 U1178 ( .A(n159), .Y(n1158) );
  INVX1 U1179 ( .A(n159), .Y(n1159) );
  OR2X2 U1180 ( .A(n390), .B(n403), .Y(n171) );
  INVX1 U1181 ( .A(n171), .Y(n1160) );
  INVX1 U1182 ( .A(n171), .Y(n1161) );
  AND2X1 U1183 ( .A(n500), .B(n489), .Y(n205) );
  OR2X1 U1184 ( .A(n569), .B(n1239), .Y(n361) );
  INVX1 U1185 ( .A(n361), .Y(n1163) );
  BUFX2 U1186 ( .A(n137), .Y(n1165) );
  BUFX2 U1187 ( .A(n243), .Y(n1166) );
  INVX1 U1188 ( .A(n1138), .Y(n277) );
  INVX1 U1189 ( .A(n1118), .Y(n275) );
  INVX1 U1190 ( .A(n1157), .Y(n276) );
  INVX1 U1191 ( .A(n207), .Y(n206) );
  INVX1 U1192 ( .A(n1024), .Y(n197) );
  INVX1 U1193 ( .A(n1135), .Y(n163) );
  INVX1 U1194 ( .A(n1026), .Y(n219) );
  INVX1 U1195 ( .A(n1088), .Y(n273) );
  INVX1 U1196 ( .A(n1236), .Y(n1240) );
  BUFX2 U1197 ( .A(n20), .Y(n1192) );
  BUFX2 U1198 ( .A(n20), .Y(n1193) );
  INVX1 U1199 ( .A(n1237), .Y(n1235) );
  INVX1 U1200 ( .A(n1023), .Y(n237) );
  OR2X1 U1201 ( .A(n351), .B(n342), .Y(n1167) );
  OR2X1 U1202 ( .A(n352), .B(n363), .Y(n1168) );
  OR2X1 U1203 ( .A(n331), .B(n324), .Y(n1169) );
  OR2X1 U1204 ( .A(n315), .B(n310), .Y(n1170) );
  BUFX2 U1205 ( .A(n44), .Y(n1208) );
  BUFX2 U1206 ( .A(n32), .Y(n1200) );
  BUFX2 U1207 ( .A(n8), .Y(n1184) );
  BUFX2 U1208 ( .A(n26), .Y(n1196) );
  BUFX2 U1209 ( .A(n44), .Y(n1209) );
  BUFX2 U1210 ( .A(n32), .Y(n1201) );
  BUFX2 U1211 ( .A(n8), .Y(n1185) );
  BUFX2 U1212 ( .A(n26), .Y(n1197) );
  INVX1 U1213 ( .A(n116), .Y(n263) );
  INVX1 U1214 ( .A(n902), .Y(n260) );
  INVX1 U1215 ( .A(a[15]), .Y(n1237) );
  OR2X1 U1216 ( .A(n511), .B(n520), .Y(n1173) );
  OR2X1 U1217 ( .A(n501), .B(n510), .Y(n1175) );
  OR2X1 U1218 ( .A(n303), .B(n300), .Y(n1176) );
  OR2X1 U1219 ( .A(n521), .B(n528), .Y(n1177) );
  INVX1 U1220 ( .A(n1222), .Y(n1221) );
  INVX1 U1221 ( .A(n1219), .Y(n1218) );
  INVX1 U1222 ( .A(n1214), .Y(n1213) );
  BUFX2 U1223 ( .A(n38), .Y(n1204) );
  BUFX2 U1224 ( .A(n38), .Y(n1205) );
  BUFX2 U1225 ( .A(n14), .Y(n1188) );
  BUFX2 U1226 ( .A(n14), .Y(n1189) );
  INVX1 U1227 ( .A(a[13]), .Y(n1234) );
  XOR2X1 U1228 ( .A(n1232), .B(a[10]), .Y(n36) );
  INVX1 U1229 ( .A(n170), .Y(n168) );
  INVX1 U1230 ( .A(n1000), .Y(n176) );
  BUFX2 U1231 ( .A(n1125), .Y(n1181) );
  OAI21X1 U1232 ( .A(a[2]), .B(n1229), .C(n1073), .Y(n741) );
  OAI21X1 U1233 ( .A(a[4]), .B(n1230), .C(n1091), .Y(n739) );
  OAI21X1 U1234 ( .A(a[6]), .B(n1231), .C(n1102), .Y(n737) );
  OAI21X1 U1235 ( .A(a[8]), .B(n1232), .C(n1141), .Y(n735) );
  OAI21X1 U1236 ( .A(n1011), .B(n1233), .C(n1083), .Y(n733) );
  OAI21X1 U1237 ( .A(a[12]), .B(n1014), .C(n1079), .Y(n731) );
  OAI21X1 U1238 ( .A(a[14]), .B(n1239), .C(n1068), .Y(n729) );
  XOR2X1 U1239 ( .A(n1069), .B(n1082), .Y(n293) );
endmodule


module alu_DW_mult_uns_38 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n2, n8, n9, n12, n14, n18, n20, n24, n26, n30, n32, n36, n38, n42,
         n44, n48, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n114, n115, n119, n120, n121, n125, n126,
         n127, n128, n129, n133, n134, n135, n136, n137, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n186, n187, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n204, n205, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n226, n227, n231, n232, n233, n237, n238, n239, n240, n241,
         n245, n246, n247, n248, n249, n250, n254, n255, n256, n267, n285,
         n286, n287, n288, n289, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n568, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n587, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n606, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n625, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n644, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n663, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n682,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n701, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n720, n721, n723, n725, n727, n729, n731, n733, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n895, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217;

  XOR2X1 U85 ( .A(n114), .B(n85), .Y(product[31]) );
  XOR2X1 U86 ( .A(n287), .B(n286), .Y(n85) );
  FAX1 U87 ( .A(n288), .B(n291), .C(n255), .YC(n114), .YS(product[30]) );
  XNOR2X1 U89 ( .A(n120), .B(n1091), .Y(product[29]) );
  AOI21X1 U90 ( .A(n120), .B(n1138), .C(n119), .Y(n115) );
  FAX1 U97 ( .A(n296), .B(n301), .C(n256), .YC(n120), .YS(product[28]) );
  XNOR2X1 U99 ( .A(n1128), .B(n1110), .Y(product[27]) );
  AOI21X1 U100 ( .A(n126), .B(n1132), .C(n125), .Y(n121) );
  OAI21X1 U108 ( .A(n1117), .B(n992), .C(n1099), .Y(n126) );
  XNOR2X1 U113 ( .A(n134), .B(n1054), .Y(product[25]) );
  AOI21X1 U114 ( .A(n134), .B(n1131), .C(n133), .Y(n129) );
  XOR2X1 U121 ( .A(n1012), .B(n1074), .Y(product[24]) );
  OAI21X1 U122 ( .A(n1116), .B(n1013), .C(n1098), .Y(n134) );
  XNOR2X1 U127 ( .A(n1147), .B(n1040), .Y(product[23]) );
  AOI21X1 U128 ( .A(n142), .B(n1130), .C(n141), .Y(n137) );
  XOR2X1 U135 ( .A(n1010), .B(n1043), .Y(product[22]) );
  OAI21X1 U136 ( .A(n1100), .B(n1010), .C(n1079), .Y(n142) );
  XNOR2X1 U141 ( .A(n150), .B(n1001), .Y(product[21]) );
  AOI21X1 U142 ( .A(n168), .B(n998), .C(n147), .Y(n145) );
  OAI21X1 U144 ( .A(n1122), .B(n1007), .C(n1063), .Y(n147) );
  XNOR2X1 U149 ( .A(n157), .B(n1053), .Y(product[20]) );
  OAI21X1 U150 ( .A(n1008), .B(n167), .C(n1007), .Y(n150) );
  AOI21X1 U152 ( .A(n161), .B(n1129), .C(n156), .Y(n152) );
  XNOR2X1 U159 ( .A(n164), .B(n1039), .Y(product[19]) );
  OAI21X1 U160 ( .A(n158), .B(n167), .C(n159), .Y(n157) );
  OAI21X1 U164 ( .A(n1126), .B(n1105), .C(n1078), .Y(n161) );
  XOR2X1 U169 ( .A(n167), .B(n1002), .Y(product[18]) );
  OAI21X1 U170 ( .A(n1065), .B(n167), .C(n1126), .Y(n164) );
  XNOR2X1 U175 ( .A(n175), .B(n1024), .Y(product[17]) );
  OAI21X1 U177 ( .A(n1004), .B(n991), .C(n996), .Y(n168) );
  AOI21X1 U179 ( .A(n1005), .B(n180), .C(n172), .Y(n170) );
  OAI21X1 U181 ( .A(n1125), .B(n1085), .C(n1046), .Y(n172) );
  XOR2X1 U186 ( .A(n1064), .B(n1033), .Y(product[16]) );
  OAI21X1 U187 ( .A(n1104), .B(n1064), .C(n1125), .Y(n175) );
  XOR2X1 U192 ( .A(n1032), .B(n1031), .Y(product[15]) );
  AOI21X1 U193 ( .A(n1003), .B(n1050), .C(n180), .Y(n178) );
  OAI21X1 U195 ( .A(n1121), .B(n1084), .C(n1047), .Y(n180) );
  XNOR2X1 U200 ( .A(n1003), .B(n1037), .Y(product[14]) );
  AOI21X1 U201 ( .A(n1003), .B(n186), .C(n187), .Y(n183) );
  XNOR2X1 U208 ( .A(n194), .B(n1038), .Y(product[13]) );
  AOI21X1 U210 ( .A(n198), .B(n997), .C(n191), .Y(n189) );
  OAI21X1 U212 ( .A(n1124), .B(n1083), .C(n1062), .Y(n191) );
  XOR2X1 U217 ( .A(n197), .B(n1073), .Y(product[12]) );
  OAI21X1 U218 ( .A(n1103), .B(n197), .C(n1124), .Y(n194) );
  XOR2X1 U223 ( .A(n1056), .B(n1055), .Y(product[11]) );
  OAI21X1 U225 ( .A(n999), .B(n1048), .C(n994), .Y(n198) );
  AOI21X1 U227 ( .A(n1137), .B(n209), .C(n204), .Y(n200) );
  XNOR2X1 U234 ( .A(n210), .B(n1090), .Y(product[10]) );
  AOI21X1 U235 ( .A(n210), .B(n1134), .C(n209), .Y(n205) );
  XNOR2X1 U242 ( .A(n216), .B(n1030), .Y(product[9]) );
  AOI21X1 U244 ( .A(n1049), .B(n220), .C(n213), .Y(n211) );
  OAI21X1 U246 ( .A(n1123), .B(n1082), .C(n1061), .Y(n213) );
  XOR2X1 U251 ( .A(n219), .B(n1072), .Y(product[8]) );
  OAI21X1 U252 ( .A(n1102), .B(n219), .C(n1123), .Y(n216) );
  XOR2X1 U257 ( .A(n1042), .B(n1041), .Y(product[7]) );
  OAI21X1 U259 ( .A(n1080), .B(n1023), .C(n1022), .Y(n220) );
  AOI21X1 U261 ( .A(n1136), .B(n231), .C(n226), .Y(n222) );
  XNOR2X1 U268 ( .A(n1089), .B(n232), .Y(product[6]) );
  AOI21X1 U269 ( .A(n232), .B(n1135), .C(n231), .Y(n227) );
  XNOR2X1 U276 ( .A(n1029), .B(n238), .Y(product[5]) );
  AOI21X1 U278 ( .A(n238), .B(n1139), .C(n237), .Y(n233) );
  XOR2X1 U285 ( .A(n1070), .B(n1101), .Y(product[4]) );
  OAI21X1 U286 ( .A(n1115), .B(n1101), .C(n1059), .Y(n238) );
  XNOR2X1 U291 ( .A(n1028), .B(n246), .Y(product[3]) );
  AOI21X1 U292 ( .A(n246), .B(n1133), .C(n245), .Y(n241) );
  XOR2X1 U299 ( .A(n1036), .B(n1120), .Y(product[2]) );
  OAI21X1 U300 ( .A(n1120), .B(n1081), .C(n1060), .Y(n246) );
  XOR2X1 U315 ( .A(n753), .B(n285), .Y(n286) );
  FAX1 U317 ( .A(n289), .B(n754), .C(n293), .YC(n287), .YS(n288) );
  FAX1 U319 ( .A(n755), .B(n294), .C(n297), .YC(n291), .YS(n292) );
  FAX1 U320 ( .A(n771), .B(n1051), .C(n1016), .YC(n293), .YS(n294) );
  FAX1 U321 ( .A(n305), .B(n298), .C(n303), .YC(n295), .YS(n296) );
  FAX1 U322 ( .A(n299), .B(n772), .C(n756), .YC(n297), .YS(n298) );
  FAX1 U324 ( .A(n311), .B(n304), .C(n309), .YC(n301), .YS(n302) );
  FAX1 U325 ( .A(n773), .B(n757), .C(n306), .YC(n303), .YS(n304) );
  FAX1 U326 ( .A(n789), .B(n1066), .C(n1018), .YC(n305), .YS(n306) );
  FAX1 U327 ( .A(n319), .B(n310), .C(n317), .YC(n307), .YS(n308) );
  FAX1 U328 ( .A(n758), .B(n321), .C(n312), .YC(n309), .YS(n310) );
  FAX1 U329 ( .A(n313), .B(n790), .C(n774), .YC(n311), .YS(n312) );
  FAX1 U331 ( .A(n320), .B(n318), .C(n325), .YC(n315), .YS(n316) );
  FAX1 U332 ( .A(n322), .B(n329), .C(n327), .YC(n317), .YS(n318) );
  FAX1 U333 ( .A(n775), .B(n791), .C(n759), .YC(n319), .YS(n320) );
  FAX1 U334 ( .A(n807), .B(n1086), .C(n1017), .YC(n321), .YS(n322) );
  FAX1 U335 ( .A(n337), .B(n326), .C(n335), .YC(n323), .YS(n324) );
  FAX1 U336 ( .A(n330), .B(n339), .C(n328), .YC(n325), .YS(n326) );
  FAX1 U337 ( .A(n792), .B(n760), .C(n341), .YC(n327), .YS(n328) );
  FAX1 U338 ( .A(n331), .B(n808), .C(n776), .YC(n329), .YS(n330) );
  FAX1 U340 ( .A(n347), .B(n336), .C(n345), .YC(n333), .YS(n334) );
  FAX1 U341 ( .A(n349), .B(n340), .C(n338), .YC(n335), .YS(n336) );
  FAX1 U342 ( .A(n777), .B(n342), .C(n351), .YC(n337), .YS(n338) );
  FAX1 U343 ( .A(n809), .B(n793), .C(n761), .YC(n339), .YS(n340) );
  FAX1 U344 ( .A(n825), .B(n1106), .C(n1019), .YC(n341), .YS(n342) );
  FAX1 U345 ( .A(n359), .B(n346), .C(n357), .YC(n343), .YS(n344) );
  FAX1 U346 ( .A(n361), .B(n350), .C(n348), .YC(n345), .YS(n346) );
  FAX1 U347 ( .A(n794), .B(n352), .C(n363), .YC(n347), .YS(n348) );
  FAX1 U348 ( .A(n778), .B(n762), .C(n365), .YC(n349), .YS(n350) );
  FAX1 U349 ( .A(n353), .B(n826), .C(n810), .YC(n351), .YS(n352) );
  FAX1 U351 ( .A(n360), .B(n369), .C(n358), .YC(n355), .YS(n356) );
  FAX1 U352 ( .A(n362), .B(n373), .C(n371), .YC(n357), .YS(n358) );
  FAX1 U353 ( .A(n377), .B(n375), .C(n364), .YC(n359), .YS(n360) );
  FAX1 U354 ( .A(n779), .B(n827), .C(n366), .YC(n361), .YS(n362) );
  FAX1 U355 ( .A(n811), .B(n795), .C(n763), .YC(n363), .YS(n364) );
  FAX1 U356 ( .A(n843), .B(n1127), .C(n1020), .YC(n365), .YS(n366) );
  FAX1 U357 ( .A(n372), .B(n383), .C(n370), .YC(n367), .YS(n368) );
  FAX1 U358 ( .A(n374), .B(n387), .C(n385), .YC(n369), .YS(n370) );
  FAX1 U359 ( .A(n389), .B(n391), .C(n376), .YC(n371), .YS(n372) );
  FAX1 U360 ( .A(n828), .B(n796), .C(n378), .YC(n373), .YS(n374) );
  FAX1 U361 ( .A(n780), .B(n764), .C(n393), .YC(n375), .YS(n376) );
  FAX1 U362 ( .A(n379), .B(n844), .C(n812), .YC(n377), .YS(n378) );
  FAX1 U364 ( .A(n386), .B(n397), .C(n384), .YC(n381), .YS(n382) );
  FAX1 U365 ( .A(n401), .B(n388), .C(n399), .YC(n383), .YS(n384) );
  FAX1 U366 ( .A(n403), .B(n392), .C(n390), .YC(n385), .YS(n386) );
  FAX1 U367 ( .A(n781), .B(n407), .C(n405), .YC(n387), .YS(n388) );
  FAX1 U368 ( .A(n845), .B(n829), .C(n797), .YC(n389), .YS(n390) );
  FAX1 U369 ( .A(n813), .B(n765), .C(n394), .YC(n391), .YS(n392) );
  FAX1 U370 ( .A(n1202), .B(n9), .C(n1097), .YC(n393), .YS(n394) );
  FAX1 U371 ( .A(n400), .B(n413), .C(n398), .YC(n395), .YS(n396) );
  FAX1 U372 ( .A(n417), .B(n402), .C(n415), .YC(n397), .YS(n398) );
  FAX1 U373 ( .A(n419), .B(n406), .C(n404), .YC(n399), .YS(n400) );
  FAX1 U374 ( .A(n408), .B(n423), .C(n421), .YC(n401), .YS(n402) );
  FAX1 U375 ( .A(n846), .B(n782), .C(n830), .YC(n403), .YS(n404) );
  FAX1 U376 ( .A(n814), .B(n798), .C(n766), .YC(n405), .YS(n406) );
  FAX1 U377 ( .A(n1199), .B(n1118), .C(n862), .YC(n407), .YS(n408) );
  FAX1 U379 ( .A(n416), .B(n428), .C(n414), .YC(n411), .YS(n412) );
  FAX1 U380 ( .A(n432), .B(n418), .C(n430), .YC(n413), .YS(n414) );
  FAX1 U381 ( .A(n436), .B(n422), .C(n420), .YC(n415), .YS(n416) );
  FAX1 U382 ( .A(n438), .B(n424), .C(n434), .YC(n417), .YS(n418) );
  FAX1 U383 ( .A(n847), .B(n783), .C(n831), .YC(n419), .YS(n420) );
  FAX1 U384 ( .A(n815), .B(n799), .C(n767), .YC(n421), .YS(n422) );
  FAX1 U385 ( .A(n1199), .B(n1025), .C(n863), .YC(n423), .YS(n424) );
  FAX1 U387 ( .A(n431), .B(n442), .C(n429), .YC(n426), .YS(n427) );
  FAX1 U388 ( .A(n446), .B(n433), .C(n1095), .YC(n428), .YS(n429) );
  FAX1 U389 ( .A(n448), .B(n437), .C(n435), .YC(n430), .YS(n431) );
  FAX1 U390 ( .A(n452), .B(n439), .C(n450), .YC(n432), .YS(n433) );
  FAX1 U391 ( .A(n848), .B(n784), .C(n832), .YC(n434), .YS(n435) );
  FAX1 U392 ( .A(n816), .B(n800), .C(n768), .YC(n436), .YS(n437) );
  FAX1 U393 ( .A(n879), .B(n1021), .C(n864), .YC(n438), .YS(n439) );
  FAX1 U394 ( .A(n445), .B(n456), .C(n443), .YC(n440), .YS(n441) );
  FAX1 U395 ( .A(n460), .B(n447), .C(n458), .YC(n442), .YS(n443) );
  FAX1 U397 ( .A(n785), .B(n453), .C(n464), .YC(n446), .YS(n447) );
  FAX1 U398 ( .A(n849), .B(n833), .C(n801), .YC(n448), .YS(n449) );
  FAX1 U399 ( .A(n817), .B(n769), .C(n466), .YC(n450), .YS(n451) );
  HAX1 U400 ( .A(n880), .B(n865), .YC(n452), .YS(n453) );
  FAX1 U401 ( .A(n459), .B(n470), .C(n457), .YC(n454), .YS(n455) );
  FAX1 U402 ( .A(n474), .B(n461), .C(n472), .YC(n456), .YS(n457) );
  FAX1 U403 ( .A(n476), .B(n465), .C(n463), .YC(n458), .YS(n459) );
  FAX1 U404 ( .A(n818), .B(n850), .C(n478), .YC(n460), .YS(n461) );
  FAX1 U405 ( .A(n866), .B(n786), .C(n467), .YC(n462), .YS(n463) );
  FAX1 U406 ( .A(n770), .B(n834), .C(n802), .YC(n464), .YS(n465) );
  HAX1 U407 ( .A(n881), .B(n735), .YC(n466), .YS(n467) );
  FAX1 U408 ( .A(n473), .B(n482), .C(n471), .YC(n468), .YS(n469) );
  FAX1 U409 ( .A(n477), .B(n475), .C(n484), .YC(n470), .YS(n471) );
  FAX1 U410 ( .A(n479), .B(n488), .C(n486), .YC(n472), .YS(n473) );
  FAX1 U411 ( .A(n851), .B(n787), .C(n835), .YC(n474), .YS(n475) );
  FAX1 U412 ( .A(n819), .B(n803), .C(n490), .YC(n476), .YS(n477) );
  HAX1 U413 ( .A(n882), .B(n867), .YC(n478), .YS(n479) );
  FAX1 U414 ( .A(n485), .B(n494), .C(n483), .YC(n480), .YS(n481) );
  FAX1 U415 ( .A(n489), .B(n487), .C(n496), .YC(n482), .YS(n483) );
  FAX1 U416 ( .A(n820), .B(n500), .C(n498), .YC(n484), .YS(n485) );
  FAX1 U417 ( .A(n868), .B(n852), .C(n491), .YC(n486), .YS(n487) );
  FAX1 U418 ( .A(n788), .B(n836), .C(n804), .YC(n488), .YS(n489) );
  HAX1 U419 ( .A(n883), .B(n736), .YC(n490), .YS(n491) );
  FAX1 U420 ( .A(n497), .B(n504), .C(n495), .YC(n492), .YS(n493) );
  FAX1 U421 ( .A(n508), .B(n506), .C(n499), .YC(n494), .YS(n495) );
  FAX1 U422 ( .A(n853), .B(n837), .C(n501), .YC(n496), .YS(n497) );
  FAX1 U423 ( .A(n821), .B(n805), .C(n510), .YC(n498), .YS(n499) );
  HAX1 U424 ( .A(n884), .B(n869), .YC(n500), .YS(n501) );
  FAX1 U425 ( .A(n507), .B(n514), .C(n505), .YC(n502), .YS(n503) );
  FAX1 U426 ( .A(n518), .B(n516), .C(n509), .YC(n504), .YS(n505) );
  FAX1 U427 ( .A(n870), .B(n822), .C(n511), .YC(n506), .YS(n507) );
  FAX1 U428 ( .A(n806), .B(n854), .C(n838), .YC(n508), .YS(n509) );
  HAX1 U429 ( .A(n885), .B(n737), .YC(n510), .YS(n511) );
  FAX1 U430 ( .A(n517), .B(n522), .C(n515), .YC(n512), .YS(n513) );
  FAX1 U431 ( .A(n855), .B(n519), .C(n524), .YC(n514), .YS(n515) );
  FAX1 U432 ( .A(n823), .B(n839), .C(n526), .YC(n516), .YS(n517) );
  HAX1 U433 ( .A(n886), .B(n871), .YC(n518), .YS(n519) );
  FAX1 U434 ( .A(n530), .B(n525), .C(n523), .YC(n520), .YS(n521) );
  FAX1 U435 ( .A(n872), .B(n527), .C(n532), .YC(n522), .YS(n523) );
  FAX1 U436 ( .A(n824), .B(n856), .C(n840), .YC(n524), .YS(n525) );
  HAX1 U437 ( .A(n887), .B(n738), .YC(n526), .YS(n527) );
  FAX1 U438 ( .A(n533), .B(n536), .C(n531), .YC(n528), .YS(n529) );
  FAX1 U439 ( .A(n857), .B(n841), .C(n538), .YC(n530), .YS(n531) );
  HAX1 U440 ( .A(n888), .B(n873), .YC(n532), .YS(n533) );
  FAX1 U441 ( .A(n539), .B(n542), .C(n537), .YC(n534), .YS(n535) );
  FAX1 U442 ( .A(n842), .B(n874), .C(n858), .YC(n536), .YS(n537) );
  HAX1 U443 ( .A(n889), .B(n739), .YC(n538), .YS(n539) );
  FAX1 U444 ( .A(n859), .B(n546), .C(n543), .YC(n540), .YS(n541) );
  HAX1 U445 ( .A(n890), .B(n875), .YC(n542), .YS(n543) );
  FAX1 U446 ( .A(n860), .B(n876), .C(n547), .YC(n544), .YS(n545) );
  HAX1 U447 ( .A(n891), .B(n740), .YC(n546), .YS(n547) );
  HAX1 U448 ( .A(n892), .B(n877), .YC(n548), .YS(n549) );
  HAX1 U449 ( .A(n893), .B(n741), .YC(n550), .YS(n551) );
  MUX2X1 U451 ( .B(b[15]), .A(b[14]), .S(n1210), .Y(n552) );
  MUX2X1 U453 ( .B(b[14]), .A(b[13]), .S(n1210), .Y(n553) );
  MUX2X1 U455 ( .B(b[13]), .A(b[12]), .S(n1210), .Y(n554) );
  MUX2X1 U457 ( .B(b[12]), .A(n1195), .S(n1210), .Y(n555) );
  MUX2X1 U459 ( .B(n1195), .A(b[10]), .S(n1210), .Y(n556) );
  MUX2X1 U461 ( .B(b[10]), .A(b[9]), .S(n1210), .Y(n557) );
  MUX2X1 U463 ( .B(b[9]), .A(b[8]), .S(n1210), .Y(n558) );
  MUX2X1 U465 ( .B(b[8]), .A(b[7]), .S(n1210), .Y(n559) );
  MUX2X1 U467 ( .B(b[7]), .A(n1193), .S(n1210), .Y(n560) );
  MUX2X1 U469 ( .B(n1193), .A(n1190), .S(n1210), .Y(n561) );
  MUX2X1 U471 ( .B(n1190), .A(n1188), .S(n1210), .Y(n562) );
  MUX2X1 U473 ( .B(n1188), .A(n1185), .S(n1210), .Y(n563) );
  MUX2X1 U475 ( .B(n1185), .A(n1183), .S(n1210), .Y(n564) );
  MUX2X1 U477 ( .B(n1183), .A(n1180), .S(n1210), .Y(n565) );
  MUX2X1 U479 ( .B(n1180), .A(n1178), .S(n1210), .Y(n566) );
  MUX2X1 U486 ( .B(n1177), .A(n753), .S(n1000), .Y(n754) );
  MUX2X1 U488 ( .B(n1177), .A(n753), .S(n571), .Y(n755) );
  MUX2X1 U489 ( .B(b[15]), .A(b[14]), .S(n1175), .Y(n571) );
  MUX2X1 U490 ( .B(n1177), .A(n753), .S(n572), .Y(n756) );
  MUX2X1 U491 ( .B(b[14]), .A(b[13]), .S(n1175), .Y(n572) );
  MUX2X1 U492 ( .B(n1177), .A(n753), .S(n573), .Y(n757) );
  MUX2X1 U493 ( .B(b[13]), .A(b[12]), .S(n1175), .Y(n573) );
  MUX2X1 U494 ( .B(n1177), .A(n753), .S(n574), .Y(n758) );
  MUX2X1 U495 ( .B(b[12]), .A(n1195), .S(n1175), .Y(n574) );
  MUX2X1 U496 ( .B(n1177), .A(n753), .S(n575), .Y(n759) );
  MUX2X1 U497 ( .B(n1195), .A(b[10]), .S(n1175), .Y(n575) );
  MUX2X1 U498 ( .B(n1177), .A(n753), .S(n576), .Y(n760) );
  MUX2X1 U499 ( .B(b[10]), .A(b[9]), .S(n1175), .Y(n576) );
  MUX2X1 U500 ( .B(n1177), .A(n753), .S(n577), .Y(n761) );
  MUX2X1 U501 ( .B(b[9]), .A(b[8]), .S(n1175), .Y(n577) );
  MUX2X1 U502 ( .B(n1176), .A(n753), .S(n578), .Y(n762) );
  MUX2X1 U503 ( .B(b[8]), .A(b[7]), .S(n1174), .Y(n578) );
  MUX2X1 U504 ( .B(n1176), .A(n753), .S(n579), .Y(n763) );
  MUX2X1 U505 ( .B(b[7]), .A(n1193), .S(n1174), .Y(n579) );
  MUX2X1 U506 ( .B(n1176), .A(n753), .S(n580), .Y(n764) );
  MUX2X1 U507 ( .B(n1193), .A(n1190), .S(n1174), .Y(n580) );
  MUX2X1 U508 ( .B(n1176), .A(n753), .S(n581), .Y(n765) );
  MUX2X1 U509 ( .B(n1190), .A(n1188), .S(n1174), .Y(n581) );
  MUX2X1 U510 ( .B(n1176), .A(n753), .S(n582), .Y(n766) );
  MUX2X1 U511 ( .B(n1188), .A(n1185), .S(n1174), .Y(n582) );
  MUX2X1 U512 ( .B(n1176), .A(n753), .S(n583), .Y(n767) );
  MUX2X1 U513 ( .B(n1185), .A(n1183), .S(n1174), .Y(n583) );
  MUX2X1 U514 ( .B(n1176), .A(n753), .S(n584), .Y(n768) );
  MUX2X1 U515 ( .B(n1183), .A(n1180), .S(n1174), .Y(n584) );
  MUX2X1 U516 ( .B(n1176), .A(n753), .S(n585), .Y(n769) );
  MUX2X1 U517 ( .B(n1180), .A(n1178), .S(n1174), .Y(n585) );
  MUX2X1 U518 ( .B(n1176), .A(n753), .S(n587), .Y(n770) );
  OR2X1 U519 ( .A(n1175), .B(n1179), .Y(n587) );
  AND2X1 U521 ( .A(n1173), .B(n723), .Y(n736) );
  MUX2X1 U524 ( .B(n1173), .A(n771), .S(n1068), .Y(n772) );
  MUX2X1 U526 ( .B(n1173), .A(n771), .S(n590), .Y(n773) );
  MUX2X1 U527 ( .B(b[15]), .A(b[14]), .S(n1171), .Y(n590) );
  MUX2X1 U528 ( .B(n1173), .A(n771), .S(n591), .Y(n774) );
  MUX2X1 U529 ( .B(b[14]), .A(b[13]), .S(n1171), .Y(n591) );
  MUX2X1 U530 ( .B(n1173), .A(n771), .S(n592), .Y(n775) );
  MUX2X1 U531 ( .B(b[13]), .A(b[12]), .S(n1171), .Y(n592) );
  MUX2X1 U532 ( .B(n1173), .A(n771), .S(n593), .Y(n776) );
  MUX2X1 U533 ( .B(b[12]), .A(n1195), .S(n1171), .Y(n593) );
  MUX2X1 U534 ( .B(n1173), .A(n771), .S(n594), .Y(n777) );
  MUX2X1 U535 ( .B(n1196), .A(b[10]), .S(n1171), .Y(n594) );
  MUX2X1 U536 ( .B(n1173), .A(n771), .S(n595), .Y(n778) );
  MUX2X1 U537 ( .B(b[10]), .A(b[9]), .S(n1171), .Y(n595) );
  MUX2X1 U538 ( .B(n1173), .A(n771), .S(n596), .Y(n779) );
  MUX2X1 U539 ( .B(b[9]), .A(b[8]), .S(n1171), .Y(n596) );
  MUX2X1 U540 ( .B(n1172), .A(n771), .S(n597), .Y(n780) );
  MUX2X1 U541 ( .B(b[8]), .A(b[7]), .S(n1170), .Y(n597) );
  MUX2X1 U542 ( .B(n1172), .A(n771), .S(n598), .Y(n781) );
  MUX2X1 U543 ( .B(b[7]), .A(n1193), .S(n1170), .Y(n598) );
  MUX2X1 U544 ( .B(n1172), .A(n771), .S(n599), .Y(n782) );
  MUX2X1 U545 ( .B(b[6]), .A(n1190), .S(n1170), .Y(n599) );
  MUX2X1 U546 ( .B(n1172), .A(n771), .S(n600), .Y(n783) );
  MUX2X1 U547 ( .B(n1191), .A(n1188), .S(n1170), .Y(n600) );
  MUX2X1 U548 ( .B(n1172), .A(n771), .S(n601), .Y(n784) );
  MUX2X1 U549 ( .B(b[4]), .A(n1185), .S(n1170), .Y(n601) );
  MUX2X1 U550 ( .B(n1172), .A(n771), .S(n602), .Y(n785) );
  MUX2X1 U551 ( .B(n1186), .A(n1183), .S(n1170), .Y(n602) );
  MUX2X1 U552 ( .B(n1172), .A(n771), .S(n603), .Y(n786) );
  MUX2X1 U553 ( .B(b[2]), .A(n1180), .S(n1170), .Y(n603) );
  MUX2X1 U554 ( .B(n1172), .A(n771), .S(n604), .Y(n787) );
  MUX2X1 U555 ( .B(n1181), .A(n1178), .S(n1170), .Y(n604) );
  MUX2X1 U556 ( .B(n1172), .A(n771), .S(n606), .Y(n788) );
  OR2X1 U557 ( .A(n1171), .B(n1179), .Y(n606) );
  AND2X1 U559 ( .A(n1169), .B(n725), .Y(n737) );
  MUX2X1 U562 ( .B(n1169), .A(n789), .S(n1069), .Y(n790) );
  MUX2X1 U564 ( .B(n1169), .A(n789), .S(n609), .Y(n791) );
  MUX2X1 U565 ( .B(b[15]), .A(b[14]), .S(n1167), .Y(n609) );
  MUX2X1 U566 ( .B(n1169), .A(n789), .S(n610), .Y(n792) );
  MUX2X1 U567 ( .B(b[14]), .A(b[13]), .S(n1167), .Y(n610) );
  MUX2X1 U568 ( .B(n1169), .A(n789), .S(n611), .Y(n793) );
  MUX2X1 U569 ( .B(b[13]), .A(b[12]), .S(n1167), .Y(n611) );
  MUX2X1 U570 ( .B(n1169), .A(n789), .S(n612), .Y(n794) );
  MUX2X1 U571 ( .B(b[12]), .A(n1195), .S(n1167), .Y(n612) );
  MUX2X1 U572 ( .B(n1169), .A(n789), .S(n613), .Y(n795) );
  MUX2X1 U573 ( .B(n1196), .A(b[10]), .S(n1167), .Y(n613) );
  MUX2X1 U574 ( .B(n1169), .A(n789), .S(n614), .Y(n796) );
  MUX2X1 U575 ( .B(b[10]), .A(b[9]), .S(n1167), .Y(n614) );
  MUX2X1 U576 ( .B(n1169), .A(n789), .S(n615), .Y(n797) );
  MUX2X1 U577 ( .B(b[9]), .A(b[8]), .S(n1167), .Y(n615) );
  MUX2X1 U578 ( .B(n1168), .A(n789), .S(n616), .Y(n798) );
  MUX2X1 U579 ( .B(b[8]), .A(b[7]), .S(n1166), .Y(n616) );
  MUX2X1 U580 ( .B(n1168), .A(n789), .S(n617), .Y(n799) );
  MUX2X1 U581 ( .B(b[7]), .A(n1193), .S(n1166), .Y(n617) );
  MUX2X1 U582 ( .B(n1168), .A(n789), .S(n618), .Y(n800) );
  MUX2X1 U583 ( .B(b[6]), .A(n1190), .S(n1166), .Y(n618) );
  MUX2X1 U584 ( .B(n1168), .A(n789), .S(n619), .Y(n801) );
  MUX2X1 U585 ( .B(n1191), .A(n1188), .S(n1166), .Y(n619) );
  MUX2X1 U586 ( .B(n1168), .A(n789), .S(n620), .Y(n802) );
  MUX2X1 U587 ( .B(b[4]), .A(n1185), .S(n1166), .Y(n620) );
  MUX2X1 U588 ( .B(n1168), .A(n789), .S(n621), .Y(n803) );
  MUX2X1 U589 ( .B(n1186), .A(n1183), .S(n1166), .Y(n621) );
  MUX2X1 U590 ( .B(n1168), .A(n789), .S(n622), .Y(n804) );
  MUX2X1 U591 ( .B(b[2]), .A(n1180), .S(n1166), .Y(n622) );
  MUX2X1 U592 ( .B(n1168), .A(n789), .S(n623), .Y(n805) );
  MUX2X1 U593 ( .B(n1181), .A(n1178), .S(n1166), .Y(n623) );
  MUX2X1 U594 ( .B(n1168), .A(n789), .S(n625), .Y(n806) );
  OR2X1 U595 ( .A(n1167), .B(n1179), .Y(n625) );
  AND2X1 U597 ( .A(n1165), .B(n727), .Y(n738) );
  MUX2X1 U600 ( .B(n1165), .A(n807), .S(n1052), .Y(n808) );
  MUX2X1 U602 ( .B(n1165), .A(n807), .S(n628), .Y(n809) );
  MUX2X1 U603 ( .B(b[15]), .A(b[14]), .S(n1163), .Y(n628) );
  MUX2X1 U604 ( .B(n1165), .A(n807), .S(n629), .Y(n810) );
  MUX2X1 U605 ( .B(b[14]), .A(b[13]), .S(n1163), .Y(n629) );
  MUX2X1 U606 ( .B(n1165), .A(n807), .S(n630), .Y(n811) );
  MUX2X1 U607 ( .B(b[13]), .A(b[12]), .S(n1163), .Y(n630) );
  MUX2X1 U608 ( .B(n1165), .A(n807), .S(n631), .Y(n812) );
  MUX2X1 U609 ( .B(b[12]), .A(n1195), .S(n1163), .Y(n631) );
  MUX2X1 U610 ( .B(n1165), .A(n807), .S(n632), .Y(n813) );
  MUX2X1 U611 ( .B(n1195), .A(b[10]), .S(n1163), .Y(n632) );
  MUX2X1 U612 ( .B(n1165), .A(n807), .S(n633), .Y(n814) );
  MUX2X1 U613 ( .B(b[10]), .A(b[9]), .S(n1163), .Y(n633) );
  MUX2X1 U614 ( .B(n1165), .A(n807), .S(n634), .Y(n815) );
  MUX2X1 U615 ( .B(b[9]), .A(b[8]), .S(n1163), .Y(n634) );
  MUX2X1 U616 ( .B(n1164), .A(n807), .S(n635), .Y(n816) );
  MUX2X1 U617 ( .B(b[8]), .A(b[7]), .S(n1162), .Y(n635) );
  MUX2X1 U618 ( .B(n1164), .A(n807), .S(n636), .Y(n817) );
  MUX2X1 U619 ( .B(b[7]), .A(n1193), .S(n1162), .Y(n636) );
  MUX2X1 U620 ( .B(n1164), .A(n807), .S(n637), .Y(n818) );
  MUX2X1 U621 ( .B(n1193), .A(n1190), .S(n1162), .Y(n637) );
  MUX2X1 U622 ( .B(n1164), .A(n807), .S(n638), .Y(n819) );
  MUX2X1 U623 ( .B(n1190), .A(n1188), .S(n1162), .Y(n638) );
  MUX2X1 U624 ( .B(n1164), .A(n807), .S(n639), .Y(n820) );
  MUX2X1 U625 ( .B(n1188), .A(n1185), .S(n1162), .Y(n639) );
  MUX2X1 U626 ( .B(n1164), .A(n807), .S(n640), .Y(n821) );
  MUX2X1 U627 ( .B(n1185), .A(n1183), .S(n1162), .Y(n640) );
  MUX2X1 U628 ( .B(n1164), .A(n807), .S(n641), .Y(n822) );
  MUX2X1 U629 ( .B(n1183), .A(n1180), .S(n1162), .Y(n641) );
  MUX2X1 U630 ( .B(n1164), .A(n807), .S(n642), .Y(n823) );
  MUX2X1 U631 ( .B(n1180), .A(n1178), .S(n1162), .Y(n642) );
  MUX2X1 U632 ( .B(n1164), .A(n807), .S(n644), .Y(n824) );
  OR2X1 U633 ( .A(n1163), .B(n1179), .Y(n644) );
  AND2X1 U635 ( .A(n1161), .B(n729), .Y(n739) );
  MUX2X1 U638 ( .B(n1161), .A(n825), .S(n1109), .Y(n826) );
  MUX2X1 U640 ( .B(n1161), .A(n825), .S(n647), .Y(n827) );
  MUX2X1 U641 ( .B(b[15]), .A(b[14]), .S(n1159), .Y(n647) );
  MUX2X1 U642 ( .B(n1161), .A(n825), .S(n648), .Y(n828) );
  MUX2X1 U643 ( .B(b[14]), .A(b[13]), .S(n1159), .Y(n648) );
  MUX2X1 U644 ( .B(n1161), .A(n825), .S(n649), .Y(n829) );
  MUX2X1 U645 ( .B(b[13]), .A(b[12]), .S(n1159), .Y(n649) );
  MUX2X1 U646 ( .B(n1161), .A(n825), .S(n650), .Y(n830) );
  MUX2X1 U647 ( .B(b[12]), .A(n1195), .S(n1159), .Y(n650) );
  MUX2X1 U648 ( .B(n1161), .A(n825), .S(n651), .Y(n831) );
  MUX2X1 U649 ( .B(n1195), .A(b[10]), .S(n1159), .Y(n651) );
  MUX2X1 U650 ( .B(n1161), .A(n825), .S(n652), .Y(n832) );
  MUX2X1 U651 ( .B(b[10]), .A(b[9]), .S(n1159), .Y(n652) );
  MUX2X1 U652 ( .B(n1161), .A(n825), .S(n653), .Y(n833) );
  MUX2X1 U653 ( .B(b[9]), .A(b[8]), .S(n1159), .Y(n653) );
  MUX2X1 U654 ( .B(n1160), .A(n825), .S(n654), .Y(n834) );
  MUX2X1 U655 ( .B(b[8]), .A(b[7]), .S(n1158), .Y(n654) );
  MUX2X1 U656 ( .B(n1160), .A(n825), .S(n655), .Y(n835) );
  MUX2X1 U657 ( .B(b[7]), .A(n1193), .S(n1158), .Y(n655) );
  MUX2X1 U658 ( .B(n1160), .A(n825), .S(n656), .Y(n836) );
  MUX2X1 U659 ( .B(n1193), .A(n1190), .S(n1158), .Y(n656) );
  MUX2X1 U660 ( .B(n1160), .A(n825), .S(n657), .Y(n837) );
  MUX2X1 U661 ( .B(n1190), .A(n1188), .S(n1158), .Y(n657) );
  MUX2X1 U662 ( .B(n1160), .A(n825), .S(n658), .Y(n838) );
  MUX2X1 U663 ( .B(n1188), .A(n1185), .S(n1158), .Y(n658) );
  MUX2X1 U664 ( .B(n1160), .A(n825), .S(n659), .Y(n839) );
  MUX2X1 U665 ( .B(n1185), .A(n1183), .S(n1158), .Y(n659) );
  MUX2X1 U666 ( .B(n1160), .A(n825), .S(n660), .Y(n840) );
  MUX2X1 U667 ( .B(n1183), .A(n1180), .S(n1158), .Y(n660) );
  MUX2X1 U668 ( .B(n1160), .A(n825), .S(n661), .Y(n841) );
  MUX2X1 U669 ( .B(n1180), .A(n1178), .S(n1158), .Y(n661) );
  MUX2X1 U670 ( .B(n1160), .A(n825), .S(n663), .Y(n842) );
  OR2X1 U671 ( .A(n1159), .B(n1179), .Y(n663) );
  AND2X1 U673 ( .A(n1157), .B(n731), .Y(n740) );
  MUX2X1 U676 ( .B(n1157), .A(n843), .S(n1088), .Y(n844) );
  MUX2X1 U678 ( .B(n1157), .A(n843), .S(n666), .Y(n845) );
  MUX2X1 U679 ( .B(b[15]), .A(b[14]), .S(n1155), .Y(n666) );
  MUX2X1 U680 ( .B(n1157), .A(n843), .S(n667), .Y(n846) );
  MUX2X1 U681 ( .B(b[14]), .A(b[13]), .S(n1155), .Y(n667) );
  MUX2X1 U682 ( .B(n1157), .A(n843), .S(n668), .Y(n847) );
  MUX2X1 U683 ( .B(b[13]), .A(b[12]), .S(n1155), .Y(n668) );
  MUX2X1 U684 ( .B(n1157), .A(n843), .S(n669), .Y(n848) );
  MUX2X1 U685 ( .B(b[12]), .A(n1195), .S(n1155), .Y(n669) );
  MUX2X1 U686 ( .B(n1157), .A(n843), .S(n670), .Y(n849) );
  MUX2X1 U687 ( .B(n1196), .A(b[10]), .S(n1155), .Y(n670) );
  MUX2X1 U688 ( .B(n1157), .A(n843), .S(n671), .Y(n850) );
  MUX2X1 U689 ( .B(b[10]), .A(b[9]), .S(n1155), .Y(n671) );
  MUX2X1 U690 ( .B(n1157), .A(n843), .S(n672), .Y(n851) );
  MUX2X1 U691 ( .B(b[9]), .A(b[8]), .S(n1155), .Y(n672) );
  MUX2X1 U692 ( .B(n1156), .A(n843), .S(n673), .Y(n852) );
  MUX2X1 U693 ( .B(b[8]), .A(b[7]), .S(n1154), .Y(n673) );
  MUX2X1 U694 ( .B(n1156), .A(n843), .S(n674), .Y(n853) );
  MUX2X1 U695 ( .B(b[7]), .A(n1193), .S(n1154), .Y(n674) );
  MUX2X1 U696 ( .B(n1156), .A(n843), .S(n675), .Y(n854) );
  MUX2X1 U697 ( .B(b[6]), .A(n1190), .S(n1154), .Y(n675) );
  MUX2X1 U698 ( .B(n1156), .A(n843), .S(n676), .Y(n855) );
  MUX2X1 U699 ( .B(n1191), .A(n1188), .S(n1154), .Y(n676) );
  MUX2X1 U700 ( .B(n1156), .A(n843), .S(n677), .Y(n856) );
  MUX2X1 U701 ( .B(b[4]), .A(n1185), .S(n1154), .Y(n677) );
  MUX2X1 U702 ( .B(n1156), .A(n843), .S(n678), .Y(n857) );
  MUX2X1 U703 ( .B(n1186), .A(n1183), .S(n1154), .Y(n678) );
  MUX2X1 U704 ( .B(n1156), .A(n843), .S(n679), .Y(n858) );
  MUX2X1 U705 ( .B(b[2]), .A(n1180), .S(n1154), .Y(n679) );
  MUX2X1 U706 ( .B(n1156), .A(n843), .S(n680), .Y(n859) );
  MUX2X1 U707 ( .B(n1181), .A(n1178), .S(n1154), .Y(n680) );
  MUX2X1 U708 ( .B(n1156), .A(n843), .S(n682), .Y(n860) );
  OR2X1 U709 ( .A(n1155), .B(n1179), .Y(n682) );
  AND2X1 U711 ( .A(n1153), .B(n733), .Y(n741) );
  MUX2X1 U714 ( .B(n1153), .A(n9), .S(n1119), .Y(n862) );
  MUX2X1 U716 ( .B(n1153), .A(n9), .S(n685), .Y(n863) );
  MUX2X1 U717 ( .B(b[15]), .A(b[14]), .S(n1151), .Y(n685) );
  MUX2X1 U718 ( .B(n1153), .A(n9), .S(n686), .Y(n864) );
  MUX2X1 U719 ( .B(b[14]), .A(b[13]), .S(n1151), .Y(n686) );
  MUX2X1 U720 ( .B(n1153), .A(n9), .S(n687), .Y(n865) );
  MUX2X1 U721 ( .B(b[13]), .A(b[12]), .S(n1151), .Y(n687) );
  MUX2X1 U722 ( .B(n1153), .A(n9), .S(n688), .Y(n866) );
  MUX2X1 U723 ( .B(b[12]), .A(n1195), .S(n1151), .Y(n688) );
  MUX2X1 U724 ( .B(n1153), .A(n9), .S(n689), .Y(n867) );
  MUX2X1 U725 ( .B(n1196), .A(b[10]), .S(n1151), .Y(n689) );
  MUX2X1 U726 ( .B(n1153), .A(n9), .S(n690), .Y(n868) );
  MUX2X1 U727 ( .B(b[10]), .A(b[9]), .S(n1151), .Y(n690) );
  MUX2X1 U728 ( .B(n1153), .A(n9), .S(n691), .Y(n869) );
  MUX2X1 U729 ( .B(b[9]), .A(b[8]), .S(n1151), .Y(n691) );
  MUX2X1 U730 ( .B(n1152), .A(n9), .S(n692), .Y(n870) );
  MUX2X1 U731 ( .B(b[8]), .A(b[7]), .S(n1150), .Y(n692) );
  MUX2X1 U732 ( .B(n1152), .A(n9), .S(n693), .Y(n871) );
  MUX2X1 U733 ( .B(b[7]), .A(n1193), .S(n1150), .Y(n693) );
  MUX2X1 U734 ( .B(n1152), .A(n9), .S(n694), .Y(n872) );
  MUX2X1 U735 ( .B(b[6]), .A(n1190), .S(n1150), .Y(n694) );
  MUX2X1 U736 ( .B(n1152), .A(n9), .S(n695), .Y(n873) );
  MUX2X1 U737 ( .B(n1191), .A(n1188), .S(n1150), .Y(n695) );
  MUX2X1 U738 ( .B(n1152), .A(n9), .S(n696), .Y(n874) );
  MUX2X1 U739 ( .B(b[4]), .A(n1185), .S(n1150), .Y(n696) );
  MUX2X1 U740 ( .B(n1152), .A(n9), .S(n697), .Y(n875) );
  MUX2X1 U741 ( .B(n1186), .A(n1183), .S(n1150), .Y(n697) );
  MUX2X1 U742 ( .B(n1152), .A(n9), .S(n698), .Y(n876) );
  MUX2X1 U743 ( .B(b[2]), .A(n1180), .S(n1150), .Y(n698) );
  MUX2X1 U744 ( .B(n1152), .A(n9), .S(n699), .Y(n877) );
  MUX2X1 U745 ( .B(n1181), .A(n1178), .S(n1150), .Y(n699) );
  MUX2X1 U746 ( .B(n1152), .A(n9), .S(n701), .Y(n878) );
  OR2X1 U747 ( .A(n1151), .B(n1179), .Y(n701) );
  AND2X1 U749 ( .A(n1149), .B(n1200), .Y(n742) );
  MUX2X1 U752 ( .B(n1149), .A(n1202), .S(n1087), .Y(n879) );
  MUX2X1 U754 ( .B(n1149), .A(n1202), .S(n704), .Y(n880) );
  MUX2X1 U755 ( .B(b[15]), .A(b[14]), .S(n1198), .Y(n704) );
  MUX2X1 U756 ( .B(n1149), .A(n1202), .S(n705), .Y(n881) );
  MUX2X1 U757 ( .B(b[14]), .A(b[13]), .S(n1198), .Y(n705) );
  MUX2X1 U758 ( .B(n1149), .A(n1202), .S(n706), .Y(n882) );
  MUX2X1 U759 ( .B(b[13]), .A(b[12]), .S(n1198), .Y(n706) );
  MUX2X1 U760 ( .B(n1149), .A(n1202), .S(n707), .Y(n883) );
  MUX2X1 U761 ( .B(b[12]), .A(n1195), .S(n1198), .Y(n707) );
  MUX2X1 U762 ( .B(n1149), .A(n1202), .S(n708), .Y(n884) );
  MUX2X1 U763 ( .B(n1196), .A(b[10]), .S(n1198), .Y(n708) );
  MUX2X1 U764 ( .B(n1149), .A(n1202), .S(n709), .Y(n885) );
  MUX2X1 U765 ( .B(b[10]), .A(b[9]), .S(n1198), .Y(n709) );
  MUX2X1 U766 ( .B(n1149), .A(n1202), .S(n710), .Y(n886) );
  MUX2X1 U767 ( .B(b[9]), .A(b[8]), .S(n1198), .Y(n710) );
  MUX2X1 U768 ( .B(n1148), .A(n1202), .S(n711), .Y(n887) );
  MUX2X1 U769 ( .B(b[8]), .A(b[7]), .S(n1198), .Y(n711) );
  MUX2X1 U770 ( .B(n1148), .A(n1202), .S(n712), .Y(n888) );
  MUX2X1 U771 ( .B(b[7]), .A(n1193), .S(n1198), .Y(n712) );
  MUX2X1 U772 ( .B(n1148), .A(n1202), .S(n713), .Y(n889) );
  MUX2X1 U773 ( .B(b[6]), .A(n1190), .S(n1198), .Y(n713) );
  MUX2X1 U774 ( .B(n1148), .A(n1202), .S(n714), .Y(n890) );
  MUX2X1 U775 ( .B(n1191), .A(n1188), .S(n1198), .Y(n714) );
  MUX2X1 U776 ( .B(n1148), .A(n1202), .S(n715), .Y(n891) );
  MUX2X1 U777 ( .B(b[4]), .A(n1185), .S(n1198), .Y(n715) );
  MUX2X1 U778 ( .B(n1148), .A(n1202), .S(n716), .Y(n892) );
  MUX2X1 U779 ( .B(n1186), .A(n1183), .S(n1198), .Y(n716) );
  MUX2X1 U780 ( .B(n1148), .A(n1202), .S(n717), .Y(n893) );
  MUX2X1 U781 ( .B(b[2]), .A(n1180), .S(n1198), .Y(n717) );
  MUX2X1 U782 ( .B(n1148), .A(n1202), .S(n718), .Y(n250) );
  MUX2X1 U783 ( .B(n1181), .A(n1178), .S(n1198), .Y(n718) );
  MUX2X1 U784 ( .B(n1148), .A(n1202), .S(n720), .Y(n895) );
  OR2X1 U785 ( .A(n1198), .B(n1179), .Y(n720) );
  OAI21X1 U789 ( .A(a[13]), .B(a[14]), .C(n1210), .Y(n44) );
  XNOR2X1 U792 ( .A(a[14]), .B(a[13]), .Y(n48) );
  OAI21X1 U794 ( .A(a[12]), .B(a[11]), .C(n1209), .Y(n38) );
  XNOR2X1 U797 ( .A(a[11]), .B(a[12]), .Y(n42) );
  OAI21X1 U799 ( .A(a[10]), .B(a[9]), .C(n1208), .Y(n32) );
  XNOR2X1 U802 ( .A(a[9]), .B(a[10]), .Y(n36) );
  OAI21X1 U804 ( .A(a[8]), .B(a[7]), .C(n1207), .Y(n26) );
  XNOR2X1 U807 ( .A(a[7]), .B(a[8]), .Y(n30) );
  OAI21X1 U809 ( .A(n1204), .B(a[6]), .C(n1206), .Y(n20) );
  XNOR2X1 U812 ( .A(a[6]), .B(n1204), .Y(n24) );
  OAI21X1 U814 ( .A(a[4]), .B(a[3]), .C(n1205), .Y(n14) );
  XNOR2X1 U817 ( .A(a[3]), .B(a[4]), .Y(n18) );
  OAI21X1 U819 ( .A(a[2]), .B(n1200), .C(n1203), .Y(n8) );
  XNOR2X1 U822 ( .A(n1200), .B(a[2]), .Y(n12) );
  INVX2 U829 ( .A(a[0]), .Y(n1198) );
  AND2X2 U830 ( .A(a[0]), .B(n1202), .Y(n2) );
  INVX8 U831 ( .A(n1199), .Y(n1202) );
  INVX2 U832 ( .A(n725), .Y(n789) );
  INVX8 U833 ( .A(a[15]), .Y(n1210) );
  INVX4 U834 ( .A(n733), .Y(n9) );
  OR2X1 U835 ( .A(n566), .B(n1210), .Y(n751) );
  OR2X1 U836 ( .A(n568), .B(n1210), .Y(n752) );
  OR2X1 U837 ( .A(n1210), .B(n1179), .Y(n568) );
  INVX1 U838 ( .A(a[9]), .Y(n1207) );
  OR2X1 U839 ( .A(n562), .B(n1210), .Y(n748) );
  BUFX2 U840 ( .A(n24), .Y(n1159) );
  INVX1 U841 ( .A(n1205), .Y(n1204) );
  OR2X1 U842 ( .A(n560), .B(n1210), .Y(n747) );
  AND2X1 U843 ( .A(n449), .B(n451), .Y(n1143) );
  AND2X1 U844 ( .A(n1177), .B(n721), .Y(n735) );
  BUFX2 U845 ( .A(n48), .Y(n1174) );
  INVX1 U846 ( .A(n1184), .Y(n1183) );
  OR2X1 U847 ( .A(n558), .B(n1210), .Y(n746) );
  INVX1 U848 ( .A(a[1]), .Y(n1201) );
  OR2X1 U849 ( .A(n554), .B(n1210), .Y(n744) );
  OR2X1 U850 ( .A(n556), .B(n1210), .Y(n745) );
  OR2X1 U851 ( .A(n1082), .B(n1102), .Y(n212) );
  INVX1 U852 ( .A(n1201), .Y(n1199) );
  OR2X1 U853 ( .A(n552), .B(n1210), .Y(n743) );
  AND2X1 U854 ( .A(n411), .B(n396), .Y(n166) );
  OR2X1 U855 ( .A(n1084), .B(n1094), .Y(n179) );
  AND2X1 U856 ( .A(n1075), .B(n1132), .Y(n87) );
  AND2X1 U857 ( .A(n1044), .B(n1129), .Y(n94) );
  AND2X1 U858 ( .A(n1046), .B(n173), .Y(n97) );
  AND2X1 U859 ( .A(n1125), .B(n176), .Y(n98) );
  AND2X1 U860 ( .A(n1059), .B(n239), .Y(n110) );
  AND2X1 U861 ( .A(n1060), .B(n247), .Y(n112) );
  INVX2 U862 ( .A(n1182), .Y(n1180) );
  OR2X1 U863 ( .A(n1085), .B(n1104), .Y(n171) );
  AND2X1 U864 ( .A(n1092), .B(n1140), .Y(product[0]) );
  OR2X1 U865 ( .A(n553), .B(n1210), .Y(n289) );
  OR2X1 U866 ( .A(n559), .B(n1210), .Y(n331) );
  OR2X1 U867 ( .A(n557), .B(n1210), .Y(n313) );
  OR2X1 U868 ( .A(n563), .B(n1210), .Y(n379) );
  OR2X1 U869 ( .A(n561), .B(n1210), .Y(n353) );
  OR2X1 U870 ( .A(n555), .B(n1210), .Y(n299) );
  OR2X1 U871 ( .A(n382), .B(n395), .Y(n162) );
  AND2X1 U872 ( .A(n462), .B(n451), .Y(n1142) );
  AND2X1 U873 ( .A(n449), .B(n462), .Y(n1144) );
  INVX1 U874 ( .A(a[11]), .Y(n1208) );
  OR2X1 U875 ( .A(n396), .B(n411), .Y(n165) );
  OR2X1 U876 ( .A(n412), .B(n426), .Y(n173) );
  OR2X1 U877 ( .A(n427), .B(n440), .Y(n176) );
  OR2X1 U878 ( .A(n1065), .B(n1105), .Y(n160) );
  INVX2 U879 ( .A(n721), .Y(n753) );
  INVX2 U880 ( .A(n731), .Y(n843) );
  INVX2 U881 ( .A(n727), .Y(n807) );
  OR2X2 U882 ( .A(n1008), .B(n1122), .Y(n146) );
  INVX1 U883 ( .A(a[3]), .Y(n1203) );
  INVX1 U884 ( .A(b[6]), .Y(n1194) );
  INVX1 U885 ( .A(a[5]), .Y(n1205) );
  INVX1 U886 ( .A(n171), .Y(n990) );
  AND2X2 U887 ( .A(n1050), .B(n990), .Y(n169) );
  INVX1 U888 ( .A(n169), .Y(n991) );
  BUFX2 U889 ( .A(n129), .Y(n992) );
  INVX1 U890 ( .A(n160), .Y(n993) );
  BUFX2 U891 ( .A(n200), .Y(n994) );
  INVX1 U892 ( .A(n170), .Y(n995) );
  INVX1 U893 ( .A(n995), .Y(n996) );
  OR2X1 U894 ( .A(n1083), .B(n1103), .Y(n190) );
  INVX1 U895 ( .A(n190), .Y(n997) );
  INVX1 U896 ( .A(n146), .Y(n998) );
  AND2X1 U897 ( .A(n1134), .B(n1137), .Y(n199) );
  INVX1 U898 ( .A(n199), .Y(n999) );
  AND2X1 U899 ( .A(b[15]), .B(n1175), .Y(n570) );
  INVX1 U900 ( .A(n570), .Y(n1000) );
  AND2X1 U901 ( .A(n1063), .B(n148), .Y(n93) );
  INVX1 U902 ( .A(n93), .Y(n1001) );
  AND2X1 U903 ( .A(n1126), .B(n267), .Y(n96) );
  INVX1 U904 ( .A(n96), .Y(n1002) );
  INVX1 U905 ( .A(n189), .Y(n1003) );
  INVX1 U906 ( .A(n1003), .Y(n1004) );
  INVX1 U907 ( .A(n171), .Y(n1005) );
  INVX1 U908 ( .A(n152), .Y(n1006) );
  INVX1 U909 ( .A(n1006), .Y(n1007) );
  AND2X2 U910 ( .A(n993), .B(n1129), .Y(n151) );
  INVX1 U911 ( .A(n151), .Y(n1008) );
  INVX1 U912 ( .A(n145), .Y(n1009) );
  INVX1 U913 ( .A(n1009), .Y(n1010) );
  INVX1 U914 ( .A(n137), .Y(n1011) );
  INVX1 U915 ( .A(n1011), .Y(n1012) );
  INVX1 U916 ( .A(n1011), .Y(n1013) );
  AND2X1 U917 ( .A(a[15]), .B(n1209), .Y(n1217) );
  INVX1 U918 ( .A(n1217), .Y(n1014) );
  INVX1 U919 ( .A(n743), .Y(n1015) );
  INVX1 U920 ( .A(n744), .Y(n1016) );
  INVX1 U921 ( .A(n746), .Y(n1017) );
  INVX1 U922 ( .A(n745), .Y(n1018) );
  INVX1 U923 ( .A(n747), .Y(n1019) );
  INVX1 U924 ( .A(n748), .Y(n1020) );
  INVX1 U925 ( .A(n752), .Y(n1021) );
  OR2X2 U926 ( .A(n1142), .B(n1096), .Y(n1095) );
  OR2X2 U927 ( .A(n1144), .B(n1143), .Y(n1096) );
  BUFX2 U928 ( .A(n222), .Y(n1022) );
  AND2X1 U929 ( .A(n1135), .B(n1136), .Y(n221) );
  INVX1 U930 ( .A(n221), .Y(n1023) );
  INVX1 U931 ( .A(n97), .Y(n1024) );
  INVX1 U932 ( .A(n751), .Y(n1025) );
  AND2X1 U933 ( .A(a[3]), .B(n1202), .Y(n1211) );
  INVX1 U934 ( .A(n1211), .Y(n1026) );
  AND2X2 U935 ( .A(a[11]), .B(n1207), .Y(n1215) );
  INVX1 U936 ( .A(n1215), .Y(n1027) );
  AND2X1 U937 ( .A(n1045), .B(n1133), .Y(n111) );
  INVX1 U938 ( .A(n111), .Y(n1028) );
  AND2X1 U939 ( .A(n1093), .B(n1139), .Y(n109) );
  INVX1 U940 ( .A(n109), .Y(n1029) );
  AND2X1 U941 ( .A(n1061), .B(n214), .Y(n105) );
  INVX1 U942 ( .A(n105), .Y(n1030) );
  AND2X1 U943 ( .A(n1047), .B(n181), .Y(n99) );
  INVX1 U944 ( .A(n99), .Y(n1031) );
  BUFX2 U945 ( .A(n183), .Y(n1032) );
  INVX1 U946 ( .A(n98), .Y(n1033) );
  INVX2 U947 ( .A(n177), .Y(n1125) );
  INVX1 U948 ( .A(n289), .Y(n1034) );
  AND2X1 U949 ( .A(a[9]), .B(n1206), .Y(n1214) );
  INVX1 U950 ( .A(n1214), .Y(n1035) );
  INVX1 U951 ( .A(n112), .Y(n1036) );
  AND2X1 U952 ( .A(n1121), .B(n186), .Y(n100) );
  INVX1 U953 ( .A(n100), .Y(n1037) );
  AND2X1 U954 ( .A(n1062), .B(n192), .Y(n101) );
  INVX1 U955 ( .A(n101), .Y(n1038) );
  AND2X1 U956 ( .A(n1078), .B(n162), .Y(n95) );
  INVX1 U957 ( .A(n95), .Y(n1039) );
  AND2X1 U958 ( .A(n1058), .B(n1130), .Y(n91) );
  INVX1 U959 ( .A(n91), .Y(n1040) );
  AND2X1 U960 ( .A(n1057), .B(n1136), .Y(n107) );
  INVX1 U961 ( .A(n107), .Y(n1041) );
  BUFX2 U962 ( .A(n227), .Y(n1042) );
  AND2X1 U963 ( .A(n1079), .B(n143), .Y(n92) );
  INVX1 U964 ( .A(n92), .Y(n1043) );
  AND2X1 U965 ( .A(n381), .B(n368), .Y(n156) );
  INVX1 U966 ( .A(n156), .Y(n1044) );
  AND2X1 U967 ( .A(n550), .B(n549), .Y(n245) );
  INVX1 U968 ( .A(n245), .Y(n1045) );
  AND2X2 U969 ( .A(n426), .B(n412), .Y(n174) );
  INVX1 U970 ( .A(n174), .Y(n1046) );
  AND2X1 U971 ( .A(n454), .B(n441), .Y(n182) );
  INVX1 U972 ( .A(n182), .Y(n1047) );
  BUFX2 U973 ( .A(n211), .Y(n1048) );
  INVX1 U974 ( .A(n212), .Y(n1049) );
  INVX1 U975 ( .A(n179), .Y(n1050) );
  INVX1 U976 ( .A(n299), .Y(n1051) );
  AND2X1 U977 ( .A(b[15]), .B(n1163), .Y(n627) );
  INVX1 U978 ( .A(n627), .Y(n1052) );
  INVX1 U979 ( .A(n94), .Y(n1053) );
  AND2X1 U980 ( .A(n1076), .B(n1131), .Y(n89) );
  INVX1 U981 ( .A(n89), .Y(n1054) );
  AND2X1 U982 ( .A(n1077), .B(n1137), .Y(n103) );
  INVX1 U983 ( .A(n103), .Y(n1055) );
  BUFX2 U984 ( .A(n205), .Y(n1056) );
  AND2X1 U985 ( .A(n534), .B(n529), .Y(n226) );
  INVX1 U986 ( .A(n226), .Y(n1057) );
  AND2X1 U987 ( .A(n334), .B(n343), .Y(n141) );
  INVX1 U988 ( .A(n141), .Y(n1058) );
  AND2X1 U989 ( .A(n548), .B(n545), .Y(n240) );
  INVX1 U990 ( .A(n240), .Y(n1059) );
  AND2X2 U991 ( .A(n878), .B(n551), .Y(n248) );
  INVX1 U992 ( .A(n248), .Y(n1060) );
  AND2X1 U993 ( .A(n520), .B(n513), .Y(n215) );
  INVX1 U994 ( .A(n215), .Y(n1061) );
  AND2X1 U995 ( .A(n480), .B(n469), .Y(n193) );
  INVX1 U996 ( .A(n193), .Y(n1062) );
  AND2X1 U997 ( .A(n367), .B(n356), .Y(n149) );
  INVX1 U998 ( .A(n149), .Y(n1063) );
  BUFX2 U999 ( .A(n178), .Y(n1064) );
  INVX1 U1000 ( .A(n165), .Y(n1065) );
  INVX1 U1001 ( .A(n313), .Y(n1066) );
  AND2X1 U1002 ( .A(n1204), .B(n1203), .Y(n1212) );
  INVX1 U1003 ( .A(n1212), .Y(n1067) );
  AND2X1 U1004 ( .A(b[15]), .B(n1171), .Y(n589) );
  INVX1 U1005 ( .A(n589), .Y(n1068) );
  AND2X1 U1006 ( .A(b[15]), .B(n1167), .Y(n608) );
  INVX1 U1007 ( .A(n608), .Y(n1069) );
  INVX1 U1008 ( .A(n110), .Y(n1070) );
  AND2X1 U1009 ( .A(n1099), .B(n127), .Y(n88) );
  INVX1 U1010 ( .A(n88), .Y(n1071) );
  AND2X1 U1011 ( .A(n1123), .B(n217), .Y(n106) );
  INVX1 U1012 ( .A(n106), .Y(n1072) );
  AND2X1 U1013 ( .A(n1124), .B(n195), .Y(n102) );
  INVX1 U1014 ( .A(n102), .Y(n1073) );
  AND2X1 U1015 ( .A(n1098), .B(n135), .Y(n90) );
  INVX1 U1016 ( .A(n90), .Y(n1074) );
  AND2X1 U1017 ( .A(n302), .B(n307), .Y(n125) );
  INVX1 U1018 ( .A(n125), .Y(n1075) );
  AND2X1 U1019 ( .A(n316), .B(n323), .Y(n133) );
  INVX1 U1020 ( .A(n133), .Y(n1076) );
  AND2X1 U1021 ( .A(n502), .B(n493), .Y(n204) );
  INVX1 U1022 ( .A(n204), .Y(n1077) );
  AND2X1 U1023 ( .A(n395), .B(n382), .Y(n163) );
  INVX1 U1024 ( .A(n163), .Y(n1078) );
  AND2X1 U1025 ( .A(n355), .B(n344), .Y(n144) );
  INVX1 U1026 ( .A(n144), .Y(n1079) );
  BUFX2 U1027 ( .A(n233), .Y(n1080) );
  OR2X1 U1028 ( .A(n551), .B(n878), .Y(n247) );
  INVX1 U1029 ( .A(n247), .Y(n1081) );
  OR2X1 U1030 ( .A(n513), .B(n520), .Y(n214) );
  INVX1 U1031 ( .A(n214), .Y(n1082) );
  OR2X1 U1032 ( .A(n469), .B(n480), .Y(n192) );
  INVX1 U1033 ( .A(n192), .Y(n1083) );
  OR2X1 U1034 ( .A(n441), .B(n454), .Y(n181) );
  INVX1 U1035 ( .A(n181), .Y(n1084) );
  INVX1 U1036 ( .A(n173), .Y(n1085) );
  INVX1 U1037 ( .A(n331), .Y(n1086) );
  AND2X1 U1038 ( .A(b[15]), .B(n1198), .Y(n703) );
  INVX1 U1039 ( .A(n703), .Y(n1087) );
  AND2X1 U1040 ( .A(b[15]), .B(n1155), .Y(n665) );
  INVX1 U1041 ( .A(n665), .Y(n1088) );
  AND2X1 U1042 ( .A(n1113), .B(n1135), .Y(n108) );
  INVX1 U1043 ( .A(n108), .Y(n1089) );
  AND2X1 U1044 ( .A(n1114), .B(n1134), .Y(n104) );
  INVX1 U1045 ( .A(n104), .Y(n1090) );
  AND2X1 U1046 ( .A(n1112), .B(n1138), .Y(n86) );
  INVX1 U1047 ( .A(n86), .Y(n1091) );
  AND2X1 U1048 ( .A(n742), .B(n895), .Y(n254) );
  INVX1 U1049 ( .A(n254), .Y(n1092) );
  AND2X1 U1050 ( .A(n544), .B(n541), .Y(n237) );
  INVX1 U1051 ( .A(n237), .Y(n1093) );
  OR2X1 U1052 ( .A(n455), .B(n468), .Y(n186) );
  INVX1 U1053 ( .A(n186), .Y(n1094) );
  OR2X1 U1054 ( .A(n564), .B(n1210), .Y(n749) );
  INVX1 U1055 ( .A(n749), .Y(n1097) );
  AND2X1 U1056 ( .A(n324), .B(n333), .Y(n136) );
  INVX1 U1057 ( .A(n136), .Y(n1098) );
  AND2X1 U1058 ( .A(n308), .B(n315), .Y(n128) );
  INVX1 U1059 ( .A(n128), .Y(n1099) );
  OR2X1 U1060 ( .A(n344), .B(n355), .Y(n143) );
  INVX1 U1061 ( .A(n143), .Y(n1100) );
  BUFX2 U1062 ( .A(n241), .Y(n1101) );
  OR2X1 U1063 ( .A(n521), .B(n528), .Y(n217) );
  INVX1 U1064 ( .A(n217), .Y(n1102) );
  OR2X1 U1065 ( .A(n481), .B(n492), .Y(n195) );
  INVX1 U1066 ( .A(n195), .Y(n1103) );
  INVX1 U1067 ( .A(n176), .Y(n1104) );
  INVX1 U1068 ( .A(n162), .Y(n1105) );
  INVX1 U1069 ( .A(n353), .Y(n1106) );
  AND2X1 U1070 ( .A(a[13]), .B(n1208), .Y(n1216) );
  INVX1 U1071 ( .A(n1216), .Y(n1107) );
  AND2X1 U1072 ( .A(a[7]), .B(n1205), .Y(n1213) );
  INVX1 U1073 ( .A(n1213), .Y(n1108) );
  AND2X1 U1074 ( .A(b[15]), .B(n1159), .Y(n646) );
  INVX1 U1075 ( .A(n646), .Y(n1109) );
  INVX1 U1076 ( .A(n87), .Y(n1110) );
  INVX1 U1077 ( .A(n2), .Y(n1111) );
  AND2X1 U1078 ( .A(n292), .B(n295), .Y(n119) );
  INVX1 U1079 ( .A(n119), .Y(n1112) );
  AND2X1 U1080 ( .A(n540), .B(n535), .Y(n231) );
  INVX1 U1081 ( .A(n231), .Y(n1113) );
  AND2X1 U1082 ( .A(n512), .B(n503), .Y(n209) );
  INVX1 U1083 ( .A(n209), .Y(n1114) );
  OR2X1 U1084 ( .A(n545), .B(n548), .Y(n239) );
  INVX1 U1085 ( .A(n239), .Y(n1115) );
  OR2X1 U1086 ( .A(n333), .B(n324), .Y(n135) );
  INVX1 U1087 ( .A(n135), .Y(n1116) );
  OR2X1 U1088 ( .A(n315), .B(n308), .Y(n127) );
  INVX1 U1089 ( .A(n127), .Y(n1117) );
  OR2X1 U1090 ( .A(n565), .B(n1210), .Y(n750) );
  INVX1 U1091 ( .A(n750), .Y(n1118) );
  AND2X1 U1092 ( .A(b[15]), .B(n1151), .Y(n684) );
  INVX1 U1093 ( .A(n684), .Y(n1119) );
  AND2X1 U1094 ( .A(n250), .B(n254), .Y(n249) );
  INVX1 U1095 ( .A(n249), .Y(n1120) );
  AND2X1 U1096 ( .A(n468), .B(n455), .Y(n187) );
  INVX1 U1097 ( .A(n187), .Y(n1121) );
  OR2X1 U1098 ( .A(n356), .B(n367), .Y(n148) );
  INVX1 U1099 ( .A(n148), .Y(n1122) );
  AND2X1 U1100 ( .A(n528), .B(n521), .Y(n218) );
  INVX1 U1101 ( .A(n218), .Y(n1123) );
  AND2X1 U1102 ( .A(n492), .B(n481), .Y(n196) );
  INVX1 U1103 ( .A(n196), .Y(n1124) );
  AND2X1 U1104 ( .A(n440), .B(n427), .Y(n177) );
  INVX1 U1105 ( .A(n166), .Y(n1126) );
  INVX1 U1106 ( .A(n379), .Y(n1127) );
  INVX2 U1107 ( .A(n723), .Y(n771) );
  INVX2 U1108 ( .A(n729), .Y(n825) );
  BUFX2 U1109 ( .A(n126), .Y(n1128) );
  INVX1 U1110 ( .A(n993), .Y(n158) );
  INVX1 U1111 ( .A(n161), .Y(n159) );
  INVX1 U1112 ( .A(n1065), .Y(n267) );
  INVX1 U1113 ( .A(n168), .Y(n167) );
  INVX1 U1114 ( .A(n198), .Y(n197) );
  INVX1 U1115 ( .A(n220), .Y(n219) );
  XNOR2X1 U1116 ( .A(n1145), .B(n1071), .Y(product[26]) );
  INVX1 U1117 ( .A(n1080), .Y(n232) );
  INVX1 U1118 ( .A(n1048), .Y(n210) );
  OR2X1 U1119 ( .A(n368), .B(n381), .Y(n1129) );
  INVX1 U1120 ( .A(n121), .Y(n256) );
  OR2X1 U1121 ( .A(n343), .B(n334), .Y(n1130) );
  OR2X1 U1122 ( .A(n323), .B(n316), .Y(n1131) );
  OR2X1 U1123 ( .A(n307), .B(n302), .Y(n1132) );
  OR2X1 U1124 ( .A(n549), .B(n550), .Y(n1133) );
  BUFX2 U1125 ( .A(n36), .Y(n1167) );
  BUFX2 U1126 ( .A(n12), .Y(n1151) );
  BUFX2 U1127 ( .A(n24), .Y(n1158) );
  BUFX2 U1128 ( .A(n36), .Y(n1166) );
  BUFX2 U1129 ( .A(n12), .Y(n1150) );
  BUFX2 U1130 ( .A(n20), .Y(n1160) );
  BUFX2 U1131 ( .A(n8), .Y(n1152) );
  BUFX2 U1132 ( .A(n32), .Y(n1168) );
  BUFX2 U1133 ( .A(n20), .Y(n1161) );
  BUFX2 U1134 ( .A(n8), .Y(n1153) );
  BUFX2 U1135 ( .A(n32), .Y(n1169) );
  INVX1 U1136 ( .A(n115), .Y(n255) );
  OR2X1 U1137 ( .A(n503), .B(n512), .Y(n1134) );
  OR2X1 U1138 ( .A(n535), .B(n540), .Y(n1135) );
  OR2X1 U1139 ( .A(n529), .B(n534), .Y(n1136) );
  OR2X1 U1140 ( .A(n493), .B(n502), .Y(n1137) );
  OR2X1 U1141 ( .A(n295), .B(n292), .Y(n1138) );
  OR2X1 U1142 ( .A(n541), .B(n544), .Y(n1139) );
  XOR2X1 U1143 ( .A(n254), .B(n250), .Y(product[1]) );
  OR2X1 U1144 ( .A(n895), .B(n742), .Y(n1140) );
  BUFX2 U1145 ( .A(n48), .Y(n1175) );
  BUFX2 U1146 ( .A(n18), .Y(n1155) );
  BUFX2 U1147 ( .A(n42), .Y(n1171) );
  BUFX2 U1148 ( .A(n30), .Y(n1163) );
  BUFX2 U1149 ( .A(n18), .Y(n1154) );
  BUFX2 U1150 ( .A(n42), .Y(n1170) );
  BUFX2 U1151 ( .A(n30), .Y(n1162) );
  BUFX2 U1152 ( .A(n44), .Y(n1176) );
  BUFX2 U1153 ( .A(n14), .Y(n1156) );
  BUFX2 U1154 ( .A(n38), .Y(n1172) );
  BUFX2 U1155 ( .A(n26), .Y(n1164) );
  BUFX2 U1156 ( .A(n1111), .Y(n1148) );
  BUFX2 U1157 ( .A(n44), .Y(n1177) );
  BUFX2 U1158 ( .A(n14), .Y(n1157) );
  BUFX2 U1159 ( .A(n38), .Y(n1173) );
  BUFX2 U1160 ( .A(n26), .Y(n1165) );
  BUFX2 U1161 ( .A(n1111), .Y(n1149) );
  INVX1 U1162 ( .A(n1194), .Y(n1193) );
  INVX1 U1163 ( .A(n1187), .Y(n1185) );
  INVX1 U1164 ( .A(n1189), .Y(n1188) );
  INVX1 U1165 ( .A(n1179), .Y(n1178) );
  INVX1 U1166 ( .A(n1201), .Y(n1200) );
  INVX1 U1167 ( .A(n1187), .Y(n1186) );
  INVX1 U1168 ( .A(n1182), .Y(n1181) );
  INVX1 U1169 ( .A(a[13]), .Y(n1209) );
  INVX1 U1170 ( .A(n1197), .Y(n1195) );
  INVX1 U1171 ( .A(a[7]), .Y(n1206) );
  INVX1 U1172 ( .A(b[2]), .Y(n1184) );
  INVX1 U1173 ( .A(b[3]), .Y(n1187) );
  INVX1 U1174 ( .A(b[1]), .Y(n1182) );
  INVX1 U1175 ( .A(b[0]), .Y(n1179) );
  INVX1 U1176 ( .A(b[4]), .Y(n1189) );
  INVX1 U1177 ( .A(n1197), .Y(n1196) );
  INVX1 U1178 ( .A(b[11]), .Y(n1197) );
  INVX1 U1179 ( .A(n1192), .Y(n1190) );
  INVX1 U1180 ( .A(n1192), .Y(n1191) );
  INVX1 U1181 ( .A(b[5]), .Y(n1192) );
  XOR2X1 U1182 ( .A(n462), .B(n449), .Y(n1141) );
  XOR2X1 U1183 ( .A(n1141), .B(n451), .Y(n445) );
  INVX1 U1184 ( .A(n992), .Y(n1145) );
  INVX1 U1185 ( .A(n142), .Y(n1146) );
  INVX1 U1186 ( .A(n1146), .Y(n1147) );
  OAI21X1 U1187 ( .A(a[2]), .B(n1203), .C(n1026), .Y(n733) );
  OAI21X1 U1188 ( .A(a[4]), .B(n1205), .C(n1067), .Y(n731) );
  OAI21X1 U1189 ( .A(a[6]), .B(n1206), .C(n1108), .Y(n729) );
  OAI21X1 U1190 ( .A(a[8]), .B(n1207), .C(n1035), .Y(n727) );
  OAI21X1 U1191 ( .A(a[10]), .B(n1208), .C(n1027), .Y(n725) );
  OAI21X1 U1192 ( .A(a[12]), .B(n1209), .C(n1107), .Y(n723) );
  OAI21X1 U1193 ( .A(a[14]), .B(n1210), .C(n1014), .Y(n721) );
  XOR2X1 U1194 ( .A(n1015), .B(n1034), .Y(n285) );
endmodule


module alu_DW01_sub_17 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n36, n37, n38, n39, n40, n44, n45, n46, n47, n48, n52, n53,
         n54, n55, n56, n60, n61, n62, n63, n64, n68, n69, n70, n71, n72, n76,
         n77, n78, n79, n80, n84, n85, n86, n87, n88, n92, n93, n94, n95, n96,
         n100, n101, n102, n103, n104, n108, n110, n111, n112, n116, n117,
         n118, n119, n123, n124, n125, n126, n127, n128, n129, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n172, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461;

  XOR2X1 U1 ( .A(n29), .B(n1), .Y(DIFF[31]) );
  FAX1 U3 ( .A(n461), .B(A[30]), .C(n30), .YC(n29), .YS(DIFF[30]) );
  FAX1 U4 ( .A(n460), .B(A[29]), .C(n31), .YC(n30), .YS(DIFF[29]) );
  FAX1 U5 ( .A(n459), .B(A[28]), .C(n148), .YC(n31), .YS(DIFF[28]) );
  XNOR2X1 U7 ( .A(n409), .B(n392), .Y(DIFF[27]) );
  AOI21X1 U8 ( .A(n37), .B(n422), .C(n36), .Y(n32) );
  OAI21X1 U16 ( .A(n401), .B(n323), .C(n352), .Y(n37) );
  XNOR2X1 U21 ( .A(n45), .B(n334), .Y(DIFF[25]) );
  AOI21X1 U22 ( .A(n45), .B(n424), .C(n44), .Y(n40) );
  OAI21X1 U30 ( .A(n319), .B(n322), .C(n359), .Y(n45) );
  XNOR2X1 U35 ( .A(n408), .B(n391), .Y(DIFF[23]) );
  AOI21X1 U36 ( .A(n310), .B(n423), .C(n52), .Y(n48) );
  OAI21X1 U44 ( .A(n360), .B(n321), .C(n358), .Y(n53) );
  XNOR2X1 U49 ( .A(n430), .B(n331), .Y(DIFF[21]) );
  AOI21X1 U50 ( .A(n61), .B(n415), .C(n60), .Y(n56) );
  XOR2X1 U57 ( .A(n372), .B(n340), .Y(DIFF[20]) );
  OAI21X1 U58 ( .A(n318), .B(n372), .C(n357), .Y(n61) );
  XNOR2X1 U63 ( .A(n69), .B(n330), .Y(DIFF[19]) );
  AOI21X1 U64 ( .A(n69), .B(n416), .C(n68), .Y(n64) );
  XOR2X1 U71 ( .A(n369), .B(n339), .Y(DIFF[18]) );
  OAI21X1 U72 ( .A(n317), .B(n370), .C(n356), .Y(n69) );
  XNOR2X1 U77 ( .A(n311), .B(n329), .Y(DIFF[17]) );
  AOI21X1 U78 ( .A(n77), .B(n417), .C(n76), .Y(n72) );
  XOR2X1 U85 ( .A(n367), .B(n338), .Y(DIFF[16]) );
  OAI21X1 U86 ( .A(n316), .B(n320), .C(n355), .Y(n77) );
  XNOR2X1 U91 ( .A(n85), .B(n328), .Y(DIFF[15]) );
  AOI21X1 U92 ( .A(n85), .B(n418), .C(n84), .Y(n80) );
  XOR2X1 U99 ( .A(n365), .B(n337), .Y(DIFF[14]) );
  OAI21X1 U100 ( .A(n315), .B(n366), .C(n354), .Y(n85) );
  XNOR2X1 U105 ( .A(n93), .B(n327), .Y(DIFF[13]) );
  AOI21X1 U106 ( .A(n93), .B(n421), .C(n92), .Y(n88) );
  XOR2X1 U113 ( .A(n362), .B(n336), .Y(DIFF[12]) );
  OAI21X1 U114 ( .A(n314), .B(n363), .C(n353), .Y(n93) );
  XNOR2X1 U119 ( .A(n407), .B(n390), .Y(DIFF[11]) );
  AOI21X1 U120 ( .A(n101), .B(n420), .C(n100), .Y(n96) );
  OAI21X1 U128 ( .A(n402), .B(n388), .C(n394), .Y(n101) );
  XNOR2X1 U133 ( .A(n428), .B(n379), .Y(DIFF[9]) );
  AOI21X1 U134 ( .A(n428), .B(n414), .C(n108), .Y(n104) );
  XOR2X1 U141 ( .A(n410), .B(n380), .Y(DIFF[8]) );
  XNOR2X1 U147 ( .A(n406), .B(n389), .Y(DIFF[7]) );
  AOI21X1 U148 ( .A(n117), .B(n419), .C(n116), .Y(n112) );
  XOR2X1 U155 ( .A(n326), .B(n335), .Y(DIFF[6]) );
  OAI21X1 U156 ( .A(n313), .B(n381), .C(n325), .Y(n117) );
  AOI21X1 U158 ( .A(n126), .B(n413), .C(n123), .Y(n119) );
  XOR2X1 U165 ( .A(n377), .B(n376), .Y(DIFF[5]) );
  AOI21X1 U166 ( .A(n134), .B(n312), .C(n126), .Y(n124) );
  OAI21X1 U168 ( .A(n397), .B(n403), .C(n386), .Y(n126) );
  XNOR2X1 U173 ( .A(n134), .B(n374), .Y(DIFF[4]) );
  AOI21X1 U174 ( .A(n134), .B(n172), .C(n133), .Y(n129) );
  XNOR2X1 U181 ( .A(n140), .B(n375), .Y(DIFF[3]) );
  AOI21X1 U183 ( .A(n144), .B(n382), .C(n137), .Y(n135) );
  OAI21X1 U185 ( .A(n404), .B(n398), .C(n385), .Y(n137) );
  XOR2X1 U190 ( .A(n143), .B(n383), .Y(DIFF[2]) );
  OAI21X1 U191 ( .A(n141), .B(n143), .C(n404), .Y(n140) );
  XOR2X1 U196 ( .A(n378), .B(n396), .Y(DIFF[1]) );
  OAI21X1 U198 ( .A(n396), .B(n387), .C(n373), .Y(n144) );
  XNOR2X1 U203 ( .A(n431), .B(A[0]), .Y(DIFF[0]) );
  OR2X1 U240 ( .A(A[6]), .B(n437), .Y(n413) );
  OR2X1 U241 ( .A(A[5]), .B(n436), .Y(n127) );
  AND2X1 U242 ( .A(A[5]), .B(n436), .Y(n128) );
  OR2X1 U243 ( .A(n434), .B(A[3]), .Y(n138) );
  AND2X1 U244 ( .A(A[3]), .B(n434), .Y(n139) );
  OR2X1 U245 ( .A(n433), .B(A[2]), .Y(n411) );
  AND2X1 U246 ( .A(A[2]), .B(n433), .Y(n142) );
  AND2X1 U247 ( .A(n344), .B(n422), .Y(n2) );
  AND2X1 U248 ( .A(n352), .B(n38), .Y(n3) );
  INVX1 U249 ( .A(n371), .Y(n372) );
  AND2X1 U250 ( .A(n343), .B(n420), .Y(n18) );
  AND2X1 U251 ( .A(n394), .B(n102), .Y(n19) );
  AND2X1 U252 ( .A(n342), .B(n414), .Y(n20) );
  AND2X1 U253 ( .A(n341), .B(n419), .Y(n22) );
  OR2X1 U254 ( .A(n431), .B(A[0]), .Y(n147) );
  AND2X1 U255 ( .A(n373), .B(n145), .Y(n28) );
  INVX1 U256 ( .A(B[0]), .Y(n431) );
  OAI21X1 U257 ( .A(n360), .B(n321), .C(n358), .Y(n310) );
  BUFX2 U258 ( .A(n77), .Y(n311) );
  OR2X2 U259 ( .A(n432), .B(A[1]), .Y(n145) );
  AND2X1 U260 ( .A(n437), .B(A[6]), .Y(n123) );
  OR2X1 U261 ( .A(A[12]), .B(n443), .Y(n94) );
  OR2X1 U262 ( .A(n384), .B(n403), .Y(n125) );
  INVX1 U263 ( .A(n127), .Y(n403) );
  OR2X1 U264 ( .A(A[10]), .B(n441), .Y(n102) );
  OR2X1 U265 ( .A(n435), .B(A[4]), .Y(n132) );
  AND2X1 U266 ( .A(A[4]), .B(n435), .Y(n133) );
  AND2X2 U267 ( .A(A[1]), .B(n432), .Y(n146) );
  INVX1 U268 ( .A(n125), .Y(n312) );
  AND2X2 U269 ( .A(n441), .B(A[10]), .Y(n103) );
  AND2X2 U270 ( .A(n413), .B(n312), .Y(n118) );
  INVX1 U271 ( .A(n118), .Y(n313) );
  INVX1 U272 ( .A(n94), .Y(n314) );
  OR2X1 U273 ( .A(A[14]), .B(n445), .Y(n86) );
  INVX1 U274 ( .A(n86), .Y(n315) );
  OR2X1 U275 ( .A(A[16]), .B(n447), .Y(n78) );
  INVX1 U276 ( .A(n78), .Y(n316) );
  OR2X1 U277 ( .A(n449), .B(A[18]), .Y(n70) );
  INVX1 U278 ( .A(n70), .Y(n317) );
  OR2X1 U279 ( .A(A[20]), .B(n451), .Y(n62) );
  INVX1 U280 ( .A(n62), .Y(n318) );
  OR2X1 U281 ( .A(A[24]), .B(n455), .Y(n46) );
  INVX1 U282 ( .A(n46), .Y(n319) );
  BUFX2 U283 ( .A(n80), .Y(n320) );
  BUFX2 U284 ( .A(n56), .Y(n321) );
  BUFX2 U285 ( .A(n48), .Y(n322) );
  BUFX2 U286 ( .A(n40), .Y(n323) );
  INVX1 U287 ( .A(n119), .Y(n324) );
  INVX1 U288 ( .A(n324), .Y(n325) );
  BUFX2 U289 ( .A(n124), .Y(n326) );
  AND2X1 U290 ( .A(n346), .B(n421), .Y(n16) );
  INVX1 U291 ( .A(n16), .Y(n327) );
  AND2X1 U292 ( .A(n347), .B(n418), .Y(n14) );
  INVX1 U293 ( .A(n14), .Y(n328) );
  AND2X1 U294 ( .A(n348), .B(n417), .Y(n12) );
  INVX1 U295 ( .A(n12), .Y(n329) );
  AND2X1 U296 ( .A(n349), .B(n416), .Y(n10) );
  INVX1 U297 ( .A(n10), .Y(n330) );
  AND2X1 U298 ( .A(n350), .B(n415), .Y(n8) );
  INVX1 U299 ( .A(n8), .Y(n331) );
  AND2X1 U300 ( .A(n358), .B(n54), .Y(n7) );
  INVX1 U301 ( .A(n7), .Y(n332) );
  AND2X1 U302 ( .A(n359), .B(n46), .Y(n5) );
  INVX1 U303 ( .A(n5), .Y(n333) );
  AND2X1 U304 ( .A(n351), .B(n424), .Y(n4) );
  INVX1 U305 ( .A(n4), .Y(n334) );
  AND2X1 U306 ( .A(n345), .B(n413), .Y(n23) );
  INVX1 U307 ( .A(n23), .Y(n335) );
  AND2X1 U308 ( .A(n353), .B(n94), .Y(n17) );
  INVX1 U309 ( .A(n17), .Y(n336) );
  AND2X1 U310 ( .A(n354), .B(n86), .Y(n15) );
  INVX1 U311 ( .A(n15), .Y(n337) );
  AND2X1 U312 ( .A(n355), .B(n78), .Y(n13) );
  INVX1 U313 ( .A(n13), .Y(n338) );
  AND2X1 U314 ( .A(n356), .B(n70), .Y(n11) );
  INVX1 U315 ( .A(n11), .Y(n339) );
  AND2X1 U316 ( .A(n357), .B(n62), .Y(n9) );
  INVX1 U317 ( .A(n9), .Y(n340) );
  AND2X1 U318 ( .A(n438), .B(A[7]), .Y(n116) );
  INVX1 U319 ( .A(n116), .Y(n341) );
  AND2X1 U320 ( .A(n440), .B(A[9]), .Y(n108) );
  INVX1 U321 ( .A(n108), .Y(n342) );
  AND2X1 U322 ( .A(n442), .B(A[11]), .Y(n100) );
  INVX1 U323 ( .A(n100), .Y(n343) );
  AND2X1 U324 ( .A(n458), .B(A[27]), .Y(n36) );
  INVX1 U325 ( .A(n36), .Y(n344) );
  INVX1 U326 ( .A(n123), .Y(n345) );
  AND2X1 U327 ( .A(n444), .B(A[13]), .Y(n92) );
  INVX1 U328 ( .A(n92), .Y(n346) );
  AND2X1 U329 ( .A(n446), .B(A[15]), .Y(n84) );
  INVX1 U330 ( .A(n84), .Y(n347) );
  AND2X1 U331 ( .A(n448), .B(A[17]), .Y(n76) );
  INVX1 U332 ( .A(n76), .Y(n348) );
  AND2X1 U333 ( .A(n450), .B(A[19]), .Y(n68) );
  INVX1 U334 ( .A(n68), .Y(n349) );
  AND2X1 U335 ( .A(n452), .B(A[21]), .Y(n60) );
  INVX1 U336 ( .A(n60), .Y(n350) );
  AND2X1 U337 ( .A(n456), .B(A[25]), .Y(n44) );
  INVX1 U338 ( .A(n44), .Y(n351) );
  AND2X1 U339 ( .A(n457), .B(A[26]), .Y(n39) );
  INVX1 U340 ( .A(n39), .Y(n352) );
  AND2X1 U341 ( .A(n443), .B(A[12]), .Y(n95) );
  INVX1 U342 ( .A(n95), .Y(n353) );
  AND2X1 U343 ( .A(n445), .B(A[14]), .Y(n87) );
  INVX1 U344 ( .A(n87), .Y(n354) );
  AND2X1 U345 ( .A(n447), .B(A[16]), .Y(n79) );
  INVX1 U346 ( .A(n79), .Y(n355) );
  AND2X1 U347 ( .A(A[18]), .B(n449), .Y(n71) );
  INVX1 U348 ( .A(n71), .Y(n356) );
  AND2X1 U349 ( .A(n451), .B(A[20]), .Y(n63) );
  INVX1 U350 ( .A(n63), .Y(n357) );
  AND2X1 U351 ( .A(n453), .B(A[22]), .Y(n55) );
  INVX1 U352 ( .A(n55), .Y(n358) );
  AND2X1 U353 ( .A(n455), .B(A[24]), .Y(n47) );
  INVX1 U354 ( .A(n47), .Y(n359) );
  OR2X1 U355 ( .A(A[22]), .B(n453), .Y(n54) );
  INVX1 U356 ( .A(n54), .Y(n360) );
  INVX1 U357 ( .A(n96), .Y(n361) );
  INVX1 U358 ( .A(n361), .Y(n362) );
  INVX1 U359 ( .A(n361), .Y(n363) );
  INVX1 U360 ( .A(n88), .Y(n364) );
  INVX1 U361 ( .A(n364), .Y(n365) );
  INVX1 U362 ( .A(n364), .Y(n366) );
  BUFX2 U363 ( .A(n320), .Y(n367) );
  INVX1 U364 ( .A(n72), .Y(n368) );
  INVX1 U365 ( .A(n368), .Y(n369) );
  INVX1 U366 ( .A(n368), .Y(n370) );
  INVX1 U367 ( .A(n64), .Y(n371) );
  INVX1 U368 ( .A(n146), .Y(n373) );
  AND2X1 U369 ( .A(n397), .B(n172), .Y(n25) );
  INVX1 U370 ( .A(n25), .Y(n374) );
  AND2X1 U371 ( .A(n385), .B(n138), .Y(n26) );
  INVX1 U372 ( .A(n26), .Y(n375) );
  AND2X1 U373 ( .A(n386), .B(n127), .Y(n24) );
  INVX1 U374 ( .A(n24), .Y(n376) );
  BUFX2 U375 ( .A(n129), .Y(n377) );
  INVX1 U376 ( .A(n28), .Y(n378) );
  INVX1 U377 ( .A(n20), .Y(n379) );
  AND2X1 U378 ( .A(n395), .B(n110), .Y(n21) );
  INVX1 U379 ( .A(n21), .Y(n380) );
  BUFX2 U380 ( .A(n135), .Y(n381) );
  OR2X1 U381 ( .A(n398), .B(n141), .Y(n136) );
  INVX1 U382 ( .A(n136), .Y(n382) );
  AND2X1 U383 ( .A(n404), .B(n411), .Y(n27) );
  INVX1 U384 ( .A(n27), .Y(n383) );
  INVX1 U385 ( .A(n132), .Y(n384) );
  INVX1 U386 ( .A(n139), .Y(n385) );
  INVX1 U387 ( .A(n128), .Y(n386) );
  INVX1 U388 ( .A(n145), .Y(n387) );
  BUFX2 U389 ( .A(n104), .Y(n388) );
  INVX1 U390 ( .A(n22), .Y(n389) );
  INVX1 U391 ( .A(n18), .Y(n390) );
  AND2X1 U392 ( .A(n400), .B(n423), .Y(n6) );
  INVX1 U393 ( .A(n6), .Y(n391) );
  INVX1 U394 ( .A(n2), .Y(n392) );
  INVX1 U395 ( .A(n3), .Y(n393) );
  INVX1 U396 ( .A(n103), .Y(n394) );
  AND2X1 U397 ( .A(n439), .B(A[8]), .Y(n111) );
  INVX1 U398 ( .A(n111), .Y(n395) );
  INVX1 U399 ( .A(n147), .Y(n396) );
  INVX1 U400 ( .A(n133), .Y(n397) );
  INVX1 U401 ( .A(n138), .Y(n398) );
  INVX1 U402 ( .A(n19), .Y(n399) );
  AND2X1 U403 ( .A(n454), .B(A[23]), .Y(n52) );
  INVX1 U404 ( .A(n52), .Y(n400) );
  OR2X1 U405 ( .A(A[26]), .B(n457), .Y(n38) );
  INVX1 U406 ( .A(n38), .Y(n401) );
  INVX1 U407 ( .A(n102), .Y(n402) );
  INVX1 U408 ( .A(n142), .Y(n404) );
  OR2X1 U409 ( .A(A[8]), .B(n439), .Y(n110) );
  INVX1 U410 ( .A(n110), .Y(n405) );
  BUFX2 U411 ( .A(n117), .Y(n406) );
  BUFX2 U412 ( .A(n101), .Y(n407) );
  BUFX2 U413 ( .A(n53), .Y(n408) );
  INVX1 U414 ( .A(n411), .Y(n141) );
  BUFX2 U415 ( .A(n37), .Y(n409) );
  BUFX2 U416 ( .A(n112), .Y(n410) );
  XNOR2X1 U417 ( .A(n412), .B(n399), .Y(DIFF[10]) );
  INVX1 U418 ( .A(n388), .Y(n412) );
  INVX1 U419 ( .A(n144), .Y(n143) );
  INVX1 U420 ( .A(n381), .Y(n134) );
  XNOR2X1 U421 ( .A(n426), .B(n393), .Y(DIFF[26]) );
  XNOR2X1 U422 ( .A(n425), .B(n333), .Y(DIFF[24]) );
  XNOR2X1 U423 ( .A(n427), .B(n332), .Y(DIFF[22]) );
  OR2X1 U424 ( .A(A[9]), .B(n440), .Y(n414) );
  INVX1 U425 ( .A(n384), .Y(n172) );
  INVX1 U426 ( .A(B[18]), .Y(n449) );
  OR2X1 U427 ( .A(A[21]), .B(n452), .Y(n415) );
  INVX1 U428 ( .A(B[19]), .Y(n450) );
  OR2X1 U429 ( .A(A[19]), .B(n450), .Y(n416) );
  INVX1 U430 ( .A(B[16]), .Y(n447) );
  INVX1 U431 ( .A(B[9]), .Y(n440) );
  INVX1 U432 ( .A(B[6]), .Y(n437) );
  INVX1 U433 ( .A(B[2]), .Y(n433) );
  OR2X1 U434 ( .A(A[17]), .B(n448), .Y(n417) );
  OR2X1 U435 ( .A(A[15]), .B(n446), .Y(n418) );
  OR2X1 U436 ( .A(A[7]), .B(n438), .Y(n419) );
  OR2X1 U437 ( .A(A[11]), .B(n442), .Y(n420) );
  OR2X1 U438 ( .A(A[13]), .B(n444), .Y(n421) );
  INVX1 U439 ( .A(B[3]), .Y(n434) );
  INVX1 U440 ( .A(B[1]), .Y(n432) );
  INVX1 U441 ( .A(B[4]), .Y(n435) );
  OR2X1 U442 ( .A(A[27]), .B(n458), .Y(n422) );
  INVX1 U443 ( .A(B[26]), .Y(n457) );
  INVX1 U444 ( .A(B[24]), .Y(n455) );
  INVX1 U445 ( .A(B[25]), .Y(n456) );
  OR2X1 U446 ( .A(A[23]), .B(n454), .Y(n423) );
  OR2X1 U447 ( .A(A[25]), .B(n456), .Y(n424) );
  INVX1 U448 ( .A(B[29]), .Y(n460) );
  INVX1 U449 ( .A(B[28]), .Y(n459) );
  XNOR2X1 U450 ( .A(A[31]), .B(B[31]), .Y(n1) );
  INVX1 U451 ( .A(B[30]), .Y(n461) );
  INVX1 U452 ( .A(B[12]), .Y(n443) );
  INVX1 U453 ( .A(B[13]), .Y(n444) );
  INVX1 U454 ( .A(B[11]), .Y(n442) );
  INVX1 U455 ( .A(B[14]), .Y(n445) );
  INVX1 U456 ( .A(B[7]), .Y(n438) );
  INVX1 U457 ( .A(B[22]), .Y(n453) );
  INVX1 U458 ( .A(B[21]), .Y(n452) );
  INVX1 U459 ( .A(B[15]), .Y(n446) );
  INVX1 U460 ( .A(B[27]), .Y(n458) );
  INVX1 U461 ( .A(B[23]), .Y(n454) );
  INVX1 U462 ( .A(B[5]), .Y(n436) );
  INVX1 U463 ( .A(B[10]), .Y(n441) );
  INVX1 U464 ( .A(B[17]), .Y(n448) );
  INVX1 U465 ( .A(B[20]), .Y(n451) );
  INVX1 U466 ( .A(B[8]), .Y(n439) );
  INVX1 U467 ( .A(n322), .Y(n425) );
  INVX1 U468 ( .A(n323), .Y(n426) );
  INVX1 U469 ( .A(n321), .Y(n427) );
  OAI21X1 U470 ( .A(n405), .B(n410), .C(n395), .Y(n428) );
  INVX1 U471 ( .A(n61), .Y(n429) );
  INVX1 U472 ( .A(n429), .Y(n430) );
  INVX1 U473 ( .A(n32), .Y(n148) );
endmodule


module alu_DW01_add_16 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n29, n30, n31,
         n32, n33, n34, n35, n36, n40, n41, n42, n43, n44, n48, n49, n50, n51,
         n52, n56, n57, n58, n59, n60, n64, n66, n67, n68, n72, n73, n74, n75,
         n76, n80, n81, n82, n83, n84, n88, n89, n90, n91, n92, n96, n97, n98,
         n99, n100, n104, n105, n106, n107, n108, n112, n114, n115, n119, n120,
         n121, n122, n123, n124, n125, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n144, n167,
         n170, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398;

  FAX1 U3 ( .A(B[30]), .B(A[30]), .C(n30), .YC(n29), .YS(SUM[30]) );
  FAX1 U4 ( .A(B[29]), .B(A[29]), .C(n31), .YC(n30), .YS(SUM[29]) );
  FAX1 U5 ( .A(B[28]), .B(A[28]), .C(n32), .YC(n31), .YS(SUM[28]) );
  FAX1 U6 ( .A(B[27]), .B(A[27]), .C(n33), .YC(n32), .YS(SUM[27]) );
  XOR2X1 U7 ( .A(n350), .B(n322), .Y(SUM[26]) );
  OAI21X1 U8 ( .A(n301), .B(n303), .C(n337), .Y(n33) );
  XNOR2X1 U13 ( .A(n277), .B(n361), .Y(SUM[25]) );
  AOI21X1 U14 ( .A(n41), .B(n384), .C(n40), .Y(n36) );
  XOR2X1 U21 ( .A(n293), .B(n321), .Y(SUM[24]) );
  OAI21X1 U22 ( .A(n300), .B(n306), .C(n336), .Y(n41) );
  XNOR2X1 U27 ( .A(n285), .B(n360), .Y(SUM[23]) );
  AOI21X1 U28 ( .A(n49), .B(n388), .C(n48), .Y(n44) );
  XOR2X1 U35 ( .A(n292), .B(n320), .Y(SUM[22]) );
  OAI21X1 U36 ( .A(n343), .B(n305), .C(n335), .Y(n49) );
  XNOR2X1 U41 ( .A(n288), .B(n378), .Y(SUM[21]) );
  AOI21X1 U42 ( .A(n57), .B(n387), .C(n56), .Y(n52) );
  XOR2X1 U49 ( .A(n283), .B(n319), .Y(SUM[20]) );
  OAI21X1 U50 ( .A(n342), .B(n304), .C(n334), .Y(n57) );
  XNOR2X1 U55 ( .A(n276), .B(n377), .Y(SUM[19]) );
  AOI21X1 U56 ( .A(n398), .B(n385), .C(n64), .Y(n60) );
  XOR2X1 U63 ( .A(n291), .B(n362), .Y(SUM[18]) );
  XNOR2X1 U69 ( .A(n274), .B(n376), .Y(SUM[17]) );
  AOI21X1 U70 ( .A(n73), .B(n392), .C(n72), .Y(n68) );
  XOR2X1 U77 ( .A(n294), .B(n318), .Y(SUM[16]) );
  OAI21X1 U78 ( .A(n341), .B(n349), .C(n333), .Y(n73) );
  XNOR2X1 U83 ( .A(n278), .B(n375), .Y(SUM[15]) );
  AOI21X1 U84 ( .A(n81), .B(n386), .C(n80), .Y(n76) );
  XOR2X1 U91 ( .A(n286), .B(n317), .Y(SUM[14]) );
  OAI21X1 U92 ( .A(n299), .B(n347), .C(n332), .Y(n81) );
  XNOR2X1 U97 ( .A(n289), .B(n374), .Y(SUM[13]) );
  AOI21X1 U98 ( .A(n89), .B(n391), .C(n88), .Y(n84) );
  XOR2X1 U105 ( .A(n287), .B(n316), .Y(SUM[12]) );
  OAI21X1 U106 ( .A(n340), .B(n302), .C(n331), .Y(n89) );
  XNOR2X1 U111 ( .A(n290), .B(n373), .Y(SUM[11]) );
  AOI21X1 U112 ( .A(n97), .B(n390), .C(n96), .Y(n92) );
  XOR2X1 U119 ( .A(n284), .B(n315), .Y(SUM[10]) );
  OAI21X1 U120 ( .A(n339), .B(n359), .C(n330), .Y(n97) );
  XNOR2X1 U125 ( .A(n275), .B(n372), .Y(SUM[9]) );
  AOI21X1 U126 ( .A(n105), .B(n383), .C(n104), .Y(n100) );
  XOR2X1 U133 ( .A(n295), .B(n314), .Y(SUM[8]) );
  OAI21X1 U134 ( .A(n338), .B(n370), .C(n329), .Y(n105) );
  XNOR2X1 U139 ( .A(n279), .B(n356), .Y(SUM[7]) );
  AOI21X1 U140 ( .A(n395), .B(n389), .C(n112), .Y(n108) );
  XOR2X1 U147 ( .A(n308), .B(n313), .Y(SUM[6]) );
  AOI21X1 U150 ( .A(n122), .B(n282), .C(n119), .Y(n115) );
  XOR2X1 U157 ( .A(n307), .B(n312), .Y(SUM[5]) );
  AOI21X1 U158 ( .A(n130), .B(n345), .C(n122), .Y(n120) );
  OAI21X1 U160 ( .A(n352), .B(n351), .C(n328), .Y(n122) );
  XNOR2X1 U165 ( .A(n130), .B(n310), .Y(SUM[4]) );
  AOI21X1 U166 ( .A(n130), .B(n167), .C(n129), .Y(n125) );
  XNOR2X1 U173 ( .A(n136), .B(n355), .Y(SUM[3]) );
  AOI21X1 U175 ( .A(n140), .B(n381), .C(n133), .Y(n131) );
  OAI21X1 U177 ( .A(n354), .B(n371), .C(n353), .Y(n133) );
  XOR2X1 U182 ( .A(n139), .B(n311), .Y(SUM[2]) );
  OAI21X1 U183 ( .A(n280), .B(n139), .C(n394), .Y(n136) );
  XOR2X1 U188 ( .A(n309), .B(n281), .Y(SUM[1]) );
  OAI21X1 U190 ( .A(n281), .B(n344), .C(n327), .Y(n140) );
  AND2X2 U203 ( .A(B[25]), .B(A[25]), .Y(n40) );
  OR2X2 U204 ( .A(A[10]), .B(B[10]), .Y(n98) );
  AND2X2 U205 ( .A(B[10]), .B(A[10]), .Y(n99) );
  OR2X1 U206 ( .A(A[23]), .B(B[23]), .Y(n388) );
  OR2X1 U207 ( .A(A[21]), .B(B[21]), .Y(n387) );
  OR2X1 U208 ( .A(A[19]), .B(B[19]), .Y(n385) );
  OR2X1 U209 ( .A(A[13]), .B(B[13]), .Y(n391) );
  OR2X1 U210 ( .A(n280), .B(n371), .Y(n132) );
  AND2X1 U211 ( .A(A[2]), .B(B[2]), .Y(n138) );
  AND2X1 U212 ( .A(B[26]), .B(A[26]), .Y(n35) );
  AND2X1 U213 ( .A(B[24]), .B(A[24]), .Y(n43) );
  AND2X1 U214 ( .A(B[22]), .B(A[22]), .Y(n51) );
  AND2X1 U215 ( .A(B[18]), .B(A[18]), .Y(n67) );
  AND2X1 U216 ( .A(B[16]), .B(A[16]), .Y(n75) );
  AND2X1 U217 ( .A(B[12]), .B(A[12]), .Y(n91) );
  AND2X1 U218 ( .A(B[8]), .B(A[8]), .Y(n107) );
  AND2X1 U219 ( .A(n345), .B(n382), .Y(n114) );
  OR2X1 U220 ( .A(B[6]), .B(A[6]), .Y(n382) );
  AND2X1 U221 ( .A(A[3]), .B(B[3]), .Y(n135) );
  OR2X1 U222 ( .A(A[1]), .B(B[1]), .Y(n141) );
  AND2X1 U223 ( .A(n357), .B(n384), .Y(n3) );
  AND2X1 U224 ( .A(n324), .B(n388), .Y(n5) );
  AND2X1 U225 ( .A(n367), .B(n387), .Y(n7) );
  AND2X1 U226 ( .A(n369), .B(n385), .Y(n9) );
  AND2X1 U227 ( .A(n358), .B(n66), .Y(n10) );
  AND2X1 U228 ( .A(n368), .B(n392), .Y(n11) );
  AND2X1 U229 ( .A(n365), .B(n386), .Y(n13) );
  AND2X1 U230 ( .A(n366), .B(n391), .Y(n15) );
  AND2X1 U231 ( .A(n364), .B(n390), .Y(n17) );
  AND2X1 U232 ( .A(n363), .B(n383), .Y(n19) );
  AND2X1 U233 ( .A(n323), .B(n389), .Y(n21) );
  AND2X1 U234 ( .A(n325), .B(n282), .Y(n22) );
  AND2X1 U235 ( .A(n351), .B(n167), .Y(n24) );
  AND2X1 U236 ( .A(n353), .B(n134), .Y(n25) );
  INVX1 U237 ( .A(n141), .Y(n344) );
  AND2X2 U238 ( .A(A[4]), .B(B[4]), .Y(n129) );
  OR2X1 U239 ( .A(B[4]), .B(A[4]), .Y(n128) );
  AND2X2 U240 ( .A(B[9]), .B(A[9]), .Y(n104) );
  AND2X2 U241 ( .A(B[11]), .B(A[11]), .Y(n96) );
  AND2X1 U242 ( .A(B[7]), .B(A[7]), .Y(n112) );
  AND2X1 U243 ( .A(B[23]), .B(A[23]), .Y(n48) );
  OR2X1 U244 ( .A(A[16]), .B(B[16]), .Y(n74) );
  AND2X1 U245 ( .A(B[15]), .B(A[15]), .Y(n80) );
  OR2X1 U246 ( .A(A[26]), .B(B[26]), .Y(n34) );
  OR2X1 U247 ( .A(A[12]), .B(B[12]), .Y(n90) );
  OR2X1 U248 ( .A(A[24]), .B(B[24]), .Y(n42) );
  AND2X1 U249 ( .A(B[13]), .B(A[13]), .Y(n88) );
  AND2X1 U250 ( .A(B[17]), .B(A[17]), .Y(n72) );
  AND2X1 U251 ( .A(B[19]), .B(A[19]), .Y(n64) );
  AND2X1 U252 ( .A(B[21]), .B(A[21]), .Y(n56) );
  OR2X1 U253 ( .A(A[14]), .B(B[14]), .Y(n82) );
  OR2X1 U254 ( .A(n326), .B(n352), .Y(n121) );
  AND2X1 U255 ( .A(A[0]), .B(B[0]), .Y(n144) );
  OR2X1 U256 ( .A(B[2]), .B(A[2]), .Y(n137) );
  OR2X1 U257 ( .A(A[8]), .B(B[8]), .Y(n106) );
  OR2X1 U258 ( .A(A[22]), .B(B[22]), .Y(n50) );
  OR2X1 U259 ( .A(B[3]), .B(A[3]), .Y(n134) );
  AND2X1 U260 ( .A(n281), .B(n393), .Y(SUM[0]) );
  OR2X2 U261 ( .A(A[11]), .B(B[11]), .Y(n390) );
  OR2X1 U262 ( .A(A[5]), .B(B[5]), .Y(n123) );
  AND2X1 U263 ( .A(B[5]), .B(A[5]), .Y(n124) );
  BUFX2 U264 ( .A(n73), .Y(n274) );
  OAI21X1 U265 ( .A(n338), .B(n370), .C(n329), .Y(n275) );
  BUFX2 U266 ( .A(n398), .Y(n276) );
  OAI21X1 U267 ( .A(n300), .B(n306), .C(n336), .Y(n277) );
  BUFX2 U268 ( .A(n81), .Y(n278) );
  OAI21X1 U269 ( .A(n380), .B(n298), .C(n297), .Y(n279) );
  INVX1 U270 ( .A(n137), .Y(n280) );
  INVX1 U271 ( .A(n144), .Y(n281) );
  OR2X2 U272 ( .A(B[6]), .B(A[6]), .Y(n282) );
  BUFX2 U273 ( .A(n304), .Y(n283) );
  BUFX2 U274 ( .A(n359), .Y(n284) );
  OAI21X1 U275 ( .A(n343), .B(n292), .C(n335), .Y(n285) );
  BUFX2 U276 ( .A(n347), .Y(n286) );
  BUFX2 U277 ( .A(n302), .Y(n287) );
  AND2X1 U278 ( .A(A[1]), .B(B[1]), .Y(n142) );
  OAI21X1 U279 ( .A(n342), .B(n283), .C(n334), .Y(n288) );
  OAI21X1 U280 ( .A(n340), .B(n287), .C(n331), .Y(n289) );
  OAI21X1 U281 ( .A(n339), .B(n284), .C(n330), .Y(n290) );
  AND2X2 U282 ( .A(B[6]), .B(A[6]), .Y(n119) );
  BUFX2 U283 ( .A(n397), .Y(n291) );
  INVX1 U284 ( .A(n396), .Y(n397) );
  BUFX2 U285 ( .A(n305), .Y(n292) );
  BUFX2 U286 ( .A(n306), .Y(n293) );
  BUFX2 U287 ( .A(n349), .Y(n294) );
  BUFX2 U288 ( .A(n370), .Y(n295) );
  XNOR2X1 U289 ( .A(n29), .B(n296), .Y(SUM[31]) );
  XNOR2X1 U290 ( .A(A[31]), .B(B[31]), .Y(n296) );
  OR2X2 U291 ( .A(A[25]), .B(B[25]), .Y(n384) );
  BUFX2 U292 ( .A(n115), .Y(n297) );
  INVX1 U293 ( .A(n114), .Y(n298) );
  INVX1 U294 ( .A(n82), .Y(n299) );
  INVX1 U295 ( .A(n42), .Y(n300) );
  INVX1 U296 ( .A(n34), .Y(n301) );
  BUFX2 U297 ( .A(n92), .Y(n302) );
  BUFX2 U298 ( .A(n36), .Y(n303) );
  BUFX2 U299 ( .A(n60), .Y(n304) );
  BUFX2 U300 ( .A(n52), .Y(n305) );
  BUFX2 U301 ( .A(n44), .Y(n306) );
  BUFX2 U302 ( .A(n125), .Y(n307) );
  BUFX2 U303 ( .A(n120), .Y(n308) );
  AND2X1 U304 ( .A(n327), .B(n170), .Y(n27) );
  INVX1 U305 ( .A(n27), .Y(n309) );
  INVX1 U306 ( .A(n24), .Y(n310) );
  AND2X1 U307 ( .A(n394), .B(n137), .Y(n26) );
  INVX1 U308 ( .A(n26), .Y(n311) );
  AND2X1 U309 ( .A(n328), .B(n123), .Y(n23) );
  INVX1 U310 ( .A(n23), .Y(n312) );
  INVX1 U311 ( .A(n22), .Y(n313) );
  AND2X1 U312 ( .A(n329), .B(n106), .Y(n20) );
  INVX1 U313 ( .A(n20), .Y(n314) );
  AND2X1 U314 ( .A(n330), .B(n98), .Y(n18) );
  INVX1 U315 ( .A(n18), .Y(n315) );
  AND2X1 U316 ( .A(n331), .B(n90), .Y(n16) );
  INVX1 U317 ( .A(n16), .Y(n316) );
  AND2X1 U318 ( .A(n332), .B(n82), .Y(n14) );
  INVX1 U319 ( .A(n14), .Y(n317) );
  AND2X1 U320 ( .A(n333), .B(n74), .Y(n12) );
  INVX1 U321 ( .A(n12), .Y(n318) );
  AND2X1 U322 ( .A(n334), .B(n58), .Y(n8) );
  INVX1 U323 ( .A(n8), .Y(n319) );
  AND2X1 U324 ( .A(n335), .B(n50), .Y(n6) );
  INVX1 U325 ( .A(n6), .Y(n320) );
  AND2X1 U326 ( .A(n336), .B(n42), .Y(n4) );
  INVX1 U327 ( .A(n4), .Y(n321) );
  AND2X1 U328 ( .A(n337), .B(n34), .Y(n2) );
  INVX1 U329 ( .A(n2), .Y(n322) );
  INVX1 U330 ( .A(n112), .Y(n323) );
  INVX1 U331 ( .A(n48), .Y(n324) );
  INVX1 U332 ( .A(n119), .Y(n325) );
  INVX1 U333 ( .A(n128), .Y(n326) );
  INVX1 U334 ( .A(n142), .Y(n327) );
  INVX1 U335 ( .A(n124), .Y(n328) );
  INVX1 U336 ( .A(n107), .Y(n329) );
  INVX1 U337 ( .A(n99), .Y(n330) );
  INVX1 U338 ( .A(n91), .Y(n331) );
  AND2X1 U339 ( .A(B[14]), .B(A[14]), .Y(n83) );
  INVX1 U340 ( .A(n83), .Y(n332) );
  INVX1 U341 ( .A(n75), .Y(n333) );
  AND2X1 U342 ( .A(B[20]), .B(A[20]), .Y(n59) );
  INVX1 U343 ( .A(n59), .Y(n334) );
  INVX1 U344 ( .A(n51), .Y(n335) );
  INVX1 U345 ( .A(n43), .Y(n336) );
  INVX1 U346 ( .A(n35), .Y(n337) );
  INVX1 U347 ( .A(n106), .Y(n338) );
  INVX1 U348 ( .A(n98), .Y(n339) );
  INVX1 U349 ( .A(n90), .Y(n340) );
  INVX1 U350 ( .A(n74), .Y(n341) );
  INVX1 U351 ( .A(n58), .Y(n342) );
  OR2X1 U352 ( .A(A[20]), .B(B[20]), .Y(n58) );
  INVX1 U353 ( .A(n50), .Y(n343) );
  INVX1 U354 ( .A(n121), .Y(n345) );
  INVX1 U355 ( .A(n84), .Y(n346) );
  INVX1 U356 ( .A(n346), .Y(n347) );
  INVX1 U357 ( .A(n76), .Y(n348) );
  INVX1 U358 ( .A(n348), .Y(n349) );
  BUFX2 U359 ( .A(n303), .Y(n350) );
  INVX1 U360 ( .A(n129), .Y(n351) );
  INVX1 U361 ( .A(n123), .Y(n352) );
  OR2X2 U362 ( .A(A[9]), .B(B[9]), .Y(n383) );
  INVX1 U363 ( .A(n135), .Y(n353) );
  INVX1 U364 ( .A(n138), .Y(n354) );
  OR2X2 U365 ( .A(B[0]), .B(A[0]), .Y(n393) );
  INVX1 U366 ( .A(n25), .Y(n355) );
  INVX1 U367 ( .A(n21), .Y(n356) );
  OR2X2 U368 ( .A(A[7]), .B(B[7]), .Y(n389) );
  INVX1 U369 ( .A(n40), .Y(n357) );
  INVX1 U370 ( .A(n67), .Y(n358) );
  BUFX2 U371 ( .A(n100), .Y(n359) );
  INVX1 U372 ( .A(n5), .Y(n360) );
  INVX1 U373 ( .A(n3), .Y(n361) );
  INVX1 U374 ( .A(n10), .Y(n362) );
  INVX1 U375 ( .A(n104), .Y(n363) );
  INVX1 U376 ( .A(n96), .Y(n364) );
  INVX1 U377 ( .A(n80), .Y(n365) );
  INVX1 U378 ( .A(n88), .Y(n366) );
  INVX1 U379 ( .A(n56), .Y(n367) );
  INVX1 U380 ( .A(n72), .Y(n368) );
  INVX1 U381 ( .A(n64), .Y(n369) );
  BUFX2 U382 ( .A(n108), .Y(n370) );
  INVX1 U383 ( .A(n134), .Y(n371) );
  INVX1 U384 ( .A(n19), .Y(n372) );
  INVX1 U385 ( .A(n17), .Y(n373) );
  INVX1 U386 ( .A(n15), .Y(n374) );
  INVX1 U387 ( .A(n13), .Y(n375) );
  INVX1 U388 ( .A(n11), .Y(n376) );
  INVX1 U389 ( .A(n9), .Y(n377) );
  INVX1 U390 ( .A(n7), .Y(n378) );
  OR2X1 U391 ( .A(A[18]), .B(B[18]), .Y(n66) );
  INVX1 U392 ( .A(n66), .Y(n379) );
  BUFX2 U393 ( .A(n131), .Y(n380) );
  INVX1 U394 ( .A(n132), .Y(n381) );
  OR2X2 U395 ( .A(A[17]), .B(B[17]), .Y(n392) );
  INVX1 U396 ( .A(n326), .Y(n167) );
  OR2X1 U397 ( .A(A[15]), .B(B[15]), .Y(n386) );
  BUFX2 U398 ( .A(n354), .Y(n394) );
  INVX1 U399 ( .A(n344), .Y(n170) );
  INVX1 U400 ( .A(n140), .Y(n139) );
  INVX1 U401 ( .A(n380), .Y(n130) );
  OAI21X1 U402 ( .A(n380), .B(n298), .C(n297), .Y(n395) );
  INVX1 U403 ( .A(n68), .Y(n396) );
  OAI21X1 U404 ( .A(n379), .B(n397), .C(n358), .Y(n398) );
endmodule


module alu_DW01_add_17 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n29, n30, n31,
         n32, n33, n34, n35, n36, n40, n41, n42, n43, n44, n48, n49, n50, n51,
         n52, n56, n57, n58, n59, n60, n64, n65, n66, n67, n68, n72, n73, n74,
         n75, n76, n80, n81, n82, n83, n84, n88, n89, n90, n91, n92, n96, n97,
         n98, n99, n100, n104, n105, n106, n107, n108, n112, n113, n114, n115,
         n119, n120, n121, n122, n123, n124, n125, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n144, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399;

  FAX1 U3 ( .A(B[30]), .B(A[30]), .C(n30), .YC(n29), .YS(SUM[30]) );
  FAX1 U4 ( .A(B[29]), .B(A[29]), .C(n31), .YC(n30), .YS(SUM[29]) );
  FAX1 U5 ( .A(B[28]), .B(A[28]), .C(n32), .YC(n31), .YS(SUM[28]) );
  FAX1 U6 ( .A(B[27]), .B(A[27]), .C(n33), .YC(n32), .YS(SUM[27]) );
  XOR2X1 U7 ( .A(n336), .B(n308), .Y(SUM[26]) );
  OAI21X1 U8 ( .A(n324), .B(n337), .C(n319), .Y(n33) );
  XNOR2X1 U13 ( .A(n41), .B(n378), .Y(SUM[25]) );
  AOI21X1 U14 ( .A(n41), .B(n386), .C(n40), .Y(n36) );
  XOR2X1 U21 ( .A(n334), .B(n307), .Y(SUM[24]) );
  OAI21X1 U22 ( .A(n323), .B(n334), .C(n318), .Y(n41) );
  XNOR2X1 U27 ( .A(n279), .B(n377), .Y(SUM[23]) );
  AOI21X1 U28 ( .A(n49), .B(n392), .C(n48), .Y(n44) );
  XOR2X1 U35 ( .A(n332), .B(n306), .Y(SUM[22]) );
  OAI21X1 U36 ( .A(n322), .B(n332), .C(n317), .Y(n49) );
  XNOR2X1 U41 ( .A(n57), .B(n376), .Y(SUM[21]) );
  AOI21X1 U42 ( .A(n275), .B(n388), .C(n56), .Y(n52) );
  XOR2X1 U49 ( .A(n330), .B(n305), .Y(SUM[20]) );
  OAI21X1 U50 ( .A(n291), .B(n293), .C(n316), .Y(n57) );
  XNOR2X1 U55 ( .A(n274), .B(n375), .Y(SUM[19]) );
  AOI21X1 U56 ( .A(n65), .B(n384), .C(n64), .Y(n60) );
  XOR2X1 U63 ( .A(n284), .B(n304), .Y(SUM[18]) );
  OAI21X1 U64 ( .A(n290), .B(n329), .C(n315), .Y(n65) );
  XNOR2X1 U69 ( .A(n73), .B(n374), .Y(SUM[17]) );
  AOI21X1 U70 ( .A(n276), .B(n383), .C(n72), .Y(n68) );
  XOR2X1 U77 ( .A(n396), .B(n303), .Y(SUM[16]) );
  OAI21X1 U78 ( .A(n289), .B(n292), .C(n314), .Y(n73) );
  XNOR2X1 U83 ( .A(n286), .B(n373), .Y(SUM[15]) );
  AOI21X1 U84 ( .A(n81), .B(n387), .C(n80), .Y(n76) );
  XOR2X1 U91 ( .A(n285), .B(n352), .Y(SUM[14]) );
  OAI21X1 U92 ( .A(n369), .B(n397), .C(n348), .Y(n81) );
  XNOR2X1 U97 ( .A(n89), .B(n357), .Y(SUM[13]) );
  AOI21X1 U98 ( .A(n89), .B(n391), .C(n88), .Y(n84) );
  XOR2X1 U105 ( .A(n399), .B(n346), .Y(SUM[12]) );
  OAI21X1 U106 ( .A(n368), .B(n355), .C(n344), .Y(n89) );
  XNOR2X1 U111 ( .A(n97), .B(n372), .Y(SUM[11]) );
  AOI21X1 U112 ( .A(n277), .B(n390), .C(n96), .Y(n92) );
  XOR2X1 U119 ( .A(n398), .B(n351), .Y(SUM[10]) );
  OAI21X1 U120 ( .A(n367), .B(n398), .C(n347), .Y(n97) );
  XNOR2X1 U125 ( .A(n280), .B(n356), .Y(SUM[9]) );
  AOI21X1 U126 ( .A(n105), .B(n381), .C(n104), .Y(n100) );
  XOR2X1 U133 ( .A(n327), .B(n302), .Y(SUM[8]) );
  OAI21X1 U134 ( .A(n321), .B(n327), .C(n313), .Y(n105) );
  XNOR2X1 U139 ( .A(n278), .B(n371), .Y(SUM[7]) );
  AOI21X1 U140 ( .A(n113), .B(n389), .C(n112), .Y(n108) );
  XOR2X1 U147 ( .A(n298), .B(n301), .Y(SUM[6]) );
  OAI21X1 U148 ( .A(n294), .B(n288), .C(n296), .Y(n113) );
  AOI21X1 U150 ( .A(n122), .B(n382), .C(n119), .Y(n115) );
  XOR2X1 U157 ( .A(n297), .B(n300), .Y(SUM[5]) );
  AOI21X1 U158 ( .A(n130), .B(n325), .C(n122), .Y(n120) );
  OAI21X1 U160 ( .A(n338), .B(n340), .C(n312), .Y(n122) );
  XNOR2X1 U165 ( .A(n130), .B(n299), .Y(SUM[4]) );
  AOI21X1 U166 ( .A(n130), .B(n310), .C(n129), .Y(n125) );
  XNOR2X1 U173 ( .A(n136), .B(n350), .Y(SUM[3]) );
  AOI21X1 U175 ( .A(n287), .B(n140), .C(n133), .Y(n131) );
  OAI21X1 U177 ( .A(n320), .B(n370), .C(n349), .Y(n133) );
  XOR2X1 U182 ( .A(n139), .B(n358), .Y(SUM[2]) );
  OAI21X1 U183 ( .A(n379), .B(n139), .C(n395), .Y(n136) );
  XOR2X1 U188 ( .A(n343), .B(n380), .Y(SUM[1]) );
  OAI21X1 U190 ( .A(n380), .B(n345), .C(n342), .Y(n140) );
  BUFX2 U203 ( .A(n65), .Y(n274) );
  AND2X2 U204 ( .A(B[16]), .B(A[16]), .Y(n75) );
  OR2X2 U205 ( .A(A[16]), .B(B[16]), .Y(n74) );
  AND2X1 U206 ( .A(n382), .B(n325), .Y(n114) );
  OR2X1 U207 ( .A(A[9]), .B(B[9]), .Y(n381) );
  OR2X1 U208 ( .A(n370), .B(n379), .Y(n132) );
  AND2X1 U209 ( .A(A[2]), .B(B[2]), .Y(n138) );
  AND2X1 U210 ( .A(B[14]), .B(A[14]), .Y(n83) );
  AND2X1 U211 ( .A(B[10]), .B(A[10]), .Y(n99) );
  OR2X1 U212 ( .A(n341), .B(n311), .Y(n121) );
  AND2X1 U213 ( .A(A[5]), .B(B[5]), .Y(n124) );
  AND2X1 U214 ( .A(A[3]), .B(B[3]), .Y(n135) );
  INVX1 U215 ( .A(n141), .Y(n345) );
  OR2X1 U216 ( .A(B[1]), .B(A[1]), .Y(n141) );
  AND2X1 U217 ( .A(A[1]), .B(B[1]), .Y(n142) );
  AND2X1 U218 ( .A(n364), .B(n386), .Y(n3) );
  INVX1 U219 ( .A(n333), .Y(n334) );
  AND2X1 U220 ( .A(n363), .B(n392), .Y(n5) );
  INVX1 U221 ( .A(n331), .Y(n332) );
  AND2X1 U222 ( .A(n362), .B(n388), .Y(n7) );
  AND2X1 U223 ( .A(n361), .B(n384), .Y(n9) );
  AND2X1 U224 ( .A(n360), .B(n383), .Y(n11) );
  AND2X1 U225 ( .A(n366), .B(n387), .Y(n13) );
  AND2X1 U226 ( .A(n348), .B(n82), .Y(n14) );
  AND2X1 U227 ( .A(n354), .B(n391), .Y(n15) );
  AND2X1 U228 ( .A(n344), .B(n90), .Y(n16) );
  AND2X1 U229 ( .A(n365), .B(n390), .Y(n17) );
  AND2X1 U230 ( .A(n347), .B(n98), .Y(n18) );
  AND2X1 U231 ( .A(n353), .B(n381), .Y(n19) );
  INVX1 U232 ( .A(n326), .Y(n327) );
  AND2X1 U233 ( .A(n359), .B(n389), .Y(n21) );
  AND2X1 U234 ( .A(n349), .B(n134), .Y(n25) );
  AND2X1 U235 ( .A(n342), .B(n141), .Y(n27) );
  AND2X1 U236 ( .A(A[0]), .B(B[0]), .Y(n144) );
  OAI21X1 U237 ( .A(n291), .B(n293), .C(n316), .Y(n275) );
  OAI21X1 U238 ( .A(n289), .B(n292), .C(n314), .Y(n276) );
  OAI21X1 U239 ( .A(n367), .B(n398), .C(n347), .Y(n277) );
  BUFX2 U240 ( .A(n113), .Y(n278) );
  INVX1 U241 ( .A(n144), .Y(n380) );
  AND2X1 U242 ( .A(B[21]), .B(A[21]), .Y(n56) );
  OR2X1 U243 ( .A(A[5]), .B(B[5]), .Y(n123) );
  AND2X1 U244 ( .A(B[9]), .B(A[9]), .Y(n104) );
  AND2X1 U245 ( .A(B[17]), .B(A[17]), .Y(n72) );
  AND2X1 U246 ( .A(A[4]), .B(B[4]), .Y(n129) );
  OR2X1 U247 ( .A(A[20]), .B(B[20]), .Y(n58) );
  INVX1 U248 ( .A(n137), .Y(n379) );
  OR2X1 U249 ( .A(A[2]), .B(B[2]), .Y(n137) );
  OR2X1 U250 ( .A(A[3]), .B(B[3]), .Y(n134) );
  BUFX2 U251 ( .A(n49), .Y(n279) );
  BUFX2 U252 ( .A(n105), .Y(n280) );
  OR2X2 U253 ( .A(A[17]), .B(B[17]), .Y(n383) );
  BUFX2 U254 ( .A(n311), .Y(n281) );
  OR2X1 U255 ( .A(B[4]), .B(A[4]), .Y(n128) );
  OAI21X1 U256 ( .A(n380), .B(n345), .C(n342), .Y(n282) );
  INVX1 U257 ( .A(n337), .Y(n283) );
  OR2X1 U258 ( .A(A[6]), .B(B[6]), .Y(n382) );
  BUFX2 U259 ( .A(n329), .Y(n284) );
  BUFX2 U260 ( .A(n397), .Y(n285) );
  OAI21X1 U261 ( .A(n369), .B(n285), .C(n348), .Y(n286) );
  AND2X2 U262 ( .A(B[20]), .B(A[20]), .Y(n59) );
  OR2X2 U263 ( .A(A[21]), .B(B[21]), .Y(n388) );
  INVX1 U264 ( .A(n132), .Y(n287) );
  INVX1 U265 ( .A(n114), .Y(n288) );
  INVX1 U266 ( .A(n74), .Y(n289) );
  OR2X1 U267 ( .A(A[18]), .B(B[18]), .Y(n66) );
  INVX1 U268 ( .A(n66), .Y(n290) );
  INVX1 U269 ( .A(n58), .Y(n291) );
  BUFX2 U270 ( .A(n76), .Y(n292) );
  BUFX2 U271 ( .A(n60), .Y(n293) );
  BUFX2 U272 ( .A(n131), .Y(n294) );
  INVX1 U273 ( .A(n115), .Y(n295) );
  INVX1 U274 ( .A(n295), .Y(n296) );
  BUFX2 U275 ( .A(n125), .Y(n297) );
  BUFX2 U276 ( .A(n120), .Y(n298) );
  AND2X1 U277 ( .A(n338), .B(n310), .Y(n24) );
  INVX1 U278 ( .A(n24), .Y(n299) );
  AND2X1 U279 ( .A(n312), .B(n339), .Y(n23) );
  INVX1 U280 ( .A(n23), .Y(n300) );
  AND2X1 U281 ( .A(n309), .B(n382), .Y(n22) );
  INVX1 U282 ( .A(n22), .Y(n301) );
  AND2X1 U283 ( .A(n313), .B(n106), .Y(n20) );
  INVX1 U284 ( .A(n20), .Y(n302) );
  AND2X1 U285 ( .A(n314), .B(n74), .Y(n12) );
  INVX1 U286 ( .A(n12), .Y(n303) );
  AND2X1 U287 ( .A(n315), .B(n66), .Y(n10) );
  INVX1 U288 ( .A(n10), .Y(n304) );
  AND2X1 U289 ( .A(n316), .B(n58), .Y(n8) );
  INVX1 U290 ( .A(n8), .Y(n305) );
  AND2X1 U291 ( .A(n317), .B(n50), .Y(n6) );
  INVX1 U292 ( .A(n6), .Y(n306) );
  AND2X1 U293 ( .A(n318), .B(n42), .Y(n4) );
  INVX1 U294 ( .A(n4), .Y(n307) );
  AND2X1 U295 ( .A(n319), .B(n34), .Y(n2) );
  INVX1 U296 ( .A(n2), .Y(n308) );
  AND2X1 U297 ( .A(B[6]), .B(A[6]), .Y(n119) );
  INVX1 U298 ( .A(n119), .Y(n309) );
  INVX1 U299 ( .A(n281), .Y(n310) );
  INVX1 U300 ( .A(n128), .Y(n311) );
  INVX1 U301 ( .A(n124), .Y(n312) );
  AND2X1 U302 ( .A(B[8]), .B(A[8]), .Y(n107) );
  INVX1 U303 ( .A(n107), .Y(n313) );
  INVX1 U304 ( .A(n75), .Y(n314) );
  AND2X1 U305 ( .A(B[18]), .B(A[18]), .Y(n67) );
  INVX1 U306 ( .A(n67), .Y(n315) );
  INVX1 U307 ( .A(n59), .Y(n316) );
  AND2X1 U308 ( .A(B[22]), .B(A[22]), .Y(n51) );
  INVX1 U309 ( .A(n51), .Y(n317) );
  AND2X1 U310 ( .A(B[24]), .B(A[24]), .Y(n43) );
  INVX1 U311 ( .A(n43), .Y(n318) );
  AND2X1 U312 ( .A(B[26]), .B(A[26]), .Y(n35) );
  INVX1 U313 ( .A(n35), .Y(n319) );
  INVX1 U314 ( .A(n138), .Y(n320) );
  OR2X1 U315 ( .A(A[8]), .B(B[8]), .Y(n106) );
  INVX1 U316 ( .A(n106), .Y(n321) );
  OR2X1 U317 ( .A(A[22]), .B(B[22]), .Y(n50) );
  INVX1 U318 ( .A(n50), .Y(n322) );
  OR2X1 U319 ( .A(A[24]), .B(B[24]), .Y(n42) );
  INVX1 U320 ( .A(n42), .Y(n323) );
  OR2X1 U321 ( .A(A[26]), .B(B[26]), .Y(n34) );
  INVX1 U322 ( .A(n34), .Y(n324) );
  INVX1 U323 ( .A(n121), .Y(n325) );
  INVX1 U324 ( .A(n108), .Y(n326) );
  INVX1 U325 ( .A(n68), .Y(n328) );
  INVX1 U326 ( .A(n328), .Y(n329) );
  BUFX2 U327 ( .A(n293), .Y(n330) );
  INVX1 U328 ( .A(n52), .Y(n331) );
  INVX1 U329 ( .A(n44), .Y(n333) );
  INVX1 U330 ( .A(n36), .Y(n335) );
  INVX1 U331 ( .A(n283), .Y(n336) );
  INVX1 U332 ( .A(n335), .Y(n337) );
  INVX1 U333 ( .A(n129), .Y(n338) );
  INVX1 U334 ( .A(n341), .Y(n339) );
  INVX1 U335 ( .A(n339), .Y(n340) );
  INVX1 U336 ( .A(n123), .Y(n341) );
  INVX1 U337 ( .A(n142), .Y(n342) );
  INVX1 U338 ( .A(n27), .Y(n343) );
  AND2X1 U339 ( .A(B[12]), .B(A[12]), .Y(n91) );
  INVX1 U340 ( .A(n91), .Y(n344) );
  INVX1 U341 ( .A(n16), .Y(n346) );
  INVX1 U342 ( .A(n99), .Y(n347) );
  INVX1 U343 ( .A(n83), .Y(n348) );
  INVX1 U344 ( .A(n135), .Y(n349) );
  AND2X1 U345 ( .A(n380), .B(n385), .Y(SUM[0]) );
  INVX1 U346 ( .A(n25), .Y(n350) );
  INVX1 U347 ( .A(n18), .Y(n351) );
  INVX1 U348 ( .A(n14), .Y(n352) );
  INVX1 U349 ( .A(n104), .Y(n353) );
  AND2X1 U350 ( .A(B[13]), .B(A[13]), .Y(n88) );
  INVX1 U351 ( .A(n88), .Y(n354) );
  BUFX2 U352 ( .A(n92), .Y(n355) );
  INVX1 U353 ( .A(n19), .Y(n356) );
  INVX1 U354 ( .A(n15), .Y(n357) );
  AND2X1 U355 ( .A(n395), .B(n137), .Y(n26) );
  INVX1 U356 ( .A(n26), .Y(n358) );
  AND2X1 U357 ( .A(B[7]), .B(A[7]), .Y(n112) );
  INVX1 U358 ( .A(n112), .Y(n359) );
  INVX1 U359 ( .A(n72), .Y(n360) );
  AND2X1 U360 ( .A(B[19]), .B(A[19]), .Y(n64) );
  INVX1 U361 ( .A(n64), .Y(n361) );
  INVX1 U362 ( .A(n56), .Y(n362) );
  AND2X1 U363 ( .A(B[23]), .B(A[23]), .Y(n48) );
  INVX1 U364 ( .A(n48), .Y(n363) );
  AND2X1 U365 ( .A(B[25]), .B(A[25]), .Y(n40) );
  INVX1 U366 ( .A(n40), .Y(n364) );
  AND2X1 U367 ( .A(B[11]), .B(A[11]), .Y(n96) );
  INVX1 U368 ( .A(n96), .Y(n365) );
  AND2X1 U369 ( .A(B[15]), .B(A[15]), .Y(n80) );
  INVX1 U370 ( .A(n80), .Y(n366) );
  OR2X1 U371 ( .A(A[10]), .B(B[10]), .Y(n98) );
  INVX1 U372 ( .A(n98), .Y(n367) );
  OR2X1 U373 ( .A(A[12]), .B(B[12]), .Y(n90) );
  INVX1 U374 ( .A(n90), .Y(n368) );
  OR2X1 U375 ( .A(A[14]), .B(B[14]), .Y(n82) );
  INVX1 U376 ( .A(n82), .Y(n369) );
  INVX1 U377 ( .A(n134), .Y(n370) );
  INVX1 U378 ( .A(n21), .Y(n371) );
  INVX1 U379 ( .A(n17), .Y(n372) );
  INVX1 U380 ( .A(n13), .Y(n373) );
  INVX1 U381 ( .A(n11), .Y(n374) );
  INVX1 U382 ( .A(n9), .Y(n375) );
  INVX1 U383 ( .A(n7), .Y(n376) );
  INVX1 U384 ( .A(n5), .Y(n377) );
  INVX1 U385 ( .A(n3), .Y(n378) );
  OR2X1 U386 ( .A(A[19]), .B(B[19]), .Y(n384) );
  OR2X1 U387 ( .A(B[0]), .B(A[0]), .Y(n385) );
  OR2X1 U388 ( .A(A[25]), .B(B[25]), .Y(n386) );
  OR2X1 U389 ( .A(A[15]), .B(B[15]), .Y(n387) );
  OR2X1 U390 ( .A(A[7]), .B(B[7]), .Y(n389) );
  OR2X1 U391 ( .A(A[11]), .B(B[11]), .Y(n390) );
  OR2X1 U392 ( .A(A[13]), .B(B[13]), .Y(n391) );
  OR2X1 U393 ( .A(A[23]), .B(B[23]), .Y(n392) );
  INVX1 U394 ( .A(n294), .Y(n130) );
  INVX1 U395 ( .A(n282), .Y(n139) );
  XNOR2X1 U396 ( .A(n29), .B(n393), .Y(SUM[31]) );
  XNOR2X1 U397 ( .A(A[31]), .B(B[31]), .Y(n393) );
  INVX1 U398 ( .A(n320), .Y(n394) );
  INVX1 U399 ( .A(n394), .Y(n395) );
  BUFX2 U400 ( .A(n292), .Y(n396) );
  BUFX2 U401 ( .A(n84), .Y(n397) );
  BUFX2 U402 ( .A(n100), .Y(n398) );
  BUFX2 U403 ( .A(n355), .Y(n399) );
endmodule


module alu_DW01_sub_16 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n39, n40, n41, n42, n43, n47, n48, n49, n50,
         n51, n55, n56, n57, n58, n59, n63, n64, n65, n66, n67, n71, n72, n73,
         n74, n75, n79, n80, n81, n82, n83, n87, n88, n89, n90, n91, n95, n96,
         n97, n98, n99, n103, n104, n105, n106, n107, n111, n112, n113, n114,
         n118, n119, n120, n121, n122, n123, n124, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n165, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460;

  XOR2X1 U1 ( .A(n28), .B(n1), .Y(DIFF[31]) );
  FAX1 U3 ( .A(n460), .B(A[30]), .C(n29), .YC(n28), .YS(DIFF[30]) );
  FAX1 U4 ( .A(n459), .B(A[29]), .C(n30), .YC(n29), .YS(DIFF[29]) );
  FAX1 U5 ( .A(n458), .B(A[28]), .C(n31), .YC(n30), .YS(DIFF[28]) );
  FAX1 U6 ( .A(n457), .B(A[27]), .C(n32), .YC(n31), .YS(DIFF[27]) );
  OAI21X1 U8 ( .A(n377), .B(n330), .C(n372), .Y(n32) );
  XNOR2X1 U13 ( .A(n307), .B(n341), .Y(DIFF[25]) );
  AOI21X1 U14 ( .A(n40), .B(n427), .C(n39), .Y(n35) );
  XOR2X1 U21 ( .A(n398), .B(n352), .Y(DIFF[24]) );
  OAI21X1 U22 ( .A(n326), .B(n329), .C(n371), .Y(n40) );
  XNOR2X1 U27 ( .A(n304), .B(n340), .Y(DIFF[23]) );
  AOI21X1 U28 ( .A(n48), .B(n419), .C(n47), .Y(n43) );
  XOR2X1 U35 ( .A(n315), .B(n351), .Y(DIFF[22]) );
  OAI21X1 U36 ( .A(n331), .B(n397), .C(n370), .Y(n48) );
  XNOR2X1 U41 ( .A(n309), .B(n339), .Y(DIFF[21]) );
  AOI21X1 U42 ( .A(n56), .B(n421), .C(n55), .Y(n51) );
  XOR2X1 U49 ( .A(n394), .B(n350), .Y(DIFF[20]) );
  OAI21X1 U50 ( .A(n376), .B(n395), .C(n369), .Y(n56) );
  XNOR2X1 U55 ( .A(n314), .B(n338), .Y(DIFF[19]) );
  AOI21X1 U56 ( .A(n64), .B(n426), .C(n63), .Y(n59) );
  XOR2X1 U63 ( .A(n392), .B(n349), .Y(DIFF[18]) );
  OAI21X1 U64 ( .A(n325), .B(n328), .C(n368), .Y(n64) );
  XNOR2X1 U69 ( .A(n305), .B(n337), .Y(DIFF[17]) );
  AOI21X1 U70 ( .A(n72), .B(n428), .C(n71), .Y(n67) );
  XOR2X1 U77 ( .A(n390), .B(n348), .Y(DIFF[16]) );
  OAI21X1 U78 ( .A(n375), .B(n391), .C(n367), .Y(n72) );
  XNOR2X1 U83 ( .A(n310), .B(n336), .Y(DIFF[15]) );
  AOI21X1 U84 ( .A(n80), .B(n420), .C(n79), .Y(n75) );
  XOR2X1 U91 ( .A(n387), .B(n347), .Y(DIFF[14]) );
  OAI21X1 U92 ( .A(n374), .B(n388), .C(n366), .Y(n80) );
  XNOR2X1 U97 ( .A(n311), .B(n335), .Y(DIFF[13]) );
  AOI21X1 U98 ( .A(n88), .B(n424), .C(n87), .Y(n83) );
  XOR2X1 U105 ( .A(n385), .B(n346), .Y(DIFF[12]) );
  OAI21X1 U106 ( .A(n324), .B(n327), .C(n365), .Y(n88) );
  XNOR2X1 U111 ( .A(n306), .B(n334), .Y(DIFF[11]) );
  AOI21X1 U112 ( .A(n96), .B(n423), .C(n95), .Y(n91) );
  XOR2X1 U119 ( .A(n383), .B(n345), .Y(DIFF[10]) );
  OAI21X1 U120 ( .A(n373), .B(n384), .C(n364), .Y(n96) );
  XNOR2X1 U125 ( .A(n312), .B(n333), .Y(DIFF[9]) );
  AOI21X1 U126 ( .A(n104), .B(n425), .C(n103), .Y(n99) );
  XOR2X1 U133 ( .A(n380), .B(n344), .Y(DIFF[8]) );
  OAI21X1 U134 ( .A(n323), .B(n381), .C(n363), .Y(n104) );
  XNOR2X1 U139 ( .A(n313), .B(n414), .Y(DIFF[7]) );
  AOI21X1 U140 ( .A(n112), .B(n422), .C(n111), .Y(n107) );
  XOR2X1 U147 ( .A(n332), .B(n343), .Y(DIFF[6]) );
  OAI21X1 U148 ( .A(n322), .B(n405), .C(n321), .Y(n112) );
  AOI21X1 U150 ( .A(n121), .B(n418), .C(n118), .Y(n114) );
  XOR2X1 U157 ( .A(n403), .B(n402), .Y(DIFF[5]) );
  AOI21X1 U158 ( .A(n129), .B(n378), .C(n121), .Y(n119) );
  OAI21X1 U160 ( .A(n412), .B(n417), .C(n407), .Y(n121) );
  XNOR2X1 U165 ( .A(n129), .B(n399), .Y(DIFF[4]) );
  AOI21X1 U166 ( .A(n129), .B(n165), .C(n128), .Y(n124) );
  XNOR2X1 U173 ( .A(n135), .B(n400), .Y(DIFF[3]) );
  AOI21X1 U175 ( .A(n406), .B(n303), .C(n132), .Y(n130) );
  OAI21X1 U177 ( .A(n413), .B(n316), .C(n362), .Y(n132) );
  XOR2X1 U182 ( .A(n138), .B(n401), .Y(DIFF[2]) );
  OAI21X1 U183 ( .A(n409), .B(n138), .C(n413), .Y(n135) );
  XOR2X1 U188 ( .A(n404), .B(n416), .Y(DIFF[1]) );
  OAI21X1 U190 ( .A(n416), .B(n411), .C(n408), .Y(n139) );
  XNOR2X1 U195 ( .A(n430), .B(A[0]), .Y(DIFF[0]) );
  OAI21X1 U232 ( .A(n416), .B(n411), .C(n408), .Y(n303) );
  OR2X2 U233 ( .A(A[5]), .B(n435), .Y(n122) );
  AND2X2 U234 ( .A(n435), .B(A[5]), .Y(n123) );
  OR2X1 U235 ( .A(n308), .B(n417), .Y(n120) );
  OR2X1 U236 ( .A(A[6]), .B(n436), .Y(n418) );
  AND2X1 U237 ( .A(n436), .B(A[6]), .Y(n118) );
  OR2X1 U238 ( .A(n409), .B(n316), .Y(n131) );
  OR2X1 U239 ( .A(A[25]), .B(n455), .Y(n427) );
  AND2X1 U240 ( .A(n454), .B(A[24]), .Y(n42) );
  AND2X1 U241 ( .A(n442), .B(A[12]), .Y(n90) );
  AND2X1 U242 ( .A(n440), .B(A[10]), .Y(n98) );
  AND2X1 U243 ( .A(n410), .B(n422), .Y(n21) );
  AND2X1 U244 ( .A(n412), .B(n165), .Y(n24) );
  AND2X1 U245 ( .A(n362), .B(n133), .Y(n25) );
  INVX1 U246 ( .A(n133), .Y(n316) );
  OR2X1 U247 ( .A(A[10]), .B(n440), .Y(n97) );
  OR2X1 U248 ( .A(A[12]), .B(n442), .Y(n89) );
  AND2X1 U249 ( .A(n455), .B(A[25]), .Y(n39) );
  INVX1 U250 ( .A(n128), .Y(n412) );
  OR2X1 U251 ( .A(A[8]), .B(n438), .Y(n105) );
  OR2X1 U252 ( .A(A[24]), .B(n454), .Y(n41) );
  OR2X1 U253 ( .A(A[3]), .B(n433), .Y(n133) );
  BUFX2 U254 ( .A(n48), .Y(n304) );
  BUFX2 U255 ( .A(n72), .Y(n305) );
  BUFX2 U256 ( .A(n96), .Y(n306) );
  OAI21X1 U257 ( .A(n326), .B(n329), .C(n371), .Y(n307) );
  INVX1 U258 ( .A(n127), .Y(n308) );
  BUFX2 U259 ( .A(n56), .Y(n309) );
  BUFX2 U260 ( .A(n80), .Y(n310) );
  OAI21X1 U261 ( .A(n324), .B(n327), .C(n365), .Y(n311) );
  BUFX2 U262 ( .A(n104), .Y(n312) );
  BUFX2 U263 ( .A(n112), .Y(n313) );
  OAI21X1 U264 ( .A(n325), .B(n328), .C(n368), .Y(n314) );
  OR2X2 U265 ( .A(A[4]), .B(n434), .Y(n127) );
  INVX2 U266 ( .A(n142), .Y(n416) );
  BUFX2 U267 ( .A(n397), .Y(n315) );
  OR2X2 U268 ( .A(n430), .B(A[0]), .Y(n142) );
  INVX1 U269 ( .A(n388), .Y(n317) );
  BUFX2 U270 ( .A(n405), .Y(n318) );
  INVX1 U271 ( .A(n391), .Y(n319) );
  BUFX2 U272 ( .A(n330), .Y(n320) );
  INVX1 U273 ( .A(n137), .Y(n413) );
  BUFX2 U274 ( .A(n114), .Y(n321) );
  AND2X2 U275 ( .A(n418), .B(n378), .Y(n113) );
  INVX1 U276 ( .A(n113), .Y(n322) );
  INVX1 U277 ( .A(n105), .Y(n323) );
  INVX1 U278 ( .A(n89), .Y(n324) );
  OR2X1 U279 ( .A(n448), .B(A[18]), .Y(n65) );
  INVX1 U280 ( .A(n65), .Y(n325) );
  INVX1 U281 ( .A(n41), .Y(n326) );
  BUFX2 U282 ( .A(n91), .Y(n327) );
  BUFX2 U283 ( .A(n67), .Y(n328) );
  BUFX2 U284 ( .A(n43), .Y(n329) );
  BUFX2 U285 ( .A(n35), .Y(n330) );
  OR2X1 U286 ( .A(A[22]), .B(n452), .Y(n49) );
  INVX1 U287 ( .A(n49), .Y(n331) );
  BUFX2 U288 ( .A(n119), .Y(n332) );
  AND2X1 U289 ( .A(n354), .B(n425), .Y(n19) );
  INVX1 U290 ( .A(n19), .Y(n333) );
  AND2X1 U291 ( .A(n355), .B(n423), .Y(n17) );
  INVX1 U292 ( .A(n17), .Y(n334) );
  AND2X1 U293 ( .A(n356), .B(n424), .Y(n15) );
  INVX1 U294 ( .A(n15), .Y(n335) );
  AND2X1 U295 ( .A(n357), .B(n420), .Y(n13) );
  INVX1 U296 ( .A(n13), .Y(n336) );
  AND2X1 U297 ( .A(n358), .B(n428), .Y(n11) );
  INVX1 U298 ( .A(n11), .Y(n337) );
  AND2X1 U299 ( .A(n359), .B(n426), .Y(n9) );
  INVX1 U300 ( .A(n9), .Y(n338) );
  AND2X1 U301 ( .A(n360), .B(n421), .Y(n7) );
  INVX1 U302 ( .A(n7), .Y(n339) );
  AND2X1 U303 ( .A(n361), .B(n419), .Y(n5) );
  INVX1 U304 ( .A(n5), .Y(n340) );
  AND2X1 U305 ( .A(n415), .B(n427), .Y(n3) );
  INVX1 U306 ( .A(n3), .Y(n341) );
  AND2X1 U307 ( .A(n372), .B(n33), .Y(n2) );
  INVX1 U308 ( .A(n2), .Y(n342) );
  AND2X1 U309 ( .A(n353), .B(n418), .Y(n22) );
  INVX1 U310 ( .A(n22), .Y(n343) );
  AND2X1 U311 ( .A(n363), .B(n105), .Y(n20) );
  INVX1 U312 ( .A(n20), .Y(n344) );
  AND2X1 U313 ( .A(n364), .B(n97), .Y(n18) );
  INVX1 U314 ( .A(n18), .Y(n345) );
  AND2X1 U315 ( .A(n365), .B(n89), .Y(n16) );
  INVX1 U316 ( .A(n16), .Y(n346) );
  AND2X1 U317 ( .A(n366), .B(n81), .Y(n14) );
  INVX1 U318 ( .A(n14), .Y(n347) );
  AND2X1 U319 ( .A(n367), .B(n73), .Y(n12) );
  INVX1 U320 ( .A(n12), .Y(n348) );
  AND2X1 U321 ( .A(n368), .B(n65), .Y(n10) );
  INVX1 U322 ( .A(n10), .Y(n349) );
  AND2X1 U323 ( .A(n369), .B(n57), .Y(n8) );
  INVX1 U324 ( .A(n8), .Y(n350) );
  AND2X1 U325 ( .A(n370), .B(n49), .Y(n6) );
  INVX1 U326 ( .A(n6), .Y(n351) );
  AND2X1 U327 ( .A(n371), .B(n41), .Y(n4) );
  INVX1 U328 ( .A(n4), .Y(n352) );
  INVX1 U329 ( .A(n118), .Y(n353) );
  AND2X1 U330 ( .A(n439), .B(A[9]), .Y(n103) );
  INVX1 U331 ( .A(n103), .Y(n354) );
  AND2X1 U332 ( .A(n441), .B(A[11]), .Y(n95) );
  INVX1 U333 ( .A(n95), .Y(n355) );
  AND2X1 U334 ( .A(n443), .B(A[13]), .Y(n87) );
  INVX1 U335 ( .A(n87), .Y(n356) );
  AND2X1 U336 ( .A(n445), .B(A[15]), .Y(n79) );
  INVX1 U337 ( .A(n79), .Y(n357) );
  AND2X1 U338 ( .A(n447), .B(A[17]), .Y(n71) );
  INVX1 U339 ( .A(n71), .Y(n358) );
  AND2X1 U340 ( .A(n449), .B(A[19]), .Y(n63) );
  INVX1 U341 ( .A(n63), .Y(n359) );
  AND2X1 U342 ( .A(n451), .B(A[21]), .Y(n55) );
  INVX1 U343 ( .A(n55), .Y(n360) );
  AND2X1 U344 ( .A(n453), .B(A[23]), .Y(n47) );
  INVX1 U345 ( .A(n47), .Y(n361) );
  AND2X1 U346 ( .A(A[3]), .B(n433), .Y(n134) );
  INVX1 U347 ( .A(n134), .Y(n362) );
  AND2X1 U348 ( .A(n438), .B(A[8]), .Y(n106) );
  INVX1 U349 ( .A(n106), .Y(n363) );
  INVX1 U350 ( .A(n98), .Y(n364) );
  INVX1 U351 ( .A(n90), .Y(n365) );
  AND2X1 U352 ( .A(n444), .B(A[14]), .Y(n82) );
  INVX1 U353 ( .A(n82), .Y(n366) );
  AND2X1 U354 ( .A(A[16]), .B(n446), .Y(n74) );
  INVX1 U355 ( .A(n74), .Y(n367) );
  AND2X1 U356 ( .A(A[18]), .B(n448), .Y(n66) );
  INVX1 U357 ( .A(n66), .Y(n368) );
  AND2X1 U358 ( .A(n450), .B(A[20]), .Y(n58) );
  INVX1 U359 ( .A(n58), .Y(n369) );
  AND2X1 U360 ( .A(n452), .B(A[22]), .Y(n50) );
  INVX1 U361 ( .A(n50), .Y(n370) );
  INVX1 U362 ( .A(n42), .Y(n371) );
  AND2X1 U363 ( .A(n456), .B(A[26]), .Y(n34) );
  INVX1 U364 ( .A(n34), .Y(n372) );
  INVX1 U365 ( .A(n97), .Y(n373) );
  OR2X1 U366 ( .A(A[14]), .B(n444), .Y(n81) );
  INVX1 U367 ( .A(n81), .Y(n374) );
  OR2X1 U368 ( .A(n446), .B(A[16]), .Y(n73) );
  INVX1 U369 ( .A(n73), .Y(n375) );
  INVX1 U370 ( .A(n57), .Y(n376) );
  OR2X1 U371 ( .A(A[20]), .B(n450), .Y(n57) );
  OR2X1 U372 ( .A(A[26]), .B(n456), .Y(n33) );
  INVX1 U373 ( .A(n33), .Y(n377) );
  INVX1 U374 ( .A(n120), .Y(n378) );
  INVX1 U375 ( .A(n107), .Y(n379) );
  INVX1 U376 ( .A(n379), .Y(n380) );
  INVX1 U377 ( .A(n379), .Y(n381) );
  INVX1 U378 ( .A(n99), .Y(n382) );
  INVX1 U379 ( .A(n382), .Y(n383) );
  INVX1 U380 ( .A(n382), .Y(n384) );
  BUFX2 U381 ( .A(n327), .Y(n385) );
  INVX1 U382 ( .A(n83), .Y(n386) );
  INVX1 U383 ( .A(n317), .Y(n387) );
  INVX1 U384 ( .A(n386), .Y(n388) );
  INVX1 U385 ( .A(n75), .Y(n389) );
  INVX1 U386 ( .A(n319), .Y(n390) );
  INVX1 U387 ( .A(n389), .Y(n391) );
  BUFX2 U388 ( .A(n328), .Y(n392) );
  INVX1 U389 ( .A(n59), .Y(n393) );
  INVX1 U390 ( .A(n393), .Y(n394) );
  INVX1 U391 ( .A(n393), .Y(n395) );
  INVX1 U392 ( .A(n51), .Y(n396) );
  INVX1 U393 ( .A(n396), .Y(n397) );
  BUFX2 U394 ( .A(n329), .Y(n398) );
  INVX1 U395 ( .A(n24), .Y(n399) );
  INVX1 U396 ( .A(n25), .Y(n400) );
  AND2X1 U397 ( .A(n413), .B(n136), .Y(n26) );
  INVX1 U398 ( .A(n26), .Y(n401) );
  AND2X1 U399 ( .A(n407), .B(n122), .Y(n23) );
  INVX1 U400 ( .A(n23), .Y(n402) );
  BUFX2 U401 ( .A(n124), .Y(n403) );
  AND2X1 U402 ( .A(n408), .B(n140), .Y(n27) );
  INVX1 U403 ( .A(n27), .Y(n404) );
  BUFX2 U404 ( .A(n130), .Y(n405) );
  INVX1 U405 ( .A(n131), .Y(n406) );
  INVX1 U406 ( .A(n123), .Y(n407) );
  AND2X1 U407 ( .A(A[1]), .B(n431), .Y(n141) );
  INVX1 U408 ( .A(n141), .Y(n408) );
  OR2X1 U409 ( .A(n432), .B(A[2]), .Y(n136) );
  INVX1 U410 ( .A(n136), .Y(n409) );
  AND2X1 U411 ( .A(n437), .B(A[7]), .Y(n111) );
  INVX1 U412 ( .A(n111), .Y(n410) );
  OR2X1 U413 ( .A(n431), .B(A[1]), .Y(n140) );
  INVX1 U414 ( .A(n140), .Y(n411) );
  AND2X2 U415 ( .A(A[4]), .B(n434), .Y(n128) );
  AND2X1 U416 ( .A(A[2]), .B(n432), .Y(n137) );
  INVX1 U417 ( .A(n21), .Y(n414) );
  INVX1 U418 ( .A(n39), .Y(n415) );
  INVX1 U419 ( .A(n122), .Y(n417) );
  INVX1 U420 ( .A(n139), .Y(n138) );
  INVX1 U421 ( .A(n318), .Y(n129) );
  XNOR2X1 U422 ( .A(n429), .B(n342), .Y(DIFF[26]) );
  INVX1 U423 ( .A(B[3]), .Y(n433) );
  INVX1 U424 ( .A(B[2]), .Y(n432) );
  INVX1 U425 ( .A(n308), .Y(n165) );
  INVX1 U426 ( .A(B[18]), .Y(n448) );
  INVX1 U427 ( .A(B[1]), .Y(n431) );
  OR2X1 U428 ( .A(A[23]), .B(n453), .Y(n419) );
  INVX1 U429 ( .A(B[19]), .Y(n449) );
  INVX1 U430 ( .A(B[10]), .Y(n440) );
  INVX1 U431 ( .A(B[4]), .Y(n434) );
  INVX1 U432 ( .A(B[8]), .Y(n438) );
  INVX1 U433 ( .A(B[9]), .Y(n439) );
  INVX1 U434 ( .A(B[24]), .Y(n454) );
  INVX1 U435 ( .A(B[17]), .Y(n447) );
  INVX1 U436 ( .A(B[16]), .Y(n446) );
  INVX1 U437 ( .A(B[14]), .Y(n444) );
  INVX1 U438 ( .A(B[6]), .Y(n436) );
  OR2X1 U439 ( .A(A[15]), .B(n445), .Y(n420) );
  OR2X1 U440 ( .A(A[21]), .B(n451), .Y(n421) );
  OR2X1 U441 ( .A(A[7]), .B(n437), .Y(n422) );
  OR2X1 U442 ( .A(A[11]), .B(n441), .Y(n423) );
  OR2X1 U443 ( .A(A[13]), .B(n443), .Y(n424) );
  OR2X1 U444 ( .A(A[9]), .B(n439), .Y(n425) );
  OR2X1 U445 ( .A(A[19]), .B(n449), .Y(n426) );
  INVX1 U446 ( .A(B[26]), .Y(n456) );
  INVX1 U447 ( .A(B[25]), .Y(n455) );
  INVX1 U448 ( .A(B[28]), .Y(n458) );
  INVX1 U449 ( .A(B[29]), .Y(n459) );
  INVX1 U450 ( .A(B[27]), .Y(n457) );
  XNOR2X1 U451 ( .A(A[31]), .B(B[31]), .Y(n1) );
  INVX1 U452 ( .A(B[0]), .Y(n430) );
  INVX1 U453 ( .A(B[30]), .Y(n460) );
  INVX1 U454 ( .A(B[12]), .Y(n442) );
  INVX1 U455 ( .A(B[13]), .Y(n443) );
  INVX1 U456 ( .A(B[11]), .Y(n441) );
  INVX1 U457 ( .A(B[7]), .Y(n437) );
  INVX1 U458 ( .A(B[23]), .Y(n453) );
  INVX1 U459 ( .A(B[22]), .Y(n452) );
  INVX1 U460 ( .A(B[20]), .Y(n450) );
  INVX1 U461 ( .A(B[21]), .Y(n451) );
  INVX1 U462 ( .A(B[15]), .Y(n445) );
  INVX1 U463 ( .A(B[5]), .Y(n435) );
  OR2X1 U464 ( .A(A[17]), .B(n447), .Y(n428) );
  INVX1 U465 ( .A(n320), .Y(n429) );
endmodule


module alu_DW_mult_uns_25 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n26, n27, n28, n29, n33, n34, n35,
         n36, n37, n41, n42, n43, n44, n45, n49, n50, n51, n52, n53, n57, n58,
         n59, n60, n61, n65, n66, n67, n68, n69, n73, n74, n75, n76, n77, n81,
         n82, n83, n84, n87, n88, n89, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n109, n110, n111, n115, n116,
         n117, n121, n122, n123, n124, n125, n129, n130, n131, n132, n133,
         n134, n136, n137, n138, n139, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n465, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796;
  assign product[0] = b[0];

  FAX1 U2 ( .A(a[15]), .B(n652), .C(n26), .YC(product[31]), .YS(product[30])
         );
  FAX1 U3 ( .A(n750), .B(n164), .C(n27), .YC(n26), .YS(product[29]) );
  FAX1 U4 ( .A(n165), .B(n166), .C(n28), .YC(n27), .YS(product[28]) );
  FAX1 U5 ( .A(n167), .B(n168), .C(n139), .YC(n28), .YS(product[27]) );
  XNOR2X1 U7 ( .A(n771), .B(n577), .Y(product[26]) );
  AOI21X1 U8 ( .A(n34), .B(n767), .C(n33), .Y(n29) );
  XOR2X1 U15 ( .A(n604), .B(n585), .Y(product[25]) );
  OAI21X1 U16 ( .A(n729), .B(n605), .C(n710), .Y(n34) );
  XNOR2X1 U21 ( .A(n551), .B(n576), .Y(product[24]) );
  AOI21X1 U22 ( .A(n42), .B(n768), .C(n41), .Y(n37) );
  XOR2X1 U29 ( .A(n602), .B(n584), .Y(product[23]) );
  OAI21X1 U30 ( .A(n558), .B(n746), .C(n726), .Y(n42) );
  XNOR2X1 U35 ( .A(n552), .B(n575), .Y(product[22]) );
  AOI21X1 U36 ( .A(n50), .B(n762), .C(n49), .Y(n45) );
  XOR2X1 U43 ( .A(n600), .B(n583), .Y(product[21]) );
  OAI21X1 U44 ( .A(n745), .B(n601), .C(n725), .Y(n50) );
  XNOR2X1 U49 ( .A(n549), .B(n574), .Y(product[20]) );
  AOI21X1 U50 ( .A(n58), .B(n765), .C(n57), .Y(n53) );
  XOR2X1 U57 ( .A(n597), .B(n582), .Y(product[19]) );
  OAI21X1 U58 ( .A(n747), .B(n598), .C(n727), .Y(n58) );
  XNOR2X1 U63 ( .A(n66), .B(n573), .Y(product[18]) );
  AOI21X1 U64 ( .A(n66), .B(n764), .C(n65), .Y(n61) );
  XOR2X1 U71 ( .A(n595), .B(n581), .Y(product[17]) );
  OAI21X1 U72 ( .A(n748), .B(n560), .C(n728), .Y(n66) );
  XNOR2X1 U77 ( .A(n548), .B(n671), .Y(product[16]) );
  AOI21X1 U78 ( .A(n74), .B(n760), .C(n73), .Y(n69) );
  XOR2X1 U85 ( .A(n738), .B(n682), .Y(product[15]) );
  OAI21X1 U86 ( .A(n711), .B(n738), .C(n744), .Y(n74) );
  XNOR2X1 U91 ( .A(n550), .B(n572), .Y(product[14]) );
  AOI21X1 U92 ( .A(n82), .B(n763), .C(n81), .Y(n77) );
  XOR2X1 U99 ( .A(n567), .B(n580), .Y(product[13]) );
  OAI21X1 U100 ( .A(n556), .B(n590), .C(n564), .Y(n82) );
  AOI21X1 U102 ( .A(n93), .B(n87), .C(n88), .Y(n84) );
  XNOR2X1 U109 ( .A(n94), .B(n571), .Y(product[12]) );
  AOI21X1 U110 ( .A(n94), .B(n778), .C(n93), .Y(n89) );
  XNOR2X1 U117 ( .A(n100), .B(n570), .Y(product[11]) );
  AOI21X1 U119 ( .A(n104), .B(n555), .C(n97), .Y(n95) );
  OAI21X1 U121 ( .A(n554), .B(n740), .C(n693), .Y(n97) );
  XOR2X1 U126 ( .A(n103), .B(n579), .Y(product[10]) );
  OAI21X1 U127 ( .A(n758), .B(n103), .C(n554), .Y(n100) );
  XOR2X1 U132 ( .A(n566), .B(n578), .Y(product[9]) );
  OAI21X1 U134 ( .A(n559), .B(n557), .C(n562), .Y(n104) );
  AOI21X1 U136 ( .A(n109), .B(n115), .C(n110), .Y(n106) );
  XNOR2X1 U143 ( .A(n116), .B(n569), .Y(product[8]) );
  AOI21X1 U144 ( .A(n116), .B(n766), .C(n115), .Y(n111) );
  XNOR2X1 U151 ( .A(n122), .B(n705), .Y(product[7]) );
  AOI21X1 U153 ( .A(n122), .B(n759), .C(n121), .Y(n117) );
  XOR2X1 U160 ( .A(n568), .B(n607), .Y(product[6]) );
  OAI21X1 U161 ( .A(n553), .B(n607), .C(n588), .Y(n122) );
  XNOR2X1 U166 ( .A(n130), .B(n670), .Y(product[5]) );
  AOI21X1 U167 ( .A(n130), .B(n769), .C(n129), .Y(n125) );
  XOR2X1 U174 ( .A(n660), .B(n739), .Y(product[4]) );
  OAI21X1 U175 ( .A(n739), .B(n712), .C(n683), .Y(n130) );
  XNOR2X1 U180 ( .A(n134), .B(n136), .Y(product[3]) );
  FAX1 U190 ( .A(a[14]), .B(n594), .C(n587), .YC(n164), .YS(n165) );
  FAX1 U191 ( .A(n730), .B(n731), .C(n170), .YC(n166), .YS(n167) );
  FAX1 U192 ( .A(n713), .B(n174), .C(n171), .YC(n168), .YS(n169) );
  FAX1 U193 ( .A(a[13]), .B(n662), .C(n661), .YC(n170), .YS(n171) );
  FAX1 U194 ( .A(n180), .B(n175), .C(n178), .YC(n172), .YS(n173) );
  FAX1 U195 ( .A(n609), .B(n610), .C(n608), .YC(n174), .YS(n175) );
  FAX1 U196 ( .A(n181), .B(n184), .C(n179), .YC(n176), .YS(n177) );
  FAX1 U197 ( .A(n685), .B(n684), .C(n186), .YC(n178), .YS(n179) );
  FAX1 U198 ( .A(a[12]), .B(n593), .C(n586), .YC(n180), .YS(n181) );
  FAX1 U199 ( .A(n187), .B(n185), .C(n190), .YC(n182), .YS(n183) );
  FAX1 U200 ( .A(n749), .B(n194), .C(n192), .YC(n184), .YS(n185) );
  FAX1 U201 ( .A(n642), .B(n643), .C(n641), .YC(n186), .YS(n187) );
  FAX1 U202 ( .A(n200), .B(n191), .C(n198), .YC(n188), .YS(n189) );
  FAX1 U203 ( .A(n202), .B(n195), .C(n193), .YC(n190), .YS(n191) );
  FAX1 U204 ( .A(n616), .B(n614), .C(n615), .YC(n192), .YS(n193) );
  FAX1 U205 ( .A(a[11]), .B(n647), .C(n646), .YC(n194), .YS(n195) );
  FAX1 U206 ( .A(n208), .B(n199), .C(n206), .YC(n196), .YS(n197) );
  FAX1 U207 ( .A(n210), .B(n203), .C(n201), .YC(n198), .YS(n199) );
  FAX1 U208 ( .A(n664), .B(n663), .C(n212), .YC(n200), .YS(n201) );
  FAX1 U209 ( .A(n620), .B(n619), .C(n621), .YC(n202), .YS(n203) );
  FAX1 U210 ( .A(n209), .B(n216), .C(n207), .YC(n204), .YS(n205) );
  FAX1 U211 ( .A(n213), .B(n211), .C(n218), .YC(n206), .YS(n207) );
  FAX1 U212 ( .A(n714), .B(n222), .C(n220), .YC(n208), .YS(n209) );
  FAX1 U213 ( .A(n628), .B(n627), .C(n626), .YC(n210), .YS(n211) );
  FAX1 U214 ( .A(a[10]), .B(n625), .C(n624), .YC(n212), .YS(n213) );
  FAX1 U215 ( .A(n219), .B(n226), .C(n217), .YC(n214), .YS(n215) );
  FAX1 U216 ( .A(n223), .B(n230), .C(n228), .YC(n216), .YS(n217) );
  FAX1 U217 ( .A(n234), .B(n232), .C(n221), .YC(n218), .YS(n219) );
  FAX1 U218 ( .A(n673), .B(n674), .C(n672), .YC(n220), .YS(n221) );
  FAX1 U219 ( .A(n632), .B(n633), .C(n631), .YC(n222), .YS(n223) );
  FAX1 U220 ( .A(n229), .B(n238), .C(n227), .YC(n224), .YS(n225) );
  FAX1 U221 ( .A(n242), .B(n231), .C(n240), .YC(n226), .YS(n227) );
  FAX1 U222 ( .A(n244), .B(n235), .C(n233), .YC(n228), .YS(n229) );
  FAX1 U223 ( .A(n698), .B(n697), .C(n246), .YC(n230), .YS(n231) );
  FAX1 U224 ( .A(n638), .B(n637), .C(n636), .YC(n232), .YS(n233) );
  FAX1 U225 ( .A(a[9]), .B(n696), .C(n695), .YC(n234), .YS(n235) );
  FAX1 U226 ( .A(n241), .B(n250), .C(n239), .YC(n236), .YS(n237) );
  FAX1 U227 ( .A(n254), .B(n243), .C(n252), .YC(n238), .YS(n239) );
  FAX1 U228 ( .A(n256), .B(n247), .C(n245), .YC(n240), .YS(n241) );
  FAX1 U229 ( .A(n751), .B(n260), .C(n258), .YC(n242), .YS(n243) );
  FAX1 U230 ( .A(n734), .B(n733), .C(n732), .YC(n244), .YS(n245) );
  FAX1 U231 ( .A(n654), .B(n655), .C(n653), .YC(n246), .YS(n247) );
  FAX1 U232 ( .A(n253), .B(n264), .C(n251), .YC(n248), .YS(n249) );
  FAX1 U233 ( .A(n268), .B(n255), .C(n266), .YC(n250), .YS(n251) );
  FAX1 U234 ( .A(n270), .B(n259), .C(n257), .YC(n252), .YS(n253) );
  FAX1 U235 ( .A(n701), .B(n272), .C(n261), .YC(n254), .YS(n255) );
  FAX1 U236 ( .A(n650), .B(n648), .C(n649), .YC(n256), .YS(n257) );
  FAX1 U237 ( .A(n721), .B(n719), .C(n720), .YC(n258), .YS(n259) );
  HAX1 U238 ( .A(a[8]), .B(n680), .YC(n260), .YS(n261) );
  FAX1 U239 ( .A(n267), .B(n276), .C(n265), .YC(n262), .YS(n263) );
  FAX1 U240 ( .A(n271), .B(n269), .C(n278), .YC(n264), .YS(n265) );
  FAX1 U241 ( .A(n273), .B(n282), .C(n280), .YC(n266), .YS(n267) );
  FAX1 U242 ( .A(n657), .B(n656), .C(n284), .YC(n268), .YS(n269) );
  FAX1 U243 ( .A(n666), .B(n667), .C(n665), .YC(n270), .YS(n271) );
  HAX1 U244 ( .A(n629), .B(n630), .YC(n272), .YS(n273) );
  FAX1 U245 ( .A(n279), .B(n288), .C(n277), .YC(n274), .YS(n275) );
  FAX1 U246 ( .A(n283), .B(n281), .C(n290), .YC(n276), .YS(n277) );
  FAX1 U247 ( .A(n294), .B(n285), .C(n292), .YC(n278), .YS(n279) );
  FAX1 U248 ( .A(n704), .B(n703), .C(n702), .YC(n280), .YS(n281) );
  FAX1 U249 ( .A(n754), .B(n753), .C(n752), .YC(n282), .YS(n283) );
  HAX1 U250 ( .A(n547), .B(n565), .YC(n284), .YS(n285) );
  FAX1 U251 ( .A(n291), .B(n298), .C(n289), .YC(n286), .YS(n287) );
  FAX1 U252 ( .A(n302), .B(n293), .C(n300), .YC(n288), .YS(n289) );
  FAX1 U253 ( .A(n700), .B(n304), .C(n295), .YC(n290), .YS(n291) );
  FAX1 U254 ( .A(n717), .B(n718), .C(n716), .YC(n292), .YS(n293) );
  HAX1 U255 ( .A(n617), .B(n618), .YC(n294), .YS(n295) );
  FAX1 U256 ( .A(n301), .B(n308), .C(n299), .YC(n296), .YS(n297) );
  FAX1 U257 ( .A(n305), .B(n310), .C(n303), .YC(n298), .YS(n299) );
  FAX1 U258 ( .A(n659), .B(n658), .C(n312), .YC(n300), .YS(n301) );
  FAX1 U259 ( .A(n688), .B(n686), .C(n687), .YC(n302), .YS(n303) );
  HAX1 U260 ( .A(a[6]), .B(n611), .YC(n304), .YS(n305) );
  FAX1 U261 ( .A(n311), .B(n316), .C(n309), .YC(n306), .YS(n307) );
  FAX1 U262 ( .A(n320), .B(n313), .C(n318), .YC(n308), .YS(n309) );
  FAX1 U263 ( .A(n679), .B(n677), .C(n678), .YC(n310), .YS(n311) );
  HAX1 U264 ( .A(n612), .B(n613), .YC(n312), .YS(n313) );
  FAX1 U265 ( .A(n319), .B(n324), .C(n317), .YC(n314), .YS(n315) );
  FAX1 U266 ( .A(n715), .B(n326), .C(n321), .YC(n316), .YS(n317) );
  FAX1 U267 ( .A(n676), .B(n442), .C(n675), .YC(n318), .YS(n319) );
  HAX1 U268 ( .A(a[5]), .B(n722), .YC(n320), .YS(n321) );
  FAX1 U270 ( .A(n669), .B(n668), .C(n332), .YC(n324), .YS(n325) );
  HAX1 U271 ( .A(n634), .B(n635), .YC(n326), .YS(n327) );
  FAX1 U272 ( .A(n336), .B(n333), .C(n331), .YC(n328), .YS(n329) );
  FAX1 U273 ( .A(n737), .B(n736), .C(n735), .YC(n330), .YS(n331) );
  HAX1 U274 ( .A(a[4]), .B(n644), .YC(n332), .YS(n333) );
  FAX1 U275 ( .A(n699), .B(n340), .C(n337), .YC(n334), .YS(n335) );
  HAX1 U276 ( .A(n622), .B(n623), .YC(n336), .YS(n337) );
  FAX1 U277 ( .A(n756), .B(n755), .C(n342), .YC(n338), .YS(n339) );
  HAX1 U278 ( .A(a[3]), .B(n681), .YC(n340), .YS(n341) );
  HAX1 U279 ( .A(n639), .B(n640), .YC(n342), .YS(n343) );
  HAX1 U280 ( .A(a[2]), .B(n462), .YC(n344), .YS(n345) );
  INVX8 U434 ( .A(b[8]), .Y(n788) );
  INVX1 U435 ( .A(n787), .Y(n547) );
  INVX8 U436 ( .A(b[7]), .Y(n787) );
  OR2X1 U437 ( .A(n796), .B(n792), .Y(n348) );
  OR2X1 U438 ( .A(n781), .B(n783), .Y(n461) );
  OR2X1 U439 ( .A(n796), .B(n793), .Y(n347) );
  OR2X1 U440 ( .A(n780), .B(n779), .Y(n465) );
  OR2X1 U441 ( .A(n793), .B(n784), .Y(n382) );
  OR2X1 U442 ( .A(n796), .B(n783), .Y(n357) );
  OR2X1 U443 ( .A(n793), .B(n782), .Y(n385) );
  OR2X1 U444 ( .A(n796), .B(n779), .Y(n360) );
  OR2X1 U445 ( .A(n786), .B(n793), .Y(n381) );
  OR2X1 U446 ( .A(n795), .B(n782), .Y(n372) );
  OR2X1 U447 ( .A(n790), .B(n784), .Y(n415) );
  OR2X1 U448 ( .A(n789), .B(n784), .Y(n424) );
  OR2X1 U449 ( .A(n791), .B(n782), .Y(n408) );
  OR2X1 U450 ( .A(n787), .B(n783), .Y(n441) );
  OR2X1 U451 ( .A(n791), .B(n793), .Y(n376) );
  OR2X1 U452 ( .A(n795), .B(n790), .Y(n364) );
  OR2X1 U453 ( .A(n795), .B(n789), .Y(n365) );
  OR2X1 U454 ( .A(n795), .B(n784), .Y(n369) );
  OR2X1 U455 ( .A(n784), .B(n792), .Y(n394) );
  OR2X1 U456 ( .A(n791), .B(n784), .Y(n405) );
  OR2X1 U457 ( .A(n792), .B(n782), .Y(n397) );
  OR2X1 U458 ( .A(n791), .B(n783), .Y(n407) );
  INVX1 U459 ( .A(n433), .Y(n717) );
  INVX1 U460 ( .A(n410), .Y(n688) );
  INVX1 U461 ( .A(n419), .Y(n687) );
  OR2X1 U462 ( .A(n784), .B(n776), .Y(n451) );
  OR2X1 U463 ( .A(n784), .B(n783), .Y(n452) );
  OR2X1 U464 ( .A(n788), .B(n779), .Y(n437) );
  OR2X1 U465 ( .A(n780), .B(n784), .Y(n454) );
  OR2X1 U466 ( .A(n796), .B(n791), .Y(n349) );
  OR2X1 U467 ( .A(n740), .B(n758), .Y(n96) );
  AND2X1 U468 ( .A(b[7]), .B(b[2]), .Y(n442) );
  INVX1 U469 ( .A(n429), .Y(n676) );
  AND2X1 U470 ( .A(n327), .B(n325), .Y(n774) );
  AND2X1 U471 ( .A(n766), .B(n109), .Y(n105) );
  AND2X1 U472 ( .A(n761), .B(n87), .Y(n83) );
  OR2X1 U473 ( .A(n287), .B(n296), .Y(n87) );
  AND2X1 U474 ( .A(n314), .B(n307), .Y(n99) );
  AND2X1 U475 ( .A(n341), .B(n339), .Y(n124) );
  OR2X1 U476 ( .A(n776), .B(n779), .Y(n459) );
  AND2X1 U477 ( .A(b[3]), .B(b[0]), .Y(n462) );
  AND2X1 U478 ( .A(n651), .B(n138), .Y(n133) );
  OR2X1 U479 ( .A(n796), .B(n795), .Y(n346) );
  AND2X1 U480 ( .A(n554), .B(n101), .Y(n17) );
  AND2X1 U481 ( .A(n137), .B(n757), .Y(product[2]) );
  OR2X1 U482 ( .A(n784), .B(n782), .Y(n453) );
  INVX8 U483 ( .A(b[2]), .Y(n782) );
  OR2X1 U484 ( .A(n788), .B(n782), .Y(n435) );
  OR2X1 U485 ( .A(n785), .B(n782), .Y(n448) );
  OR2X1 U486 ( .A(n789), .B(n782), .Y(n427) );
  OR2X1 U487 ( .A(n776), .B(n782), .Y(n457) );
  OR2X1 U488 ( .A(n783), .B(n782), .Y(n460) );
  OR2X1 U489 ( .A(n790), .B(n782), .Y(n418) );
  INVX2 U490 ( .A(b[4]), .Y(n776) );
  INVX2 U491 ( .A(b[11]), .Y(n791) );
  INVX8 U492 ( .A(b[10]), .Y(n790) );
  INVX1 U493 ( .A(b[14]), .Y(n795) );
  INVX2 U494 ( .A(b[9]), .Y(n789) );
  INVX2 U495 ( .A(b[3]), .Y(n783) );
  OR2X1 U496 ( .A(n307), .B(n314), .Y(n98) );
  AND2X1 U497 ( .A(n296), .B(n287), .Y(n88) );
  OR2X1 U498 ( .A(n263), .B(n274), .Y(n75) );
  AND2X1 U499 ( .A(a[1]), .B(n645), .Y(n138) );
  INVX1 U500 ( .A(n101), .Y(n758) );
  OR2X1 U501 ( .A(n315), .B(n591), .Y(n101) );
  OR2X1 U502 ( .A(n345), .B(n694), .Y(n131) );
  OR2X1 U503 ( .A(n796), .B(n790), .Y(n350) );
  OR2X1 U504 ( .A(n796), .B(n784), .Y(n355) );
  OR2X1 U505 ( .A(n796), .B(n782), .Y(n358) );
  INVX1 U506 ( .A(b[1]), .Y(n780) );
  OAI21X1 U507 ( .A(n711), .B(n738), .C(n744), .Y(n548) );
  BUFX2 U508 ( .A(n58), .Y(n549) );
  BUFX2 U509 ( .A(n82), .Y(n550) );
  OAI21X1 U510 ( .A(n558), .B(n746), .C(n726), .Y(n551) );
  BUFX2 U511 ( .A(n50), .Y(n552) );
  OR2X1 U512 ( .A(n339), .B(n341), .Y(n123) );
  INVX8 U513 ( .A(b[0]), .Y(n779) );
  OR2X2 U514 ( .A(n787), .B(n784), .Y(n439) );
  OR2X2 U515 ( .A(n785), .B(n784), .Y(n445) );
  INVX1 U516 ( .A(n123), .Y(n553) );
  OR2X2 U517 ( .A(n773), .B(n592), .Y(n591) );
  OR2X2 U518 ( .A(n775), .B(n774), .Y(n592) );
  AND2X2 U519 ( .A(n591), .B(n315), .Y(n102) );
  INVX1 U520 ( .A(n102), .Y(n554) );
  INVX1 U521 ( .A(n96), .Y(n555) );
  INVX1 U522 ( .A(n83), .Y(n556) );
  INVX1 U523 ( .A(n105), .Y(n557) );
  BUFX2 U524 ( .A(n45), .Y(n558) );
  BUFX2 U525 ( .A(n117), .Y(n559) );
  BUFX2 U526 ( .A(n69), .Y(n560) );
  AND2X1 U527 ( .A(n330), .B(n325), .Y(n773) );
  AND2X1 U528 ( .A(n327), .B(n330), .Y(n775) );
  OR2X1 U529 ( .A(n645), .B(a[1]), .Y(n137) );
  INVX1 U530 ( .A(n106), .Y(n561) );
  INVX1 U531 ( .A(n561), .Y(n562) );
  INVX1 U532 ( .A(n84), .Y(n563) );
  INVX1 U533 ( .A(n563), .Y(n564) );
  OR2X1 U534 ( .A(n784), .B(n788), .Y(n432) );
  INVX1 U535 ( .A(n432), .Y(n565) );
  BUFX2 U536 ( .A(n111), .Y(n566) );
  BUFX2 U537 ( .A(n89), .Y(n567) );
  AND2X1 U538 ( .A(n588), .B(n123), .Y(n21) );
  INVX1 U539 ( .A(n21), .Y(n568) );
  AND2X1 U540 ( .A(n742), .B(n766), .Y(n19) );
  INVX1 U541 ( .A(n19), .Y(n569) );
  AND2X1 U542 ( .A(n693), .B(n98), .Y(n16) );
  INVX1 U543 ( .A(n16), .Y(n570) );
  AND2X1 U544 ( .A(n743), .B(n778), .Y(n15) );
  INVX1 U545 ( .A(n15), .Y(n571) );
  AND2X1 U546 ( .A(n692), .B(n763), .Y(n13) );
  INVX1 U547 ( .A(n13), .Y(n572) );
  AND2X1 U548 ( .A(n709), .B(n764), .Y(n9) );
  INVX1 U549 ( .A(n9), .Y(n573) );
  AND2X1 U550 ( .A(n708), .B(n765), .Y(n7) );
  INVX1 U551 ( .A(n7), .Y(n574) );
  AND2X1 U552 ( .A(n690), .B(n762), .Y(n5) );
  INVX1 U553 ( .A(n5), .Y(n575) );
  AND2X1 U554 ( .A(n689), .B(n768), .Y(n3) );
  INVX1 U555 ( .A(n3), .Y(n576) );
  AND2X1 U556 ( .A(n741), .B(n767), .Y(n1) );
  INVX1 U557 ( .A(n1), .Y(n577) );
  AND2X1 U558 ( .A(n707), .B(n109), .Y(n18) );
  INVX1 U559 ( .A(n18), .Y(n578) );
  INVX1 U560 ( .A(n17), .Y(n579) );
  AND2X1 U561 ( .A(n706), .B(n87), .Y(n14) );
  INVX1 U562 ( .A(n14), .Y(n580) );
  AND2X1 U563 ( .A(n728), .B(n67), .Y(n10) );
  INVX1 U564 ( .A(n10), .Y(n581) );
  AND2X1 U565 ( .A(n727), .B(n59), .Y(n8) );
  INVX1 U566 ( .A(n8), .Y(n582) );
  AND2X1 U567 ( .A(n725), .B(n51), .Y(n6) );
  INVX1 U568 ( .A(n6), .Y(n583) );
  AND2X1 U569 ( .A(n726), .B(n43), .Y(n4) );
  INVX1 U570 ( .A(n4), .Y(n584) );
  AND2X1 U571 ( .A(n710), .B(n35), .Y(n2) );
  INVX1 U572 ( .A(n2), .Y(n585) );
  OR2X1 U573 ( .A(n793), .B(n790), .Y(n377) );
  INVX1 U574 ( .A(n377), .Y(n586) );
  INVX1 U575 ( .A(n348), .Y(n587) );
  INVX1 U576 ( .A(n124), .Y(n588) );
  INVX1 U577 ( .A(n95), .Y(n589) );
  INVX1 U578 ( .A(n589), .Y(n590) );
  OR2X1 U579 ( .A(n791), .B(n792), .Y(n388) );
  INVX1 U580 ( .A(n388), .Y(n593) );
  OR2X1 U581 ( .A(n795), .B(n793), .Y(n361) );
  INVX1 U582 ( .A(n361), .Y(n594) );
  BUFX2 U583 ( .A(n560), .Y(n595) );
  INVX1 U584 ( .A(n61), .Y(n596) );
  INVX1 U585 ( .A(n596), .Y(n597) );
  INVX1 U586 ( .A(n596), .Y(n598) );
  INVX1 U587 ( .A(n53), .Y(n599) );
  INVX1 U588 ( .A(n599), .Y(n600) );
  INVX1 U589 ( .A(n599), .Y(n601) );
  BUFX2 U590 ( .A(n558), .Y(n602) );
  INVX1 U591 ( .A(n37), .Y(n603) );
  INVX1 U592 ( .A(n603), .Y(n604) );
  INVX1 U593 ( .A(n603), .Y(n605) );
  INVX1 U594 ( .A(n125), .Y(n606) );
  INVX1 U595 ( .A(n606), .Y(n607) );
  OR2X1 U596 ( .A(n796), .B(n789), .Y(n351) );
  INVX1 U597 ( .A(n351), .Y(n608) );
  INVX1 U598 ( .A(n364), .Y(n609) );
  INVX1 U599 ( .A(n376), .Y(n610) );
  OR2X1 U600 ( .A(n783), .B(n788), .Y(n434) );
  INVX1 U601 ( .A(n434), .Y(n611) );
  INVX1 U602 ( .A(n435), .Y(n612) );
  OR2X1 U603 ( .A(n780), .B(n789), .Y(n428) );
  INVX1 U604 ( .A(n428), .Y(n613) );
  OR2X1 U605 ( .A(n795), .B(n787), .Y(n367) );
  INVX1 U606 ( .A(n367), .Y(n614) );
  OR2X1 U607 ( .A(n796), .B(n786), .Y(n354) );
  INVX1 U608 ( .A(n354), .Y(n615) );
  OR2X1 U609 ( .A(n791), .B(n790), .Y(n400) );
  INVX1 U610 ( .A(n400), .Y(n616) );
  OR2X1 U611 ( .A(n792), .B(n779), .Y(n399) );
  INVX1 U612 ( .A(n399), .Y(n617) );
  OR2X1 U613 ( .A(n780), .B(n791), .Y(n409) );
  INVX1 U614 ( .A(n409), .Y(n618) );
  OR2X1 U615 ( .A(n795), .B(n786), .Y(n368) );
  INVX1 U616 ( .A(n368), .Y(n619) );
  OR2X1 U617 ( .A(n792), .B(n788), .Y(n391) );
  INVX1 U618 ( .A(n391), .Y(n620) );
  INVX1 U619 ( .A(n355), .Y(n621) );
  INVX1 U620 ( .A(n457), .Y(n622) );
  INVX1 U621 ( .A(n454), .Y(n623) );
  OR2X1 U622 ( .A(n787), .B(n792), .Y(n392) );
  INVX1 U623 ( .A(n392), .Y(n624) );
  OR2X1 U624 ( .A(n791), .B(n788), .Y(n402) );
  INVX1 U625 ( .A(n402), .Y(n625) );
  OR2X1 U626 ( .A(n796), .B(n776), .Y(n356) );
  INVX1 U627 ( .A(n356), .Y(n626) );
  INVX1 U628 ( .A(n381), .Y(n627) );
  OR2X1 U629 ( .A(n789), .B(n790), .Y(n411) );
  INVX1 U630 ( .A(n411), .Y(n628) );
  INVX1 U631 ( .A(n397), .Y(n629) );
  OR2X1 U632 ( .A(n780), .B(n793), .Y(n386) );
  INVX1 U633 ( .A(n386), .Y(n630) );
  INVX1 U634 ( .A(n357), .Y(n631) );
  OR2X1 U635 ( .A(n790), .B(n788), .Y(n412) );
  INVX1 U636 ( .A(n412), .Y(n632) );
  OR2X1 U637 ( .A(n787), .B(n791), .Y(n403) );
  INVX1 U638 ( .A(n403), .Y(n633) );
  INVX1 U639 ( .A(n437), .Y(n634) );
  OR2X1 U640 ( .A(n780), .B(n787), .Y(n443) );
  INVX1 U641 ( .A(n443), .Y(n635) );
  INVX1 U642 ( .A(n358), .Y(n636) );
  OR2X1 U643 ( .A(n786), .B(n791), .Y(n404) );
  INVX1 U644 ( .A(n404), .Y(n637) );
  OR2X1 U645 ( .A(n789), .B(n788), .Y(n421) );
  INVX1 U646 ( .A(n421), .Y(n638) );
  INVX1 U647 ( .A(n459), .Y(n639) );
  INVX1 U648 ( .A(n461), .Y(n640) );
  OR2X1 U649 ( .A(n796), .B(n787), .Y(n353) );
  INVX1 U650 ( .A(n353), .Y(n641) );
  OR2X1 U651 ( .A(n790), .B(n792), .Y(n389) );
  INVX1 U652 ( .A(n389), .Y(n642) );
  OR2X1 U653 ( .A(n789), .B(n793), .Y(n378) );
  INVX1 U654 ( .A(n378), .Y(n643) );
  INVX1 U655 ( .A(n453), .Y(n644) );
  INVX1 U656 ( .A(n465), .Y(n645) );
  OR2X1 U657 ( .A(n789), .B(n792), .Y(n390) );
  INVX1 U658 ( .A(n390), .Y(n646) );
  OR2X1 U659 ( .A(n793), .B(n788), .Y(n379) );
  INVX1 U660 ( .A(n379), .Y(n647) );
  INVX1 U661 ( .A(n415), .Y(n648) );
  OR2X1 U662 ( .A(n786), .B(n789), .Y(n423) );
  INVX1 U663 ( .A(n423), .Y(n649) );
  OR2X1 U664 ( .A(n791), .B(n776), .Y(n406) );
  INVX1 U665 ( .A(n406), .Y(n650) );
  OR2X1 U666 ( .A(n782), .B(n779), .Y(n134) );
  INVX1 U667 ( .A(n134), .Y(n651) );
  INVX1 U668 ( .A(n346), .Y(n652) );
  OR2X1 U669 ( .A(n796), .B(n780), .Y(n359) );
  INVX1 U670 ( .A(n359), .Y(n653) );
  OR2X1 U671 ( .A(n792), .B(n776), .Y(n395) );
  INVX1 U672 ( .A(n395), .Y(n654) );
  OR2X1 U673 ( .A(n787), .B(n789), .Y(n422) );
  INVX1 U674 ( .A(n422), .Y(n655) );
  OR2X1 U675 ( .A(n786), .B(n788), .Y(n431) );
  INVX1 U676 ( .A(n431), .Y(n656) );
  INVX1 U677 ( .A(n407), .Y(n657) );
  OR2X1 U678 ( .A(n787), .B(n776), .Y(n440) );
  INVX1 U679 ( .A(n440), .Y(n658) );
  INVX1 U680 ( .A(n427), .Y(n659) );
  AND2X1 U681 ( .A(n683), .B(n131), .Y(n23) );
  INVX1 U682 ( .A(n23), .Y(n660) );
  OR2X1 U683 ( .A(n795), .B(n791), .Y(n363) );
  INVX1 U684 ( .A(n363), .Y(n661) );
  OR2X1 U685 ( .A(n794), .B(n792), .Y(n375) );
  INVX1 U686 ( .A(n375), .Y(n662) );
  OR2X1 U687 ( .A(n789), .B(n791), .Y(n401) );
  INVX1 U688 ( .A(n401), .Y(n663) );
  OR2X1 U689 ( .A(n787), .B(n793), .Y(n380) );
  INVX1 U690 ( .A(n380), .Y(n664) );
  OR2X1 U691 ( .A(n795), .B(n779), .Y(n374) );
  INVX1 U692 ( .A(n374), .Y(n665) );
  OR2X1 U693 ( .A(n790), .B(n776), .Y(n416) );
  INVX1 U694 ( .A(n416), .Y(n666) );
  INVX1 U695 ( .A(n424), .Y(n667) );
  INVX1 U696 ( .A(n448), .Y(n668) );
  INVX1 U697 ( .A(n452), .Y(n669) );
  AND2X1 U698 ( .A(n724), .B(n769), .Y(n22) );
  INVX1 U699 ( .A(n22), .Y(n670) );
  AND2X1 U700 ( .A(n691), .B(n760), .Y(n11) );
  INVX1 U701 ( .A(n11), .Y(n671) );
  OR2X1 U702 ( .A(n795), .B(n776), .Y(n370) );
  INVX1 U703 ( .A(n370), .Y(n672) );
  OR2X1 U704 ( .A(n786), .B(n792), .Y(n393) );
  INVX1 U705 ( .A(n393), .Y(n673) );
  INVX1 U706 ( .A(n382), .Y(n674) );
  OR2X1 U707 ( .A(n780), .B(n788), .Y(n436) );
  INVX1 U708 ( .A(n436), .Y(n675) );
  OR2X1 U709 ( .A(n789), .B(n779), .Y(n429) );
  OR2X1 U710 ( .A(n785), .B(n776), .Y(n446) );
  INVX1 U711 ( .A(n446), .Y(n677) );
  INVX1 U712 ( .A(n441), .Y(n678) );
  OR2X1 U713 ( .A(n790), .B(n779), .Y(n420) );
  INVX1 U714 ( .A(n420), .Y(n679) );
  OR2X1 U715 ( .A(n792), .B(n783), .Y(n396) );
  INVX1 U716 ( .A(n396), .Y(n680) );
  INVX1 U717 ( .A(n460), .Y(n681) );
  AND2X1 U718 ( .A(n744), .B(n75), .Y(n12) );
  INVX1 U719 ( .A(n12), .Y(n682) );
  AND2X1 U720 ( .A(n694), .B(n345), .Y(n132) );
  INVX1 U721 ( .A(n132), .Y(n683) );
  OR2X1 U722 ( .A(n796), .B(n788), .Y(n352) );
  INVX1 U723 ( .A(n352), .Y(n684) );
  INVX1 U724 ( .A(n365), .Y(n685) );
  INVX1 U725 ( .A(n445), .Y(n686) );
  OR2X1 U726 ( .A(n780), .B(n790), .Y(n419) );
  OR2X1 U727 ( .A(n791), .B(n779), .Y(n410) );
  OR2X1 U728 ( .A(n323), .B(n328), .Y(n109) );
  AND2X1 U729 ( .A(n182), .B(n177), .Y(n41) );
  INVX1 U730 ( .A(n41), .Y(n689) );
  AND2X1 U731 ( .A(n189), .B(n196), .Y(n49) );
  INVX1 U732 ( .A(n49), .Y(n690) );
  AND2X1 U733 ( .A(n262), .B(n249), .Y(n73) );
  INVX1 U734 ( .A(n73), .Y(n691) );
  AND2X1 U735 ( .A(n286), .B(n275), .Y(n81) );
  INVX1 U736 ( .A(n81), .Y(n692) );
  INVX1 U737 ( .A(n99), .Y(n693) );
  OR2X1 U738 ( .A(n780), .B(n782), .Y(n463) );
  INVX1 U739 ( .A(n463), .Y(n694) );
  INVX1 U740 ( .A(n394), .Y(n695) );
  OR2X1 U741 ( .A(n793), .B(n776), .Y(n383) );
  INVX1 U742 ( .A(n383), .Y(n696) );
  OR2X1 U743 ( .A(n795), .B(n783), .Y(n371) );
  INVX1 U744 ( .A(n371), .Y(n697) );
  OR2X1 U745 ( .A(n787), .B(n790), .Y(n413) );
  INVX1 U746 ( .A(n413), .Y(n698) );
  OR2X1 U747 ( .A(n786), .B(n779), .Y(n450) );
  INVX1 U748 ( .A(n450), .Y(n699) );
  INVX1 U749 ( .A(n418), .Y(n700) );
  OR2X1 U750 ( .A(n787), .B(n788), .Y(n430) );
  INVX1 U751 ( .A(n430), .Y(n701) );
  OR2X1 U752 ( .A(n789), .B(n776), .Y(n425) );
  INVX1 U753 ( .A(n425), .Y(n702) );
  INVX1 U754 ( .A(n408), .Y(n703) );
  OR2X1 U755 ( .A(n794), .B(n779), .Y(n387) );
  INVX1 U756 ( .A(n387), .Y(n704) );
  AND2X1 U757 ( .A(n723), .B(n759), .Y(n20) );
  INVX1 U758 ( .A(n20), .Y(n705) );
  INVX1 U759 ( .A(n88), .Y(n706) );
  AND2X1 U760 ( .A(n328), .B(n323), .Y(n110) );
  INVX1 U761 ( .A(n110), .Y(n707) );
  AND2X1 U762 ( .A(n214), .B(n205), .Y(n57) );
  INVX1 U763 ( .A(n57), .Y(n708) );
  AND2X1 U764 ( .A(n236), .B(n225), .Y(n65) );
  INVX1 U765 ( .A(n65), .Y(n709) );
  AND2X1 U766 ( .A(n173), .B(n176), .Y(n36) );
  INVX1 U767 ( .A(n36), .Y(n710) );
  INVX1 U768 ( .A(n75), .Y(n711) );
  INVX1 U769 ( .A(n131), .Y(n712) );
  INVX1 U770 ( .A(n350), .Y(n713) );
  INVX1 U771 ( .A(n369), .Y(n714) );
  OR2X1 U772 ( .A(n785), .B(n783), .Y(n447) );
  INVX1 U773 ( .A(n447), .Y(n715) );
  INVX1 U774 ( .A(n439), .Y(n716) );
  OR2X1 U775 ( .A(n776), .B(n788), .Y(n433) );
  OR2X1 U776 ( .A(n789), .B(n783), .Y(n426) );
  INVX1 U777 ( .A(n426), .Y(n718) );
  OR2X1 U778 ( .A(n780), .B(n795), .Y(n373) );
  INVX1 U779 ( .A(n373), .Y(n719) );
  INVX1 U780 ( .A(n360), .Y(n720) );
  INVX1 U781 ( .A(n385), .Y(n721) );
  INVX1 U782 ( .A(n451), .Y(n722) );
  AND2X1 U783 ( .A(n338), .B(n335), .Y(n121) );
  INVX1 U784 ( .A(n121), .Y(n723) );
  AND2X1 U785 ( .A(n344), .B(n343), .Y(n129) );
  INVX1 U786 ( .A(n129), .Y(n724) );
  AND2X1 U787 ( .A(n197), .B(n204), .Y(n52) );
  INVX1 U788 ( .A(n52), .Y(n725) );
  AND2X1 U789 ( .A(n183), .B(n188), .Y(n44) );
  INVX1 U790 ( .A(n44), .Y(n726) );
  AND2X1 U791 ( .A(n224), .B(n215), .Y(n60) );
  INVX1 U792 ( .A(n60), .Y(n727) );
  AND2X1 U793 ( .A(n248), .B(n237), .Y(n68) );
  INVX1 U794 ( .A(n68), .Y(n728) );
  OR2X1 U795 ( .A(n176), .B(n173), .Y(n35) );
  INVX1 U796 ( .A(n35), .Y(n729) );
  OR2X1 U797 ( .A(n795), .B(n792), .Y(n362) );
  INVX1 U798 ( .A(n362), .Y(n730) );
  INVX1 U799 ( .A(n349), .Y(n731) );
  INVX1 U800 ( .A(n372), .Y(n732) );
  OR2X1 U801 ( .A(n786), .B(n790), .Y(n414) );
  INVX1 U802 ( .A(n414), .Y(n733) );
  OR2X1 U803 ( .A(n793), .B(n783), .Y(n384) );
  INVX1 U804 ( .A(n384), .Y(n734) );
  OR2X1 U805 ( .A(n780), .B(n785), .Y(n449) );
  INVX1 U806 ( .A(n449), .Y(n735) );
  OR2X1 U807 ( .A(n787), .B(n779), .Y(n444) );
  INVX1 U808 ( .A(n444), .Y(n736) );
  OR2X1 U809 ( .A(n783), .B(n776), .Y(n456) );
  INVX1 U810 ( .A(n456), .Y(n737) );
  BUFX2 U811 ( .A(n77), .Y(n738) );
  INVX1 U812 ( .A(n133), .Y(n739) );
  INVX1 U813 ( .A(n98), .Y(n740) );
  AND2X1 U814 ( .A(n169), .B(n172), .Y(n33) );
  INVX1 U815 ( .A(n33), .Y(n741) );
  AND2X1 U816 ( .A(n334), .B(n329), .Y(n115) );
  INVX1 U817 ( .A(n115), .Y(n742) );
  AND2X1 U818 ( .A(n306), .B(n297), .Y(n93) );
  INVX1 U819 ( .A(n93), .Y(n743) );
  AND2X1 U820 ( .A(n274), .B(n263), .Y(n76) );
  INVX1 U821 ( .A(n76), .Y(n744) );
  OR2X1 U822 ( .A(n204), .B(n197), .Y(n51) );
  INVX1 U823 ( .A(n51), .Y(n745) );
  OR2X1 U824 ( .A(n188), .B(n183), .Y(n43) );
  INVX1 U825 ( .A(n43), .Y(n746) );
  OR2X1 U826 ( .A(n215), .B(n224), .Y(n59) );
  INVX1 U827 ( .A(n59), .Y(n747) );
  OR2X1 U828 ( .A(n237), .B(n248), .Y(n67) );
  INVX1 U829 ( .A(n67), .Y(n748) );
  OR2X1 U830 ( .A(n795), .B(n788), .Y(n366) );
  INVX1 U831 ( .A(n366), .Y(n749) );
  INVX1 U832 ( .A(n347), .Y(n750) );
  INVX1 U833 ( .A(n405), .Y(n751) );
  OR2X1 U834 ( .A(n787), .B(n786), .Y(n438) );
  INVX1 U835 ( .A(n438), .Y(n752) );
  OR2X1 U836 ( .A(n780), .B(n792), .Y(n398) );
  INVX1 U837 ( .A(n398), .Y(n753) );
  OR2X1 U838 ( .A(n790), .B(n783), .Y(n417) );
  INVX1 U839 ( .A(n417), .Y(n754) );
  OR2X1 U840 ( .A(n781), .B(n776), .Y(n458) );
  INVX1 U841 ( .A(n458), .Y(n755) );
  OR2X1 U842 ( .A(n784), .B(n779), .Y(n455) );
  INVX1 U843 ( .A(n455), .Y(n756) );
  INVX1 U844 ( .A(n138), .Y(n757) );
  OR2X1 U845 ( .A(n335), .B(n338), .Y(n759) );
  OR2X1 U846 ( .A(n249), .B(n262), .Y(n760) );
  OR2X1 U847 ( .A(n306), .B(n297), .Y(n761) );
  OR2X1 U848 ( .A(n196), .B(n189), .Y(n762) );
  OR2X1 U849 ( .A(n275), .B(n286), .Y(n763) );
  OR2X1 U850 ( .A(n225), .B(n236), .Y(n764) );
  OR2X1 U851 ( .A(n205), .B(n214), .Y(n765) );
  INVX1 U852 ( .A(n29), .Y(n139) );
  OR2X1 U853 ( .A(n329), .B(n334), .Y(n766) );
  OR2X1 U854 ( .A(n172), .B(n169), .Y(n767) );
  OR2X1 U855 ( .A(n177), .B(n182), .Y(n768) );
  OR2X1 U856 ( .A(n343), .B(n344), .Y(n769) );
  INVX1 U857 ( .A(b[13]), .Y(n793) );
  INVX1 U858 ( .A(b[15]), .Y(n796) );
  INVX1 U859 ( .A(b[13]), .Y(n794) );
  INVX1 U860 ( .A(b[6]), .Y(n785) );
  INVX1 U861 ( .A(b[12]), .Y(n792) );
  INVX1 U862 ( .A(b[1]), .Y(n781) );
  BUFX2 U863 ( .A(n34), .Y(n771) );
  XOR2X1 U864 ( .A(n330), .B(n327), .Y(n772) );
  XOR2X1 U865 ( .A(n325), .B(n772), .Y(n323) );
  INVX1 U866 ( .A(n761), .Y(n777) );
  INVX1 U867 ( .A(n777), .Y(n778) );
  INVX1 U868 ( .A(n757), .Y(n136) );
  INVX1 U869 ( .A(n559), .Y(n116) );
  INVX1 U870 ( .A(b[5]), .Y(n784) );
  INVX1 U871 ( .A(n590), .Y(n94) );
  INVX1 U872 ( .A(b[6]), .Y(n786) );
  INVX1 U873 ( .A(n104), .Y(n103) );
endmodule


module alu_DW_mult_uns_24 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n26, n27, n28, n29, n33, n34, n35,
         n36, n41, n42, n43, n44, n45, n49, n50, n51, n52, n53, n57, n58, n59,
         n60, n61, n65, n66, n67, n68, n69, n73, n74, n75, n76, n77, n81, n82,
         n83, n84, n85, n87, n88, n89, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n105, n106, n110, n111, n115, n116, n117, n121,
         n122, n123, n124, n125, n129, n130, n131, n132, n133, n134, n138,
         n139, n155, n160, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n420, n421, n422, n423, n424, n425, n426, n427,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n462,
         n463, n465, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833;
  assign product[0] = b[0];

  FAX1 U2 ( .A(a[15]), .B(n675), .C(n26), .YC(product[31]), .YS(product[30])
         );
  FAX1 U3 ( .A(n719), .B(n164), .C(n27), .YC(n26), .YS(product[29]) );
  FAX1 U4 ( .A(n165), .B(n166), .C(n28), .YC(n27), .YS(product[28]) );
  FAX1 U5 ( .A(n167), .B(n168), .C(n139), .YC(n28), .YS(product[27]) );
  XNOR2X1 U7 ( .A(n778), .B(n715), .Y(product[26]) );
  AOI21X1 U8 ( .A(n551), .B(n787), .C(n33), .Y(n29) );
  XOR2X1 U15 ( .A(n631), .B(n608), .Y(product[25]) );
  OAI21X1 U16 ( .A(n762), .B(n575), .C(n744), .Y(n34) );
  XNOR2X1 U21 ( .A(n779), .B(n700), .Y(product[24]) );
  XOR2X1 U29 ( .A(n629), .B(n607), .Y(product[23]) );
  OAI21X1 U30 ( .A(n763), .B(n630), .C(n745), .Y(n42) );
  XNOR2X1 U35 ( .A(n565), .B(n693), .Y(product[22]) );
  AOI21X1 U36 ( .A(n50), .B(n780), .C(n49), .Y(n45) );
  XOR2X1 U43 ( .A(n559), .B(n606), .Y(product[21]) );
  OAI21X1 U44 ( .A(n576), .B(n764), .C(n746), .Y(n50) );
  XNOR2X1 U49 ( .A(n634), .B(n601), .Y(product[20]) );
  AOI21X1 U50 ( .A(n58), .B(n784), .C(n57), .Y(n53) );
  XOR2X1 U57 ( .A(n626), .B(n605), .Y(product[19]) );
  OAI21X1 U58 ( .A(n765), .B(n627), .C(n748), .Y(n58) );
  XNOR2X1 U63 ( .A(n564), .B(n714), .Y(product[18]) );
  AOI21X1 U64 ( .A(n66), .B(n783), .C(n65), .Y(n61) );
  XOR2X1 U71 ( .A(n557), .B(n604), .Y(product[17]) );
  OAI21X1 U72 ( .A(n766), .B(n579), .C(n747), .Y(n66) );
  XNOR2X1 U77 ( .A(n566), .B(n682), .Y(product[16]) );
  AOI21X1 U78 ( .A(n550), .B(n781), .C(n73), .Y(n69) );
  XOR2X1 U85 ( .A(n560), .B(n701), .Y(product[15]) );
  OAI21X1 U86 ( .A(n554), .B(n758), .C(n734), .Y(n74) );
  XNOR2X1 U91 ( .A(n552), .B(n600), .Y(product[14]) );
  AOI21X1 U92 ( .A(n549), .B(n782), .C(n81), .Y(n77) );
  XOR2X1 U99 ( .A(n593), .B(n603), .Y(product[13]) );
  OAI21X1 U100 ( .A(n574), .B(n578), .C(n586), .Y(n82) );
  AOI21X1 U102 ( .A(n799), .B(n85), .C(n88), .Y(n84) );
  XNOR2X1 U109 ( .A(n94), .B(n599), .Y(product[12]) );
  AOI21X1 U110 ( .A(n94), .B(n798), .C(n799), .Y(n89) );
  XNOR2X1 U117 ( .A(n100), .B(n674), .Y(product[11]) );
  AOI21X1 U119 ( .A(n567), .B(n590), .C(n589), .Y(n95) );
  XOR2X1 U126 ( .A(n103), .B(n728), .Y(product[10]) );
  OAI21X1 U127 ( .A(n777), .B(n103), .C(n759), .Y(n100) );
  XOR2X1 U132 ( .A(n592), .B(n602), .Y(product[9]) );
  AOI21X1 U136 ( .A(n790), .B(n115), .C(n110), .Y(n106) );
  XNOR2X1 U143 ( .A(n116), .B(n598), .Y(product[8]) );
  AOI21X1 U144 ( .A(n116), .B(n789), .C(n115), .Y(n111) );
  XNOR2X1 U151 ( .A(n568), .B(n597), .Y(product[7]) );
  AOI21X1 U153 ( .A(n122), .B(n792), .C(n121), .Y(n117) );
  XOR2X1 U160 ( .A(n595), .B(n633), .Y(product[6]) );
  OAI21X1 U161 ( .A(n618), .B(n633), .C(n615), .Y(n122) );
  XNOR2X1 U166 ( .A(n130), .B(n596), .Y(product[5]) );
  AOI21X1 U167 ( .A(n130), .B(n791), .C(n129), .Y(n125) );
  XOR2X1 U174 ( .A(n594), .B(n571), .Y(product[4]) );
  OAI21X1 U175 ( .A(n571), .B(n572), .C(n583), .Y(n130) );
  XNOR2X1 U180 ( .A(n134), .B(n138), .Y(product[3]) );
  FAX1 U190 ( .A(a[14]), .B(n624), .C(n614), .YC(n164), .YS(n165) );
  FAX1 U191 ( .A(n704), .B(n703), .C(n170), .YC(n166), .YS(n167) );
  FAX1 U192 ( .A(n683), .B(n174), .C(n171), .YC(n168), .YS(n169) );
  FAX1 U193 ( .A(a[13]), .B(n643), .C(n642), .YC(n170), .YS(n171) );
  FAX1 U194 ( .A(n180), .B(n175), .C(n178), .YC(n172), .YS(n173) );
  FAX1 U195 ( .A(n656), .B(n654), .C(n655), .YC(n174), .YS(n175) );
  FAX1 U196 ( .A(n181), .B(n184), .C(n179), .YC(n176), .YS(n177) );
  FAX1 U197 ( .A(n665), .B(n664), .C(n186), .YC(n178), .YS(n179) );
  FAX1 U198 ( .A(a[12]), .B(n636), .C(n635), .YC(n180), .YS(n181) );
  FAX1 U199 ( .A(n187), .B(n185), .C(n190), .YC(n182), .YS(n183) );
  FAX1 U200 ( .A(n720), .B(n194), .C(n192), .YC(n184), .YS(n185) );
  FAX1 U201 ( .A(n752), .B(n751), .C(n750), .YC(n186), .YS(n187) );
  FAX1 U202 ( .A(n200), .B(n191), .C(n198), .YC(n188), .YS(n189) );
  FAX1 U203 ( .A(n202), .B(n195), .C(n193), .YC(n190), .YS(n191) );
  FAX1 U204 ( .A(n645), .B(n646), .C(n644), .YC(n192), .YS(n193) );
  FAX1 U205 ( .A(a[11]), .B(n623), .C(n613), .YC(n194), .YS(n195) );
  FAX1 U206 ( .A(n208), .B(n199), .C(n206), .YC(n196), .YS(n197) );
  FAX1 U207 ( .A(n210), .B(n203), .C(n201), .YC(n198), .YS(n199) );
  FAX1 U208 ( .A(n666), .B(n667), .C(n212), .YC(n200), .YS(n201) );
  FAX1 U209 ( .A(n650), .B(n651), .C(n649), .YC(n202), .YS(n203) );
  FAX1 U210 ( .A(n209), .B(n216), .C(n207), .YC(n204), .YS(n205) );
  FAX1 U211 ( .A(n213), .B(n211), .C(n218), .YC(n206), .YS(n207) );
  FAX1 U212 ( .A(n697), .B(n222), .C(n220), .YC(n208), .YS(n209) );
  FAX1 U213 ( .A(n696), .B(n694), .C(n695), .YC(n210), .YS(n211) );
  FAX1 U214 ( .A(a[10]), .B(n638), .C(n637), .YC(n212), .YS(n213) );
  FAX1 U215 ( .A(n219), .B(n226), .C(n217), .YC(n214), .YS(n215) );
  FAX1 U216 ( .A(n223), .B(n230), .C(n228), .YC(n216), .YS(n217) );
  FAX1 U217 ( .A(n234), .B(n232), .C(n221), .YC(n218), .YS(n219) );
  FAX1 U218 ( .A(n686), .B(n684), .C(n685), .YC(n220), .YS(n221) );
  FAX1 U219 ( .A(n662), .B(n661), .C(n660), .YC(n222), .YS(n223) );
  FAX1 U220 ( .A(n229), .B(n238), .C(n227), .YC(n224), .YS(n225) );
  FAX1 U221 ( .A(n242), .B(n231), .C(n240), .YC(n226), .YS(n227) );
  FAX1 U222 ( .A(n244), .B(n235), .C(n233), .YC(n228), .YS(n229) );
  FAX1 U223 ( .A(n735), .B(n736), .C(n246), .YC(n230), .YS(n231) );
  FAX1 U224 ( .A(n673), .B(n672), .C(n671), .YC(n232), .YS(n233) );
  FAX1 U225 ( .A(a[9]), .B(n658), .C(n659), .YC(n234), .YS(n235) );
  FAX1 U226 ( .A(n241), .B(n250), .C(n239), .YC(n236), .YS(n237) );
  FAX1 U227 ( .A(n254), .B(n243), .C(n252), .YC(n238), .YS(n239) );
  FAX1 U228 ( .A(n256), .B(n247), .C(n245), .YC(n240), .YS(n241) );
  FAX1 U229 ( .A(n724), .B(n260), .C(n258), .YC(n242), .YS(n243) );
  FAX1 U230 ( .A(n706), .B(n708), .C(n707), .YC(n244), .YS(n245) );
  FAX1 U231 ( .A(n678), .B(n677), .C(n676), .YC(n246), .YS(n247) );
  FAX1 U232 ( .A(n253), .B(n264), .C(n251), .YC(n248), .YS(n249) );
  FAX1 U233 ( .A(n268), .B(n255), .C(n266), .YC(n250), .YS(n251) );
  FAX1 U234 ( .A(n270), .B(n259), .C(n257), .YC(n252), .YS(n253) );
  FAX1 U235 ( .A(n769), .B(n272), .C(n261), .YC(n254), .YS(n255) );
  FAX1 U236 ( .A(n771), .B(n770), .C(n772), .YC(n256), .YS(n257) );
  FAX1 U237 ( .A(n774), .B(n775), .C(n773), .YC(n258), .YS(n259) );
  HAX1 U238 ( .A(a[8]), .B(n668), .YC(n260), .YS(n261) );
  FAX1 U239 ( .A(n267), .B(n276), .C(n265), .YC(n262), .YS(n263) );
  FAX1 U240 ( .A(n271), .B(n269), .C(n278), .YC(n264), .YS(n265) );
  FAX1 U241 ( .A(n273), .B(n282), .C(n280), .YC(n266), .YS(n267) );
  FAX1 U242 ( .A(n754), .B(n753), .C(n284), .YC(n268), .YS(n269) );
  FAX1 U243 ( .A(n757), .B(n755), .C(n756), .YC(n270), .YS(n271) );
  HAX1 U244 ( .A(n648), .B(n647), .YC(n272), .YS(n273) );
  FAX1 U245 ( .A(n279), .B(n288), .C(n277), .YC(n274), .YS(n275) );
  FAX1 U246 ( .A(n283), .B(n281), .C(n290), .YC(n276), .YS(n277) );
  FAX1 U247 ( .A(n294), .B(n285), .C(n292), .YC(n278), .YS(n279) );
  FAX1 U248 ( .A(n738), .B(n739), .C(n737), .YC(n280), .YS(n281) );
  FAX1 U249 ( .A(n723), .B(n722), .C(n721), .YC(n282), .YS(n283) );
  HAX1 U250 ( .A(a[7]), .B(n727), .YC(n284), .YS(n285) );
  FAX1 U251 ( .A(n298), .B(n291), .C(n289), .YC(n286), .YS(n287) );
  FAX1 U252 ( .A(n302), .B(n293), .C(n300), .YC(n288), .YS(n289) );
  FAX1 U253 ( .A(n768), .B(n304), .C(n295), .YC(n290), .YS(n291) );
  FAX1 U254 ( .A(n711), .B(n710), .C(n709), .YC(n292), .YS(n293) );
  HAX1 U255 ( .A(n692), .B(n691), .YC(n294), .YS(n295) );
  FAX1 U256 ( .A(n301), .B(n621), .C(n299), .YC(n296), .YS(n297) );
  FAX1 U257 ( .A(n305), .B(n310), .C(n303), .YC(n298), .YS(n299) );
  FAX1 U258 ( .A(n699), .B(n698), .C(n312), .YC(n300), .YS(n301) );
  FAX1 U259 ( .A(n410), .B(n663), .C(n553), .YC(n302), .YS(n303) );
  HAX1 U260 ( .A(a[6]), .B(n690), .YC(n304), .YS(n305) );
  FAX1 U263 ( .A(n681), .B(n680), .C(n679), .YC(n310), .YS(n311) );
  HAX1 U264 ( .A(n657), .B(n555), .YC(n312), .YS(n313) );
  FAX1 U265 ( .A(n319), .B(n324), .C(n317), .YC(n314), .YS(n315) );
  FAX1 U266 ( .A(n767), .B(n321), .C(n788), .YC(n316), .YS(n317) );
  FAX1 U267 ( .A(n687), .B(n689), .C(n688), .YC(n318), .YS(n319) );
  HAX1 U268 ( .A(a[5]), .B(n726), .YC(n320), .YS(n321) );
  FAX1 U269 ( .A(n327), .B(n330), .C(n325), .YC(n322), .YS(n323) );
  FAX1 U270 ( .A(n452), .B(n639), .C(n332), .YC(n324), .YS(n325) );
  FAX1 U272 ( .A(n336), .B(n333), .C(n331), .YC(n328), .YS(n329) );
  FAX1 U273 ( .A(n712), .B(n653), .C(n652), .YC(n330), .YS(n331) );
  HAX1 U274 ( .A(a[4]), .B(n453), .YC(n332), .YS(n333) );
  FAX1 U275 ( .A(n705), .B(n340), .C(n337), .YC(n334), .YS(n335) );
  HAX1 U276 ( .A(n641), .B(n640), .YC(n336), .YS(n337) );
  FAX1 U277 ( .A(n670), .B(n669), .C(n342), .YC(n338), .YS(n339) );
  HAX1 U278 ( .A(a[3]), .B(n743), .YC(n340), .YS(n341) );
  HAX1 U279 ( .A(n713), .B(n793), .YC(n342), .YS(n343) );
  HAX1 U280 ( .A(a[2]), .B(n462), .YC(n344), .YS(n345) );
  INVX2 U434 ( .A(n83), .Y(n574) );
  INVX2 U435 ( .A(n398), .Y(n722) );
  OR2X2 U436 ( .A(n833), .B(n831), .Y(n347) );
  OR2X2 U437 ( .A(n833), .B(n829), .Y(n348) );
  OR2X2 U438 ( .A(n833), .B(n828), .Y(n349) );
  OR2X2 U439 ( .A(n833), .B(n826), .Y(n350) );
  OR2X2 U440 ( .A(n833), .B(n825), .Y(n351) );
  OR2X2 U441 ( .A(n833), .B(n821), .Y(n353) );
  OR2X2 U442 ( .A(n833), .B(n820), .Y(n354) );
  OR2X2 U443 ( .A(n833), .B(n819), .Y(n355) );
  INVX2 U444 ( .A(n433), .Y(n711) );
  XOR2X1 U445 ( .A(n806), .B(n309), .Y(n547) );
  INVX1 U446 ( .A(n547), .Y(n307) );
  INVX1 U447 ( .A(n547), .Y(n548) );
  OAI21X1 U448 ( .A(n574), .B(n578), .C(n586), .Y(n549) );
  OAI21X1 U449 ( .A(n554), .B(n758), .C(n734), .Y(n550) );
  OAI21X1 U450 ( .A(n762), .B(n575), .C(n744), .Y(n551) );
  OR2X2 U451 ( .A(n819), .B(n816), .Y(n794) );
  INVX8 U452 ( .A(b[3]), .Y(n816) );
  OR2X1 U453 ( .A(n826), .B(n816), .Y(n417) );
  OR2X2 U454 ( .A(n828), .B(n816), .Y(n407) );
  AND2X2 U455 ( .A(n573), .B(n582), .Y(n806) );
  AND2X2 U456 ( .A(n616), .B(n297), .Y(n799) );
  OR2X2 U457 ( .A(n297), .B(n616), .Y(n786) );
  OR2X2 U458 ( .A(n810), .B(n617), .Y(n616) );
  OR2X2 U459 ( .A(n812), .B(n811), .Y(n617) );
  AND2X2 U460 ( .A(n309), .B(n311), .Y(n811) );
  INVX4 U461 ( .A(n429), .Y(n689) );
  OR2X2 U462 ( .A(n824), .B(n813), .Y(n429) );
  AND2X2 U463 ( .A(n561), .B(n309), .Y(n812) );
  AND2X1 U464 ( .A(n563), .B(n801), .Y(n802) );
  OR2X1 U465 ( .A(n225), .B(n236), .Y(n783) );
  OR2X1 U466 ( .A(n249), .B(n262), .Y(n781) );
  INVX1 U467 ( .A(n632), .Y(n633) );
  OR2X1 U468 ( .A(n329), .B(n334), .Y(n789) );
  OR2X1 U469 ( .A(n832), .B(n821), .Y(n367) );
  OR2X1 U470 ( .A(n833), .B(n815), .Y(n358) );
  OR2X1 U471 ( .A(n825), .B(n822), .Y(n421) );
  OR2X1 U472 ( .A(n820), .B(n828), .Y(n404) );
  OR2X1 U473 ( .A(n814), .B(n831), .Y(n386) );
  OR2X1 U474 ( .A(n825), .B(n818), .Y(n425) );
  OR2X1 U475 ( .A(n826), .B(n829), .Y(n389) );
  OR2X1 U476 ( .A(n825), .B(n831), .Y(n378) );
  OR2X1 U477 ( .A(n832), .B(n820), .Y(n368) );
  OR2X1 U478 ( .A(n829), .B(n822), .Y(n391) );
  OR2X1 U479 ( .A(n821), .B(n831), .Y(n380) );
  OR2X1 U480 ( .A(n832), .B(n816), .Y(n371) );
  OR2X1 U481 ( .A(n820), .B(n831), .Y(n381) );
  OR2X1 U482 ( .A(n825), .B(n826), .Y(n411) );
  OR2X1 U483 ( .A(n833), .B(n816), .Y(n357) );
  OR2X1 U484 ( .A(n826), .B(n822), .Y(n412) );
  OR2X1 U485 ( .A(n821), .B(n828), .Y(n403) );
  OR2X1 U486 ( .A(n832), .B(n818), .Y(n370) );
  OR2X1 U487 ( .A(n820), .B(n829), .Y(n393) );
  OR2X1 U488 ( .A(n831), .B(n819), .Y(n382) );
  OR2X1 U489 ( .A(n831), .B(n818), .Y(n383) );
  OR2X1 U490 ( .A(n829), .B(n818), .Y(n395) );
  OR2X1 U491 ( .A(n821), .B(n825), .Y(n422) );
  OR2X1 U492 ( .A(n820), .B(n825), .Y(n423) );
  OR2X1 U493 ( .A(n826), .B(n818), .Y(n416) );
  OR2X1 U494 ( .A(n825), .B(n819), .Y(n424) );
  INVX1 U495 ( .A(n438), .Y(n721) );
  INVX1 U496 ( .A(n426), .Y(n710) );
  AND2X1 U497 ( .A(b[11]), .B(b[0]), .Y(n410) );
  OR2X1 U498 ( .A(n832), .B(n826), .Y(n364) );
  OR2X1 U499 ( .A(n828), .B(n831), .Y(n376) );
  OR2X1 U500 ( .A(n832), .B(n825), .Y(n365) );
  OR2X1 U501 ( .A(n831), .B(n826), .Y(n377) );
  OR2X1 U502 ( .A(n832), .B(n822), .Y(n366) );
  OR2X1 U503 ( .A(n828), .B(n822), .Y(n402) );
  INVX1 U504 ( .A(n414), .Y(n708) );
  INVX1 U505 ( .A(n373), .Y(n775) );
  OR2X1 U506 ( .A(n820), .B(n822), .Y(n431) );
  OR2X1 U507 ( .A(n821), .B(n822), .Y(n430) );
  OR2X1 U508 ( .A(n826), .B(n815), .Y(n418) );
  AND2X1 U509 ( .A(n313), .B(n558), .Y(n809) );
  INVX1 U510 ( .A(n440), .Y(n698) );
  INVX1 U511 ( .A(n427), .Y(n699) );
  OR2X1 U512 ( .A(n821), .B(n818), .Y(n440) );
  OR2X1 U513 ( .A(n819), .B(n818), .Y(n451) );
  INVX2 U514 ( .A(n436), .Y(n688) );
  OR2X1 U515 ( .A(n814), .B(n822), .Y(n436) );
  INVX2 U516 ( .A(n442), .Y(n687) );
  OR2X1 U517 ( .A(n821), .B(n815), .Y(n442) );
  OR2X1 U518 ( .A(n831), .B(n829), .Y(n375) );
  OR2X1 U519 ( .A(n832), .B(n819), .Y(n369) );
  AND2X1 U520 ( .A(n786), .B(n87), .Y(n83) );
  OR2X1 U521 ( .A(n287), .B(n296), .Y(n87) );
  OR2X1 U522 ( .A(n742), .B(n777), .Y(n96) );
  AND2X1 U523 ( .A(n789), .B(n790), .Y(n105) );
  OR2X1 U524 ( .A(n814), .B(n821), .Y(n443) );
  OR2X1 U525 ( .A(n823), .B(n813), .Y(n437) );
  AND2X1 U526 ( .A(b[5]), .B(b[2]), .Y(n453) );
  INVX1 U527 ( .A(n444), .Y(n653) );
  INVX1 U528 ( .A(b[6]), .Y(n820) );
  OR2X1 U529 ( .A(n818), .B(n815), .Y(n457) );
  OR2X1 U530 ( .A(n323), .B(n328), .Y(n790) );
  AND2X1 U531 ( .A(n341), .B(n339), .Y(n124) );
  OR2X1 U532 ( .A(n818), .B(n813), .Y(n459) );
  AND2X1 U533 ( .A(n733), .B(n783), .Y(n9) );
  AND2X1 U534 ( .A(n248), .B(n237), .Y(n68) );
  AND2X1 U535 ( .A(n717), .B(n781), .Y(n11) );
  AND2X1 U536 ( .A(n612), .B(n85), .Y(n14) );
  AND2X1 U537 ( .A(n718), .B(n155), .Y(n16) );
  AND2X1 U538 ( .A(n609), .B(n138), .Y(n133) );
  OR2X1 U539 ( .A(n345), .B(n620), .Y(n131) );
  AND2X1 U540 ( .A(n620), .B(n345), .Y(n132) );
  AND2X1 U541 ( .A(n795), .B(n776), .Y(product[2]) );
  AND2X1 U542 ( .A(n611), .B(n789), .Y(n19) );
  BUFX2 U543 ( .A(n82), .Y(n552) );
  AND2X1 U544 ( .A(n334), .B(n329), .Y(n115) );
  INVX2 U545 ( .A(b[7]), .Y(n821) );
  AND2X1 U546 ( .A(n338), .B(n335), .Y(n121) );
  OR2X1 U547 ( .A(n815), .B(n813), .Y(n134) );
  AND2X1 U548 ( .A(n563), .B(n561), .Y(n810) );
  AND2X1 U549 ( .A(n286), .B(n275), .Y(n81) );
  OR2X1 U550 ( .A(n315), .B(n322), .Y(n101) );
  AND2X1 U551 ( .A(n328), .B(n323), .Y(n110) );
  AND2X1 U552 ( .A(n322), .B(n315), .Y(n102) );
  AND2X1 U553 ( .A(n262), .B(n249), .Y(n73) );
  AND2X1 U554 ( .A(n236), .B(n225), .Y(n65) );
  OR2X1 U555 ( .A(n263), .B(n274), .Y(n75) );
  AND2X1 U556 ( .A(b[1]), .B(b[10]), .Y(n553) );
  INVX2 U557 ( .A(b[10]), .Y(n826) );
  INVX8 U558 ( .A(b[11]), .Y(n828) );
  OR2X1 U559 ( .A(n828), .B(n815), .Y(n408) );
  OR2X1 U560 ( .A(n817), .B(n815), .Y(n460) );
  INVX4 U561 ( .A(n794), .Y(n452) );
  INVX1 U562 ( .A(n75), .Y(n554) );
  INVX4 U563 ( .A(n441), .Y(n679) );
  AND2X2 U564 ( .A(b[1]), .B(b[9]), .Y(n555) );
  INVX1 U565 ( .A(b[9]), .Y(n824) );
  OR2X2 U566 ( .A(n829), .B(n816), .Y(n396) );
  INVX8 U567 ( .A(b[4]), .Y(n818) );
  INVX8 U568 ( .A(b[2]), .Y(n815) );
  OR2X2 U569 ( .A(n814), .B(n815), .Y(n463) );
  INVX1 U570 ( .A(n630), .Y(n556) );
  BUFX2 U571 ( .A(n579), .Y(n557) );
  FAX1 U572 ( .A(n687), .B(n689), .C(n688), .YC(n558), .YS() );
  INVX2 U573 ( .A(b[5]), .Y(n819) );
  INVX1 U574 ( .A(n320), .Y(n562) );
  OR2X2 U575 ( .A(n823), .B(n815), .Y(n435) );
  INVX2 U576 ( .A(b[12]), .Y(n829) );
  BUFX2 U577 ( .A(n576), .Y(n559) );
  BUFX2 U578 ( .A(n758), .Y(n560) );
  INVX1 U579 ( .A(n801), .Y(n561) );
  XNOR2X1 U580 ( .A(n313), .B(n562), .Y(n805) );
  FAX1 U581 ( .A(n681), .B(n680), .C(n679), .YC(), .YS(n563) );
  INVX8 U582 ( .A(n446), .Y(n680) );
  OR2X2 U583 ( .A(n832), .B(n831), .Y(n361) );
  OR2X2 U584 ( .A(n831), .B(n816), .Y(n384) );
  INVX8 U585 ( .A(b[13]), .Y(n831) );
  OR2X2 U586 ( .A(n820), .B(n819), .Y(n445) );
  INVX8 U587 ( .A(b[0]), .Y(n813) );
  OAI21X1 U588 ( .A(n766), .B(n557), .C(n747), .Y(n564) );
  OAI21X1 U589 ( .A(n559), .B(n764), .C(n746), .Y(n565) );
  BUFX2 U590 ( .A(n74), .Y(n566) );
  OAI21X1 U591 ( .A(n591), .B(n577), .C(n584), .Y(n567) );
  BUFX2 U592 ( .A(n122), .Y(n568) );
  INVX1 U593 ( .A(n627), .Y(n569) );
  OR2X2 U594 ( .A(n833), .B(n822), .Y(n352) );
  OR2X2 U595 ( .A(n831), .B(n822), .Y(n379) );
  OR2X2 U596 ( .A(n819), .B(n822), .Y(n432) );
  OR2X2 U597 ( .A(n816), .B(n822), .Y(n434) );
  OR2X2 U598 ( .A(n818), .B(n822), .Y(n433) );
  INVX2 U599 ( .A(n308), .Y(n621) );
  AND2X2 U600 ( .A(a[3]), .B(b[0]), .Y(n462) );
  AND2X2 U601 ( .A(b[1]), .B(a[1]), .Y(n570) );
  OR2X2 U602 ( .A(n814), .B(n813), .Y(n465) );
  AND2X2 U603 ( .A(n296), .B(n287), .Y(n88) );
  INVX8 U604 ( .A(b[8]), .Y(n822) );
  AND2X2 U605 ( .A(n580), .B(n622), .Y(n308) );
  AND2X2 U606 ( .A(n588), .B(n587), .Y(n622) );
  AND2X2 U607 ( .A(n102), .B(n98), .Y(n804) );
  AND2X2 U608 ( .A(n320), .B(n558), .Y(n808) );
  INVX1 U609 ( .A(n133), .Y(n571) );
  INVX1 U610 ( .A(n131), .Y(n572) );
  INVX1 U611 ( .A(n802), .Y(n573) );
  BUFX2 U612 ( .A(n619), .Y(n575) );
  BUFX2 U613 ( .A(n53), .Y(n576) );
  BUFX2 U614 ( .A(n117), .Y(n577) );
  BUFX2 U615 ( .A(n95), .Y(n578) );
  BUFX2 U616 ( .A(n69), .Y(n579) );
  INVX1 U617 ( .A(n809), .Y(n580) );
  INVX1 U618 ( .A(n804), .Y(n581) );
  AND2X2 U619 ( .A(n800), .B(n316), .Y(n803) );
  INVX1 U620 ( .A(n803), .Y(n582) );
  INVX1 U621 ( .A(n132), .Y(n583) );
  BUFX2 U622 ( .A(n106), .Y(n584) );
  INVX1 U623 ( .A(n84), .Y(n585) );
  INVX1 U624 ( .A(n585), .Y(n586) );
  INVX1 U625 ( .A(n808), .Y(n587) );
  AND2X2 U626 ( .A(n320), .B(n313), .Y(n807) );
  INVX1 U627 ( .A(n807), .Y(n588) );
  AND2X2 U628 ( .A(n581), .B(n718), .Y(n97) );
  INVX1 U629 ( .A(n97), .Y(n589) );
  INVX1 U630 ( .A(n96), .Y(n590) );
  INVX1 U631 ( .A(n105), .Y(n591) );
  BUFX2 U632 ( .A(n111), .Y(n592) );
  BUFX2 U633 ( .A(n89), .Y(n593) );
  AND2X1 U634 ( .A(n583), .B(n131), .Y(n23) );
  INVX1 U635 ( .A(n23), .Y(n594) );
  AND2X1 U636 ( .A(n615), .B(n160), .Y(n21) );
  INVX1 U637 ( .A(n21), .Y(n595) );
  AND2X1 U638 ( .A(n761), .B(n791), .Y(n22) );
  INVX1 U639 ( .A(n22), .Y(n596) );
  AND2X1 U640 ( .A(n610), .B(n792), .Y(n20) );
  INVX1 U641 ( .A(n20), .Y(n597) );
  INVX1 U642 ( .A(n19), .Y(n598) );
  AND2X1 U643 ( .A(n93), .B(n798), .Y(n15) );
  INVX1 U644 ( .A(n15), .Y(n599) );
  AND2X1 U645 ( .A(n716), .B(n782), .Y(n13) );
  INVX1 U646 ( .A(n13), .Y(n600) );
  AND2X1 U647 ( .A(n732), .B(n784), .Y(n7) );
  INVX1 U648 ( .A(n7), .Y(n601) );
  AND2X1 U649 ( .A(n702), .B(n790), .Y(n18) );
  INVX1 U650 ( .A(n18), .Y(n602) );
  INVX1 U651 ( .A(n14), .Y(n603) );
  AND2X1 U652 ( .A(n747), .B(n67), .Y(n10) );
  INVX1 U653 ( .A(n10), .Y(n604) );
  AND2X1 U654 ( .A(n748), .B(n59), .Y(n8) );
  INVX1 U655 ( .A(n8), .Y(n605) );
  AND2X1 U656 ( .A(n746), .B(n51), .Y(n6) );
  INVX1 U657 ( .A(n6), .Y(n606) );
  AND2X1 U658 ( .A(n745), .B(n43), .Y(n4) );
  INVX1 U659 ( .A(n4), .Y(n607) );
  AND2X1 U660 ( .A(n744), .B(n35), .Y(n2) );
  INVX1 U661 ( .A(n2), .Y(n608) );
  INVX1 U662 ( .A(n134), .Y(n609) );
  INVX1 U663 ( .A(n121), .Y(n610) );
  INVX1 U664 ( .A(n115), .Y(n611) );
  INVX1 U665 ( .A(n88), .Y(n612) );
  OR2X1 U666 ( .A(n825), .B(n829), .Y(n390) );
  INVX1 U667 ( .A(n390), .Y(n613) );
  INVX1 U668 ( .A(n348), .Y(n614) );
  INVX1 U669 ( .A(n124), .Y(n615) );
  OR2X1 U670 ( .A(n339), .B(n341), .Y(n123) );
  INVX1 U671 ( .A(n123), .Y(n618) );
  AOI21X1 U672 ( .A(n42), .B(n785), .C(n41), .Y(n619) );
  INVX1 U673 ( .A(n463), .Y(n620) );
  INVX1 U674 ( .A(n379), .Y(n623) );
  INVX1 U675 ( .A(n361), .Y(n624) );
  INVX1 U676 ( .A(n61), .Y(n625) );
  INVX1 U677 ( .A(n569), .Y(n626) );
  INVX1 U678 ( .A(n625), .Y(n627) );
  INVX1 U679 ( .A(n45), .Y(n628) );
  INVX1 U680 ( .A(n556), .Y(n629) );
  INVX1 U681 ( .A(n628), .Y(n630) );
  BUFX2 U682 ( .A(n575), .Y(n631) );
  INVX1 U683 ( .A(n125), .Y(n632) );
  BUFX2 U684 ( .A(n58), .Y(n634) );
  INVX1 U685 ( .A(b[14]), .Y(n832) );
  INVX1 U686 ( .A(n377), .Y(n635) );
  OR2X1 U687 ( .A(n828), .B(n829), .Y(n388) );
  INVX1 U688 ( .A(n388), .Y(n636) );
  OR2X2 U689 ( .A(n821), .B(n829), .Y(n392) );
  INVX1 U690 ( .A(n392), .Y(n637) );
  INVX1 U691 ( .A(n402), .Y(n638) );
  OR2X2 U692 ( .A(n820), .B(n815), .Y(n448) );
  INVX4 U693 ( .A(n448), .Y(n639) );
  OR2X1 U694 ( .A(n814), .B(n819), .Y(n454) );
  INVX1 U695 ( .A(n454), .Y(n640) );
  INVX1 U696 ( .A(n457), .Y(n641) );
  OR2X1 U697 ( .A(n832), .B(n828), .Y(n363) );
  INVX1 U698 ( .A(n363), .Y(n642) );
  INVX1 U699 ( .A(n375), .Y(n643) );
  INVX1 U700 ( .A(n354), .Y(n644) );
  OR2X1 U701 ( .A(n828), .B(n826), .Y(n400) );
  INVX1 U702 ( .A(n400), .Y(n645) );
  INVX1 U703 ( .A(n367), .Y(n646) );
  INVX1 U704 ( .A(n386), .Y(n647) );
  OR2X2 U705 ( .A(n830), .B(n815), .Y(n397) );
  INVX1 U706 ( .A(n397), .Y(n648) );
  INVX1 U707 ( .A(n355), .Y(n649) );
  INVX1 U708 ( .A(n391), .Y(n650) );
  INVX1 U709 ( .A(n368), .Y(n651) );
  OR2X2 U710 ( .A(n814), .B(n820), .Y(n449) );
  INVX1 U711 ( .A(n449), .Y(n652) );
  OR2X2 U712 ( .A(n821), .B(n813), .Y(n444) );
  INVX1 U713 ( .A(n376), .Y(n654) );
  INVX1 U714 ( .A(n351), .Y(n655) );
  INVX1 U715 ( .A(n364), .Y(n656) );
  INVX1 U716 ( .A(n435), .Y(n657) );
  INVX1 U717 ( .A(n383), .Y(n658) );
  OR2X1 U718 ( .A(n819), .B(n829), .Y(n394) );
  INVX1 U719 ( .A(n394), .Y(n659) );
  INVX1 U720 ( .A(n357), .Y(n660) );
  INVX1 U721 ( .A(n403), .Y(n661) );
  INVX1 U722 ( .A(n412), .Y(n662) );
  INVX1 U723 ( .A(n445), .Y(n663) );
  INVX1 U724 ( .A(n352), .Y(n664) );
  INVX1 U725 ( .A(n365), .Y(n665) );
  INVX1 U726 ( .A(n380), .Y(n666) );
  OR2X1 U727 ( .A(n825), .B(n828), .Y(n401) );
  INVX1 U728 ( .A(n401), .Y(n667) );
  INVX1 U729 ( .A(n396), .Y(n668) );
  OR2X1 U730 ( .A(n814), .B(n818), .Y(n458) );
  INVX1 U731 ( .A(n458), .Y(n669) );
  OR2X2 U732 ( .A(n819), .B(n813), .Y(n455) );
  INVX1 U733 ( .A(n455), .Y(n670) );
  INVX1 U734 ( .A(n358), .Y(n671) );
  INVX1 U735 ( .A(n404), .Y(n672) );
  INVX1 U736 ( .A(n421), .Y(n673) );
  INVX1 U737 ( .A(n16), .Y(n674) );
  OR2X2 U738 ( .A(n833), .B(n832), .Y(n346) );
  INVX1 U739 ( .A(n346), .Y(n675) );
  INVX2 U740 ( .A(b[15]), .Y(n833) );
  OR2X1 U741 ( .A(n833), .B(n814), .Y(n359) );
  INVX1 U742 ( .A(n359), .Y(n676) );
  INVX1 U743 ( .A(n422), .Y(n677) );
  INVX1 U744 ( .A(n395), .Y(n678) );
  OR2X2 U745 ( .A(n821), .B(n816), .Y(n441) );
  OR2X2 U746 ( .A(n820), .B(n818), .Y(n446) );
  OR2X2 U747 ( .A(n827), .B(n813), .Y(n420) );
  INVX4 U748 ( .A(n420), .Y(n681) );
  INVX1 U749 ( .A(n11), .Y(n682) );
  INVX1 U750 ( .A(n350), .Y(n683) );
  INVX1 U751 ( .A(n382), .Y(n684) );
  INVX1 U752 ( .A(n370), .Y(n685) );
  INVX1 U753 ( .A(n393), .Y(n686) );
  INVX1 U754 ( .A(n434), .Y(n690) );
  OR2X1 U755 ( .A(n814), .B(n828), .Y(n409) );
  INVX1 U756 ( .A(n409), .Y(n691) );
  OR2X2 U757 ( .A(n830), .B(n813), .Y(n399) );
  INVX1 U758 ( .A(n399), .Y(n692) );
  AND2X1 U759 ( .A(n731), .B(n780), .Y(n5) );
  INVX1 U760 ( .A(n5), .Y(n693) );
  INVX1 U761 ( .A(n381), .Y(n694) );
  OR2X1 U762 ( .A(n833), .B(n818), .Y(n356) );
  INVX1 U763 ( .A(n356), .Y(n695) );
  INVX1 U764 ( .A(n411), .Y(n696) );
  INVX1 U765 ( .A(n369), .Y(n697) );
  OR2X2 U766 ( .A(n824), .B(n815), .Y(n427) );
  AND2X1 U767 ( .A(n730), .B(n785), .Y(n3) );
  INVX1 U768 ( .A(n3), .Y(n700) );
  AND2X1 U769 ( .A(n734), .B(n75), .Y(n12) );
  INVX1 U770 ( .A(n12), .Y(n701) );
  INVX1 U771 ( .A(n110), .Y(n702) );
  INVX1 U772 ( .A(n349), .Y(n703) );
  OR2X1 U773 ( .A(n832), .B(n829), .Y(n362) );
  INVX1 U774 ( .A(n362), .Y(n704) );
  OR2X2 U775 ( .A(n820), .B(n813), .Y(n450) );
  INVX1 U776 ( .A(n450), .Y(n705) );
  INVX1 U777 ( .A(n384), .Y(n706) );
  OR2X2 U778 ( .A(n832), .B(n815), .Y(n372) );
  INVX1 U779 ( .A(n372), .Y(n707) );
  OR2X2 U780 ( .A(n820), .B(n826), .Y(n414) );
  OR2X2 U781 ( .A(n821), .B(n819), .Y(n439) );
  INVX1 U782 ( .A(n439), .Y(n709) );
  OR2X2 U783 ( .A(n824), .B(n816), .Y(n426) );
  OR2X1 U784 ( .A(n817), .B(n818), .Y(n456) );
  INVX1 U785 ( .A(n456), .Y(n712) );
  INVX1 U786 ( .A(n459), .Y(n713) );
  INVX1 U787 ( .A(n9), .Y(n714) );
  AND2X1 U788 ( .A(n729), .B(n787), .Y(n1) );
  INVX1 U789 ( .A(n1), .Y(n715) );
  INVX1 U790 ( .A(n81), .Y(n716) );
  INVX1 U791 ( .A(n73), .Y(n717) );
  AND2X2 U792 ( .A(n548), .B(n314), .Y(n99) );
  INVX1 U793 ( .A(n99), .Y(n718) );
  INVX1 U794 ( .A(n347), .Y(n719) );
  INVX1 U795 ( .A(n366), .Y(n720) );
  OR2X2 U796 ( .A(n821), .B(n820), .Y(n438) );
  OR2X1 U797 ( .A(n814), .B(n829), .Y(n398) );
  INVX1 U798 ( .A(n417), .Y(n723) );
  OR2X1 U799 ( .A(n828), .B(n819), .Y(n405) );
  INVX1 U800 ( .A(n405), .Y(n724) );
  INVX1 U801 ( .A(n437), .Y(n725) );
  INVX1 U802 ( .A(n451), .Y(n726) );
  INVX1 U803 ( .A(n432), .Y(n727) );
  AND2X1 U804 ( .A(n759), .B(n101), .Y(n17) );
  INVX1 U805 ( .A(n17), .Y(n728) );
  AND2X1 U806 ( .A(n169), .B(n172), .Y(n33) );
  INVX1 U807 ( .A(n33), .Y(n729) );
  AND2X1 U808 ( .A(n182), .B(n177), .Y(n41) );
  INVX1 U809 ( .A(n41), .Y(n730) );
  AND2X1 U810 ( .A(n189), .B(n196), .Y(n49) );
  INVX1 U811 ( .A(n49), .Y(n731) );
  AND2X1 U812 ( .A(n214), .B(n205), .Y(n57) );
  INVX1 U813 ( .A(n57), .Y(n732) );
  INVX1 U814 ( .A(n65), .Y(n733) );
  AND2X1 U815 ( .A(n274), .B(n263), .Y(n76) );
  INVX1 U816 ( .A(n76), .Y(n734) );
  OR2X1 U817 ( .A(n821), .B(n826), .Y(n413) );
  INVX1 U818 ( .A(n413), .Y(n735) );
  INVX1 U819 ( .A(n371), .Y(n736) );
  INVX1 U820 ( .A(n425), .Y(n737) );
  OR2X1 U821 ( .A(n831), .B(n813), .Y(n387) );
  INVX1 U822 ( .A(n387), .Y(n738) );
  INVX1 U823 ( .A(n408), .Y(n739) );
  INVX1 U824 ( .A(n443), .Y(n740) );
  INVX1 U825 ( .A(n443), .Y(n741) );
  AND2X2 U826 ( .A(n725), .B(n740), .Y(n788) );
  OR2X2 U827 ( .A(n307), .B(n314), .Y(n98) );
  INVX1 U828 ( .A(n98), .Y(n742) );
  INVX1 U829 ( .A(n460), .Y(n743) );
  AND2X1 U830 ( .A(n173), .B(n176), .Y(n36) );
  INVX1 U831 ( .A(n36), .Y(n744) );
  AND2X1 U832 ( .A(n183), .B(n188), .Y(n44) );
  INVX1 U833 ( .A(n44), .Y(n745) );
  AND2X1 U834 ( .A(n197), .B(n204), .Y(n52) );
  INVX1 U835 ( .A(n52), .Y(n746) );
  INVX1 U836 ( .A(n68), .Y(n747) );
  AND2X1 U837 ( .A(n224), .B(n215), .Y(n60) );
  INVX1 U838 ( .A(n60), .Y(n748) );
  INVX1 U839 ( .A(n465), .Y(n749) );
  OR2X2 U840 ( .A(n749), .B(a[1]), .Y(n795) );
  INVX1 U841 ( .A(n353), .Y(n750) );
  INVX1 U842 ( .A(n378), .Y(n751) );
  INVX1 U843 ( .A(n389), .Y(n752) );
  INVX1 U844 ( .A(n431), .Y(n753) );
  INVX1 U845 ( .A(n407), .Y(n754) );
  INVX1 U846 ( .A(n424), .Y(n755) );
  OR2X1 U847 ( .A(n832), .B(n813), .Y(n374) );
  INVX1 U848 ( .A(n374), .Y(n756) );
  INVX1 U849 ( .A(n416), .Y(n757) );
  BUFX2 U850 ( .A(n77), .Y(n758) );
  INVX1 U851 ( .A(n102), .Y(n759) );
  INVX1 U852 ( .A(n87), .Y(n760) );
  AND2X1 U853 ( .A(n344), .B(n343), .Y(n129) );
  INVX1 U854 ( .A(n129), .Y(n761) );
  OR2X1 U855 ( .A(n176), .B(n173), .Y(n35) );
  INVX1 U856 ( .A(n35), .Y(n762) );
  OR2X1 U857 ( .A(n188), .B(n183), .Y(n43) );
  INVX1 U858 ( .A(n43), .Y(n763) );
  OR2X1 U859 ( .A(n204), .B(n197), .Y(n51) );
  INVX1 U860 ( .A(n51), .Y(n764) );
  OR2X1 U861 ( .A(n215), .B(n224), .Y(n59) );
  INVX1 U862 ( .A(n59), .Y(n765) );
  OR2X1 U863 ( .A(n237), .B(n248), .Y(n67) );
  INVX1 U864 ( .A(n67), .Y(n766) );
  OR2X2 U865 ( .A(n820), .B(n816), .Y(n447) );
  INVX1 U866 ( .A(n447), .Y(n767) );
  INVX1 U867 ( .A(n418), .Y(n768) );
  INVX1 U868 ( .A(n430), .Y(n769) );
  OR2X1 U869 ( .A(n826), .B(n819), .Y(n415) );
  INVX1 U870 ( .A(n415), .Y(n770) );
  OR2X1 U871 ( .A(n828), .B(n818), .Y(n406) );
  INVX1 U872 ( .A(n406), .Y(n771) );
  INVX1 U873 ( .A(n423), .Y(n772) );
  OR2X1 U874 ( .A(n833), .B(n813), .Y(n360) );
  INVX1 U875 ( .A(n360), .Y(n773) );
  OR2X2 U876 ( .A(n831), .B(n815), .Y(n385) );
  INVX1 U877 ( .A(n385), .Y(n774) );
  OR2X1 U878 ( .A(n814), .B(n832), .Y(n373) );
  AND2X2 U879 ( .A(b[0]), .B(n570), .Y(n138) );
  INVX1 U880 ( .A(n138), .Y(n776) );
  INVX1 U881 ( .A(n101), .Y(n777) );
  BUFX2 U882 ( .A(n34), .Y(n778) );
  BUFX2 U883 ( .A(n42), .Y(n779) );
  INVX2 U884 ( .A(b[1]), .Y(n814) );
  OR2X1 U885 ( .A(n196), .B(n189), .Y(n780) );
  OR2X1 U886 ( .A(n275), .B(n286), .Y(n782) );
  OR2X1 U887 ( .A(n205), .B(n214), .Y(n784) );
  OR2X1 U888 ( .A(n177), .B(n182), .Y(n785) );
  OR2X1 U889 ( .A(n172), .B(n169), .Y(n787) );
  OR2X1 U890 ( .A(n343), .B(n344), .Y(n791) );
  INVX1 U891 ( .A(b[8]), .Y(n823) );
  INVX1 U892 ( .A(a[3]), .Y(n817) );
  INVX1 U893 ( .A(b[9]), .Y(n825) );
  INVX1 U894 ( .A(b[10]), .Y(n827) );
  INVX1 U895 ( .A(b[12]), .Y(n830) );
  OR2X1 U896 ( .A(n335), .B(n338), .Y(n792) );
  AND2X1 U897 ( .A(a[1]), .B(a[3]), .Y(n793) );
  INVX1 U898 ( .A(n567), .Y(n103) );
  INVX1 U899 ( .A(n786), .Y(n797) );
  INVX1 U900 ( .A(n797), .Y(n798) );
  INVX1 U901 ( .A(n799), .Y(n93) );
  INVX1 U902 ( .A(n618), .Y(n160) );
  INVX1 U903 ( .A(n311), .Y(n800) );
  INVX1 U904 ( .A(n316), .Y(n801) );
  XOR2X1 U905 ( .A(n725), .B(n741), .Y(n327) );
  INVX1 U906 ( .A(n760), .Y(n85) );
  XOR2X1 U907 ( .A(n805), .B(n318), .Y(n309) );
  INVX1 U908 ( .A(n577), .Y(n116) );
  INVX1 U909 ( .A(n578), .Y(n94) );
  INVX1 U910 ( .A(n742), .Y(n155) );
  INVX1 U911 ( .A(n29), .Y(n139) );
endmodule


module alu_DW_mult_uns_27 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n26, n27, n29, n33, n34, n35, n36,
         n37, n41, n42, n43, n44, n45, n49, n50, n51, n52, n53, n57, n58, n59,
         n60, n61, n65, n66, n67, n68, n69, n73, n74, n75, n76, n77, n81, n82,
         n83, n84, n86, n88, n89, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n110, n111, n115, n116, n117,
         n121, n122, n123, n124, n125, n129, n130, n131, n132, n133, n134,
         n136, n138, n139, n155, n156, n162, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n465, n547, n548, n549, n550,
         n551, n552, n553, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824;
  assign product[0] = b[0];

  FAX1 U2 ( .A(a[15]), .B(n750), .C(n26), .YC(product[31]), .YS(product[30])
         );
  FAX1 U3 ( .A(n772), .B(n164), .C(n27), .YC(n26), .YS(product[29]) );
  FAX1 U4 ( .A(n165), .B(n166), .C(n593), .YC(n27), .YS(product[28]) );
  XNOR2X1 U7 ( .A(n557), .B(n615), .Y(product[26]) );
  AOI21X1 U8 ( .A(n34), .B(n791), .C(n33), .Y(n29) );
  XOR2X1 U15 ( .A(n555), .B(n729), .Y(product[25]) );
  OAI21X1 U16 ( .A(n749), .B(n590), .C(n721), .Y(n34) );
  XNOR2X1 U21 ( .A(n582), .B(n763), .Y(product[24]) );
  AOI21X1 U22 ( .A(n42), .B(n793), .C(n41), .Y(n37) );
  XOR2X1 U29 ( .A(n579), .B(n623), .Y(product[23]) );
  OAI21X1 U30 ( .A(n767), .B(n589), .C(n732), .Y(n42) );
  XNOR2X1 U35 ( .A(n558), .B(n614), .Y(product[22]) );
  AOI21X1 U36 ( .A(n50), .B(n783), .C(n49), .Y(n45) );
  XOR2X1 U43 ( .A(n567), .B(n622), .Y(product[21]) );
  OAI21X1 U44 ( .A(n768), .B(n761), .C(n722), .Y(n50) );
  XNOR2X1 U49 ( .A(n559), .B(n613), .Y(product[20]) );
  AOI21X1 U50 ( .A(n58), .B(n785), .C(n57), .Y(n53) );
  XOR2X1 U57 ( .A(n805), .B(n621), .Y(product[19]) );
  OAI21X1 U58 ( .A(n769), .B(n592), .C(n733), .Y(n58) );
  XNOR2X1 U63 ( .A(n583), .B(n612), .Y(product[18]) );
  AOI21X1 U64 ( .A(n66), .B(n786), .C(n65), .Y(n61) );
  XOR2X1 U71 ( .A(n634), .B(n620), .Y(product[17]) );
  OAI21X1 U72 ( .A(n771), .B(n588), .C(n748), .Y(n66) );
  XNOR2X1 U77 ( .A(n581), .B(n611), .Y(product[16]) );
  AOI21X1 U78 ( .A(n74), .B(n784), .C(n73), .Y(n69) );
  XOR2X1 U85 ( .A(n578), .B(n619), .Y(product[15]) );
  OAI21X1 U86 ( .A(n770), .B(n760), .C(n734), .Y(n74) );
  XNOR2X1 U91 ( .A(n782), .B(n764), .Y(product[14]) );
  AOI21X1 U92 ( .A(n82), .B(n792), .C(n81), .Y(n77) );
  XOR2X1 U99 ( .A(n605), .B(n618), .Y(product[13]) );
  OAI21X1 U100 ( .A(n599), .B(n591), .C(n597), .Y(n82) );
  AOI21X1 U102 ( .A(n790), .B(n93), .C(n86), .Y(n84) );
  XNOR2X1 U109 ( .A(n94), .B(n610), .Y(product[12]) );
  AOI21X1 U110 ( .A(n94), .B(n789), .C(n93), .Y(n89) );
  XNOR2X1 U117 ( .A(n100), .B(n609), .Y(product[11]) );
  AOI21X1 U119 ( .A(n598), .B(n549), .C(n97), .Y(n95) );
  OAI21X1 U121 ( .A(n762), .B(n746), .C(n723), .Y(n97) );
  XOR2X1 U126 ( .A(n103), .B(n617), .Y(product[10]) );
  OAI21X1 U127 ( .A(n781), .B(n103), .C(n762), .Y(n100) );
  XOR2X1 U132 ( .A(n604), .B(n616), .Y(product[9]) );
  OAI21X1 U134 ( .A(n586), .B(n587), .C(n596), .Y(n104) );
  AOI21X1 U136 ( .A(n580), .B(n115), .C(n110), .Y(n106) );
  XNOR2X1 U143 ( .A(n116), .B(n608), .Y(product[8]) );
  AOI21X1 U144 ( .A(n116), .B(n584), .C(n115), .Y(n111) );
  XNOR2X1 U151 ( .A(n569), .B(n607), .Y(product[7]) );
  AOI21X1 U153 ( .A(n122), .B(n787), .C(n121), .Y(n117) );
  OAI21X1 U161 ( .A(n572), .B(n631), .C(n629), .Y(n122) );
  XNOR2X1 U166 ( .A(n602), .B(n570), .Y(product[5]) );
  AOI21X1 U167 ( .A(n130), .B(n788), .C(n129), .Y(n125) );
  XOR2X1 U174 ( .A(n606), .B(n635), .Y(product[4]) );
  OAI21X1 U175 ( .A(n635), .B(n632), .C(n628), .Y(n130) );
  XNOR2X1 U180 ( .A(n134), .B(n136), .Y(product[3]) );
  FAX1 U190 ( .A(a[14]), .B(n671), .C(n670), .YC(n164), .YS(n165) );
  FAX1 U191 ( .A(n697), .B(n696), .C(n170), .YC(n166), .YS(n167) );
  FAX1 U192 ( .A(n684), .B(n174), .C(n171), .YC(n168), .YS(n169) );
  FAX1 U193 ( .A(a[13]), .B(n737), .C(n736), .YC(n170), .YS(n171) );
  FAX1 U194 ( .A(n180), .B(n175), .C(n178), .YC(n172), .YS(n173) );
  FAX1 U195 ( .A(n700), .B(n699), .C(n698), .YC(n174), .YS(n175) );
  FAX1 U196 ( .A(n181), .B(n184), .C(n179), .YC(n176), .YS(n177) );
  FAX1 U197 ( .A(n739), .B(n738), .C(n186), .YC(n178), .YS(n179) );
  FAX1 U198 ( .A(a[12]), .B(n637), .C(n636), .YC(n180), .YS(n181) );
  FAX1 U199 ( .A(n187), .B(n185), .C(n190), .YC(n182), .YS(n183) );
  FAX1 U200 ( .A(n773), .B(n194), .C(n192), .YC(n184), .YS(n185) );
  FAX1 U201 ( .A(n726), .B(n725), .C(n724), .YC(n186), .YS(n187) );
  FAX1 U202 ( .A(n200), .B(n191), .C(n198), .YC(n188), .YS(n189) );
  FAX1 U203 ( .A(n202), .B(n195), .C(n193), .YC(n190), .YS(n191) );
  FAX1 U204 ( .A(n648), .B(n649), .C(n647), .YC(n192), .YS(n193) );
  FAX1 U205 ( .A(a[11]), .B(n633), .C(n627), .YC(n194), .YS(n195) );
  FAX1 U206 ( .A(n208), .B(n199), .C(n206), .YC(n196), .YS(n197) );
  FAX1 U207 ( .A(n210), .B(n203), .C(n201), .YC(n198), .YS(n199) );
  FAX1 U208 ( .A(n752), .B(n751), .C(n212), .YC(n200), .YS(n201) );
  FAX1 U209 ( .A(n642), .B(n641), .C(n640), .YC(n202), .YS(n203) );
  FAX1 U210 ( .A(n209), .B(n216), .C(n207), .YC(n204), .YS(n205) );
  FAX1 U211 ( .A(n213), .B(n211), .C(n218), .YC(n206), .YS(n207) );
  FAX1 U212 ( .A(n741), .B(n222), .C(n220), .YC(n208), .YS(n209) );
  FAX1 U213 ( .A(n662), .B(n663), .C(n661), .YC(n210), .YS(n211) );
  FAX1 U214 ( .A(a[10]), .B(n660), .C(n659), .YC(n212), .YS(n213) );
  FAX1 U215 ( .A(n219), .B(n226), .C(n217), .YC(n214), .YS(n215) );
  FAX1 U216 ( .A(n223), .B(n230), .C(n228), .YC(n216), .YS(n217) );
  FAX1 U217 ( .A(n234), .B(n232), .C(n221), .YC(n218), .YS(n219) );
  FAX1 U218 ( .A(n654), .B(n653), .C(n652), .YC(n220), .YS(n221) );
  FAX1 U219 ( .A(n675), .B(n676), .C(n674), .YC(n222), .YS(n223) );
  FAX1 U220 ( .A(n229), .B(n238), .C(n227), .YC(n224), .YS(n225) );
  FAX1 U221 ( .A(n242), .B(n231), .C(n240), .YC(n226), .YS(n227) );
  FAX1 U222 ( .A(n244), .B(n235), .C(n233), .YC(n228), .YS(n229) );
  FAX1 U223 ( .A(n774), .B(n775), .C(n246), .YC(n230), .YS(n231) );
  FAX1 U224 ( .A(n666), .B(n668), .C(n667), .YC(n232), .YS(n233) );
  FAX1 U225 ( .A(a[9]), .B(n683), .C(n682), .YC(n234), .YS(n235) );
  FAX1 U226 ( .A(n241), .B(n250), .C(n239), .YC(n236), .YS(n237) );
  FAX1 U227 ( .A(n254), .B(n243), .C(n252), .YC(n238), .YS(n239) );
  FAX1 U228 ( .A(n256), .B(n247), .C(n245), .YC(n240), .YS(n241) );
  FAX1 U229 ( .A(n779), .B(n260), .C(n258), .YC(n242), .YS(n243) );
  FAX1 U230 ( .A(n694), .B(n692), .C(n693), .YC(n244), .YS(n245) );
  FAX1 U231 ( .A(n679), .B(n677), .C(n678), .YC(n246), .YS(n247) );
  FAX1 U232 ( .A(n253), .B(n264), .C(n251), .YC(n248), .YS(n249) );
  FAX1 U233 ( .A(n268), .B(n255), .C(n266), .YC(n250), .YS(n251) );
  FAX1 U234 ( .A(n270), .B(n259), .C(n257), .YC(n252), .YS(n253) );
  FAX1 U235 ( .A(n753), .B(n272), .C(n261), .YC(n254), .YS(n255) );
  FAX1 U236 ( .A(n756), .B(n755), .C(n754), .YC(n256), .YS(n257) );
  FAX1 U237 ( .A(n759), .B(n758), .C(n757), .YC(n258), .YS(n259) );
  HAX1 U238 ( .A(a[8]), .B(n644), .YC(n260), .YS(n261) );
  FAX1 U239 ( .A(n267), .B(n276), .C(n265), .YC(n262), .YS(n263) );
  FAX1 U240 ( .A(n269), .B(n278), .C(n271), .YC(n264), .YS(n265) );
  FAX1 U241 ( .A(n273), .B(n282), .C(n280), .YC(n266), .YS(n267) );
  FAX1 U242 ( .A(n709), .B(n708), .C(n284), .YC(n268), .YS(n269) );
  FAX1 U243 ( .A(n714), .B(n712), .C(n713), .YC(n270), .YS(n271) );
  HAX1 U244 ( .A(n657), .B(n658), .YC(n272), .YS(n273) );
  FAX1 U245 ( .A(n279), .B(n288), .C(n277), .YC(n274), .YS(n275) );
  FAX1 U246 ( .A(n290), .B(n281), .C(n283), .YC(n276), .YS(n277) );
  FAX1 U247 ( .A(n294), .B(n285), .C(n292), .YC(n278), .YS(n279) );
  FAX1 U248 ( .A(n743), .B(n744), .C(n742), .YC(n280), .YS(n281) );
  FAX1 U249 ( .A(n778), .B(n777), .C(n776), .YC(n282), .YS(n283) );
  HAX1 U250 ( .A(a[7]), .B(n695), .YC(n284), .YS(n285) );
  FAX1 U251 ( .A(n298), .B(n291), .C(n289), .YC(n286), .YS(n287) );
  FAX1 U252 ( .A(n302), .B(n293), .C(n300), .YC(n288), .YS(n289) );
  FAX1 U253 ( .A(n704), .B(n304), .C(n295), .YC(n290), .YS(n291) );
  FAX1 U254 ( .A(n806), .B(n639), .C(n638), .YC(n292), .YS(n293) );
  HAX1 U255 ( .A(n651), .B(n650), .YC(n294), .YS(n295) );
  FAX1 U256 ( .A(n301), .B(n308), .C(n299), .YC(n296), .YS(n297) );
  FAX1 U257 ( .A(n305), .B(n310), .C(n303), .YC(n298), .YS(n299) );
  FAX1 U258 ( .A(n710), .B(n711), .C(n312), .YC(n300), .YS(n301) );
  FAX1 U259 ( .A(n728), .B(n727), .C(n571), .YC(n302), .YS(n303) );
  HAX1 U260 ( .A(a[6]), .B(n717), .YC(n304), .YS(n305) );
  FAX1 U261 ( .A(n311), .B(n316), .C(n309), .YC(n306), .YS(n307) );
  FAX1 U262 ( .A(n320), .B(n313), .C(n318), .YC(n308), .YS(n309) );
  FAX1 U263 ( .A(n703), .B(n702), .C(n701), .YC(n310), .YS(n311) );
  HAX1 U264 ( .A(n646), .B(n645), .YC(n312), .YS(n313) );
  FAX1 U265 ( .A(n319), .B(n324), .C(n317), .YC(n314), .YS(n315) );
  FAX1 U266 ( .A(n688), .B(n321), .C(n326), .YC(n316), .YS(n317) );
  FAX1 U267 ( .A(n685), .B(n687), .C(n686), .YC(n318), .YS(n319) );
  HAX1 U268 ( .A(n573), .B(n716), .YC(n320), .YS(n321) );
  FAX1 U269 ( .A(n327), .B(n330), .C(n325), .YC(n322), .YS(n323) );
  FAX1 U270 ( .A(n681), .B(n680), .C(n803), .YC(n324), .YS(n325) );
  HAX1 U271 ( .A(n664), .B(n665), .YC(n326), .YS(n327) );
  FAX1 U272 ( .A(n336), .B(n333), .C(n331), .YC(n328), .YS(n329) );
  FAX1 U273 ( .A(n691), .B(n690), .C(n689), .YC(n330), .YS(n331) );
  FAX1 U275 ( .A(n740), .B(n340), .C(n337), .YC(n334), .YS(n335) );
  HAX1 U276 ( .A(n601), .B(n600), .YC(n336), .YS(n337) );
  FAX1 U277 ( .A(n673), .B(n672), .C(n342), .YC(n338), .YS(n339) );
  HAX1 U278 ( .A(a[3]), .B(n715), .YC(n340), .YS(n341) );
  HAX1 U279 ( .A(n655), .B(n656), .YC(n342), .YS(n343) );
  HAX1 U280 ( .A(a[2]), .B(n643), .YC(n344), .YS(n345) );
  BUFX2 U434 ( .A(n139), .Y(n547) );
  INVX4 U435 ( .A(b[5]), .Y(n548) );
  INVX4 U436 ( .A(b[5]), .Y(n565) );
  OR2X2 U437 ( .A(n808), .B(n548), .Y(n454) );
  OR2X2 U438 ( .A(n548), .B(n566), .Y(n432) );
  OR2X2 U439 ( .A(n548), .B(n811), .Y(n451) );
  OR2X2 U440 ( .A(n814), .B(n548), .Y(n439) );
  OAI21X1 U441 ( .A(n586), .B(n587), .C(n596), .Y(n549) );
  INVX2 U442 ( .A(n105), .Y(n586) );
  INVX8 U443 ( .A(b[1]), .Y(n808) );
  INVX1 U444 ( .A(n813), .Y(n550) );
  INVX1 U445 ( .A(n550), .Y(n551) );
  INVX1 U446 ( .A(n550), .Y(n552) );
  INVX1 U447 ( .A(n550), .Y(n553) );
  INVX2 U448 ( .A(n449), .Y(n689) );
  INVX1 U449 ( .A(b[11]), .Y(n563) );
  OR2X1 U450 ( .A(n563), .B(n812), .Y(n405) );
  OR2X1 U451 ( .A(n814), .B(n810), .Y(n441) );
  OR2X1 U452 ( .A(n565), .B(n810), .Y(n452) );
  OR2X1 U453 ( .A(n563), .B(n810), .Y(n407) );
  INVX1 U454 ( .A(n447), .Y(n688) );
  AND2X1 U455 ( .A(n585), .B(n796), .Y(product[2]) );
  OR2X1 U456 ( .A(n824), .B(n568), .Y(n354) );
  OR2X1 U457 ( .A(n823), .B(n814), .Y(n367) );
  OR2X1 U458 ( .A(n563), .B(n818), .Y(n400) );
  OR2X1 U459 ( .A(n822), .B(n566), .Y(n379) );
  OR2X1 U460 ( .A(n824), .B(n812), .Y(n355) );
  OR2X1 U461 ( .A(n823), .B(n568), .Y(n368) );
  OR2X1 U462 ( .A(n820), .B(n566), .Y(n391) );
  OR2X1 U463 ( .A(n814), .B(n820), .Y(n392) );
  OR2X1 U464 ( .A(n824), .B(n811), .Y(n356) );
  OR2X1 U465 ( .A(n568), .B(n822), .Y(n381) );
  OR2X1 U466 ( .A(n816), .B(n818), .Y(n411) );
  OR2X1 U467 ( .A(n823), .B(n811), .Y(n370) );
  OR2X1 U468 ( .A(n822), .B(n812), .Y(n382) );
  OR2X1 U469 ( .A(n568), .B(n820), .Y(n393) );
  OR2X1 U470 ( .A(n818), .B(n566), .Y(n412) );
  OR2X1 U471 ( .A(n814), .B(n563), .Y(n403) );
  OR2X1 U472 ( .A(n568), .B(n563), .Y(n404) );
  OR2X1 U473 ( .A(n816), .B(n566), .Y(n421) );
  OR2X1 U474 ( .A(n823), .B(n809), .Y(n372) );
  OR2X1 U475 ( .A(n822), .B(n810), .Y(n384) );
  OR2X1 U476 ( .A(n568), .B(n818), .Y(n414) );
  OR2X1 U477 ( .A(n824), .B(n808), .Y(n359) );
  OR2X1 U478 ( .A(n820), .B(n811), .Y(n395) );
  OR2X1 U479 ( .A(n814), .B(n816), .Y(n422) );
  OR2X1 U480 ( .A(n822), .B(n809), .Y(n385) );
  OR2X1 U481 ( .A(n568), .B(n816), .Y(n423) );
  OR2X1 U482 ( .A(n818), .B(n812), .Y(n415) );
  OR2X1 U483 ( .A(n563), .B(n811), .Y(n406) );
  OR2X1 U484 ( .A(n815), .B(n809), .Y(n435) );
  OR2X1 U485 ( .A(n824), .B(n814), .Y(n353) );
  OR2X1 U486 ( .A(n816), .B(n822), .Y(n378) );
  OR2X1 U487 ( .A(n818), .B(n820), .Y(n389) );
  OR2X1 U488 ( .A(n814), .B(n818), .Y(n413) );
  OR2X1 U489 ( .A(n812), .B(n820), .Y(n394) );
  OR2X1 U490 ( .A(n568), .B(n566), .Y(n431) );
  OR2X1 U491 ( .A(n823), .B(n807), .Y(n374) );
  OR2X1 U492 ( .A(n818), .B(n811), .Y(n416) );
  OR2X1 U493 ( .A(n816), .B(n812), .Y(n424) );
  OR2X1 U494 ( .A(n821), .B(n807), .Y(n399) );
  OR2X1 U495 ( .A(n818), .B(n810), .Y(n417) );
  OR2X1 U496 ( .A(n563), .B(n809), .Y(n408) );
  OR2X1 U497 ( .A(n816), .B(n811), .Y(n425) );
  INVX1 U498 ( .A(n373), .Y(n758) );
  OR2X1 U499 ( .A(n562), .B(n807), .Y(n437) );
  OR2X1 U500 ( .A(n823), .B(n818), .Y(n364) );
  OR2X1 U501 ( .A(n824), .B(n816), .Y(n351) );
  OR2X1 U502 ( .A(n563), .B(n822), .Y(n376) );
  OR2X1 U503 ( .A(n823), .B(n563), .Y(n363) );
  OR2X1 U504 ( .A(n823), .B(n816), .Y(n365) );
  OR2X1 U505 ( .A(n563), .B(n820), .Y(n388) );
  OR2X1 U506 ( .A(n823), .B(n566), .Y(n366) );
  OR2X1 U507 ( .A(n816), .B(n563), .Y(n401) );
  OR2X1 U508 ( .A(n823), .B(n812), .Y(n369) );
  OR2X1 U509 ( .A(n821), .B(n809), .Y(n397) );
  AND2X1 U510 ( .A(b[11]), .B(a[0]), .Y(n571) );
  INVX2 U511 ( .A(n419), .Y(n728) );
  INVX1 U512 ( .A(n426), .Y(n639) );
  INVX1 U513 ( .A(n439), .Y(n638) );
  INVX2 U514 ( .A(n387), .Y(n778) );
  OR2X1 U515 ( .A(n818), .B(n809), .Y(n418) );
  OR2X1 U516 ( .A(n814), .B(n811), .Y(n440) );
  INVX2 U517 ( .A(n420), .Y(n703) );
  INVX1 U518 ( .A(n452), .Y(n681) );
  INVX1 U519 ( .A(n448), .Y(n680) );
  INVX1 U520 ( .A(n456), .Y(n691) );
  INVX1 U521 ( .A(b[6]), .Y(n813) );
  OR2X1 U522 ( .A(n811), .B(n807), .Y(n459) );
  OR2X1 U523 ( .A(n824), .B(n820), .Y(n348) );
  OR2X1 U524 ( .A(n824), .B(n563), .Y(n349) );
  OR2X1 U525 ( .A(n745), .B(n781), .Y(n96) );
  AND2X1 U526 ( .A(n794), .B(n795), .Y(n105) );
  INVX1 U527 ( .A(n458), .Y(n672) );
  INVX1 U528 ( .A(n455), .Y(n673) );
  OR2X1 U529 ( .A(n808), .B(n811), .Y(n458) );
  OR2X1 U530 ( .A(n824), .B(n818), .Y(n350) );
  AND2X1 U531 ( .A(n224), .B(n215), .Y(n60) );
  AND2X1 U532 ( .A(n248), .B(n237), .Y(n68) );
  OR2X1 U533 ( .A(n345), .B(n669), .Y(n131) );
  AND2X1 U534 ( .A(n669), .B(n345), .Y(n132) );
  OR2X1 U535 ( .A(n824), .B(n822), .Y(n347) );
  AND2X1 U536 ( .A(n721), .B(n35), .Y(n2) );
  AND2X1 U537 ( .A(n705), .B(n793), .Y(n3) );
  AND2X1 U538 ( .A(n274), .B(n263), .Y(n76) );
  AND2X1 U539 ( .A(n718), .B(n792), .Y(n13) );
  AND2X1 U540 ( .A(n766), .B(n789), .Y(n15) );
  AND2X1 U541 ( .A(n730), .B(n580), .Y(n18) );
  AND2X1 U542 ( .A(n747), .B(n584), .Y(n19) );
  INVX1 U543 ( .A(n133), .Y(n635) );
  OR2X2 U544 ( .A(n814), .B(n566), .Y(n430) );
  INVX8 U545 ( .A(b[3]), .Y(n810) );
  AND2X1 U546 ( .A(n306), .B(n297), .Y(n93) );
  INVX2 U547 ( .A(b[4]), .Y(n811) );
  OR2X1 U548 ( .A(n809), .B(n807), .Y(n134) );
  INVX1 U549 ( .A(b[11]), .Y(n819) );
  AND2X1 U550 ( .A(b[4]), .B(a[8]), .Y(n806) );
  INVX1 U551 ( .A(n75), .Y(n770) );
  OR2X1 U552 ( .A(n263), .B(n274), .Y(n75) );
  INVX1 U553 ( .A(n67), .Y(n771) );
  INVX2 U554 ( .A(b[0]), .Y(n807) );
  INVX2 U555 ( .A(b[7]), .Y(n814) );
  AND2X1 U556 ( .A(n328), .B(n577), .Y(n110) );
  OR2X1 U557 ( .A(n315), .B(n322), .Y(n101) );
  AND2X1 U558 ( .A(n262), .B(n249), .Y(n73) );
  AND2X1 U559 ( .A(n286), .B(n275), .Y(n81) );
  OR2X1 U560 ( .A(n339), .B(n341), .Y(n123) );
  OR2X1 U561 ( .A(n565), .B(n809), .Y(n453) );
  BUFX2 U562 ( .A(n590), .Y(n555) );
  OR2X2 U563 ( .A(n237), .B(n248), .Y(n67) );
  OR2X2 U564 ( .A(n808), .B(n823), .Y(n373) );
  AND2X1 U565 ( .A(a[1]), .B(n735), .Y(n138) );
  BUFX2 U566 ( .A(n547), .Y(n556) );
  OAI21X1 U567 ( .A(n749), .B(n555), .C(n721), .Y(n557) );
  OAI21X1 U568 ( .A(n768), .B(n761), .C(n722), .Y(n558) );
  OAI21X1 U569 ( .A(n769), .B(n592), .C(n733), .Y(n559) );
  INVX1 U570 ( .A(b[8]), .Y(n560) );
  INVX1 U571 ( .A(b[10]), .Y(n561) );
  INVX1 U572 ( .A(b[8]), .Y(n562) );
  INVX1 U573 ( .A(n446), .Y(n702) );
  INVX1 U574 ( .A(n453), .Y(n564) );
  BUFX2 U575 ( .A(n562), .Y(n566) );
  BUFX2 U576 ( .A(n761), .Y(n567) );
  INVX2 U577 ( .A(n436), .Y(n686) );
  INVX1 U578 ( .A(b[10]), .Y(n817) );
  INVX2 U579 ( .A(b[10]), .Y(n818) );
  OR2X2 U580 ( .A(n814), .B(n822), .Y(n380) );
  OR2X2 U581 ( .A(n808), .B(n822), .Y(n386) );
  OR2X2 U582 ( .A(n560), .B(n808), .Y(n436) );
  AND2X2 U583 ( .A(n322), .B(n315), .Y(n102) );
  INVX1 U584 ( .A(a[6]), .Y(n568) );
  BUFX2 U585 ( .A(n122), .Y(n569) );
  BUFX2 U586 ( .A(n130), .Y(n570) );
  OR2X2 U587 ( .A(n808), .B(n552), .Y(n449) );
  INVX1 U588 ( .A(n573), .Y(n812) );
  INVX2 U589 ( .A(n429), .Y(n687) );
  INVX1 U590 ( .A(n123), .Y(n572) );
  INVX1 U591 ( .A(n374), .Y(n713) );
  OR2X2 U592 ( .A(n816), .B(n807), .Y(n429) );
  OR2X2 U593 ( .A(n808), .B(n816), .Y(n428) );
  OR2X2 U594 ( .A(n810), .B(n807), .Y(n462) );
  INVX1 U595 ( .A(n548), .Y(n573) );
  INVX2 U596 ( .A(b[12]), .Y(n820) );
  OR2X2 U597 ( .A(n297), .B(n306), .Y(n789) );
  INVX1 U598 ( .A(n287), .Y(n574) );
  INVX1 U599 ( .A(n574), .Y(n575) );
  INVX1 U600 ( .A(n323), .Y(n576) );
  INVX1 U601 ( .A(n576), .Y(n577) );
  BUFX2 U602 ( .A(n760), .Y(n578) );
  BUFX2 U603 ( .A(n589), .Y(n579) );
  BUFX2 U604 ( .A(n795), .Y(n580) );
  OR2X2 U605 ( .A(n552), .B(n548), .Y(n445) );
  OAI21X1 U606 ( .A(n770), .B(n578), .C(n734), .Y(n581) );
  OAI21X1 U607 ( .A(n767), .B(n579), .C(n732), .Y(n582) );
  OAI21X1 U608 ( .A(n771), .B(n588), .C(n748), .Y(n583) );
  OR2X2 U609 ( .A(n824), .B(n807), .Y(n360) );
  BUFX2 U610 ( .A(n794), .Y(n584) );
  OR2X2 U611 ( .A(n808), .B(n807), .Y(n465) );
  OR2X2 U612 ( .A(n824), .B(n823), .Y(n346) );
  OR2X2 U613 ( .A(n823), .B(n810), .Y(n371) );
  INVX8 U614 ( .A(b[14]), .Y(n823) );
  OR2X1 U615 ( .A(n810), .B(n811), .Y(n456) );
  OR2X2 U616 ( .A(n329), .B(n334), .Y(n794) );
  AND2X2 U617 ( .A(n731), .B(n790), .Y(n14) );
  OR2X2 U618 ( .A(n814), .B(n552), .Y(n438) );
  OR2X2 U619 ( .A(n553), .B(n807), .Y(n450) );
  INVX8 U620 ( .A(b[9]), .Y(n816) );
  INVX1 U621 ( .A(b[12]), .Y(n821) );
  INVX8 U622 ( .A(b[2]), .Y(n809) );
  OR2X2 U623 ( .A(n323), .B(n328), .Y(n795) );
  OR2X2 U624 ( .A(n561), .B(n807), .Y(n420) );
  OR2X2 U625 ( .A(n808), .B(n817), .Y(n419) );
  OR2X2 U626 ( .A(n287), .B(n296), .Y(n790) );
  OR2X2 U627 ( .A(n594), .B(n800), .Y(n593) );
  OR2X2 U628 ( .A(n801), .B(n802), .Y(n594) );
  AND2X2 U629 ( .A(n167), .B(n547), .Y(n800) );
  AND2X2 U630 ( .A(n168), .B(n139), .Y(n801) );
  AND2X2 U631 ( .A(a[4]), .B(n564), .Y(n803) );
  INVX1 U632 ( .A(n138), .Y(n585) );
  AND2X2 U633 ( .A(n789), .B(n790), .Y(n83) );
  BUFX2 U634 ( .A(n117), .Y(n587) );
  BUFX2 U635 ( .A(n69), .Y(n588) );
  BUFX2 U636 ( .A(n45), .Y(n589) );
  BUFX2 U637 ( .A(n37), .Y(n590) );
  BUFX2 U638 ( .A(n95), .Y(n591) );
  BUFX2 U639 ( .A(n61), .Y(n592) );
  INVX1 U640 ( .A(n106), .Y(n595) );
  INVX1 U641 ( .A(n595), .Y(n596) );
  BUFX2 U642 ( .A(n84), .Y(n597) );
  INVX1 U643 ( .A(n96), .Y(n598) );
  INVX1 U644 ( .A(n83), .Y(n599) );
  AND2X1 U645 ( .A(n168), .B(n167), .Y(n802) );
  INVX1 U646 ( .A(n454), .Y(n600) );
  OR2X1 U647 ( .A(n811), .B(n809), .Y(n457) );
  INVX1 U648 ( .A(n457), .Y(n601) );
  AND2X1 U649 ( .A(n625), .B(n788), .Y(n22) );
  INVX1 U650 ( .A(n22), .Y(n602) );
  AND2X1 U651 ( .A(n629), .B(n630), .Y(n21) );
  INVX1 U652 ( .A(n21), .Y(n603) );
  BUFX2 U653 ( .A(n111), .Y(n604) );
  BUFX2 U654 ( .A(n89), .Y(n605) );
  AND2X1 U655 ( .A(n628), .B(n162), .Y(n23) );
  INVX1 U656 ( .A(n23), .Y(n606) );
  AND2X1 U657 ( .A(n626), .B(n787), .Y(n20) );
  INVX1 U658 ( .A(n20), .Y(n607) );
  INVX1 U659 ( .A(n19), .Y(n608) );
  AND2X1 U660 ( .A(n723), .B(n155), .Y(n16) );
  INVX1 U661 ( .A(n16), .Y(n609) );
  INVX1 U662 ( .A(n15), .Y(n610) );
  AND2X1 U663 ( .A(n720), .B(n784), .Y(n11) );
  INVX1 U664 ( .A(n11), .Y(n611) );
  AND2X1 U665 ( .A(n719), .B(n786), .Y(n9) );
  INVX1 U666 ( .A(n9), .Y(n612) );
  AND2X1 U667 ( .A(n707), .B(n785), .Y(n7) );
  INVX1 U668 ( .A(n7), .Y(n613) );
  AND2X1 U669 ( .A(n706), .B(n783), .Y(n5) );
  INVX1 U670 ( .A(n5), .Y(n614) );
  AND2X1 U671 ( .A(n765), .B(n791), .Y(n1) );
  INVX1 U672 ( .A(n1), .Y(n615) );
  INVX1 U673 ( .A(n18), .Y(n616) );
  AND2X1 U674 ( .A(n762), .B(n156), .Y(n17) );
  INVX1 U675 ( .A(n17), .Y(n617) );
  INVX1 U676 ( .A(n14), .Y(n618) );
  AND2X1 U677 ( .A(n734), .B(n75), .Y(n12) );
  INVX1 U678 ( .A(n12), .Y(n619) );
  AND2X1 U679 ( .A(n748), .B(n67), .Y(n10) );
  INVX1 U680 ( .A(n10), .Y(n620) );
  AND2X1 U681 ( .A(n733), .B(n59), .Y(n8) );
  INVX1 U682 ( .A(n8), .Y(n621) );
  AND2X1 U683 ( .A(n722), .B(n51), .Y(n6) );
  INVX1 U684 ( .A(n6), .Y(n622) );
  AND2X1 U685 ( .A(n732), .B(n43), .Y(n4) );
  INVX1 U686 ( .A(n4), .Y(n623) );
  INVX1 U687 ( .A(n134), .Y(n624) );
  AND2X1 U688 ( .A(n344), .B(n343), .Y(n129) );
  INVX1 U689 ( .A(n129), .Y(n625) );
  AND2X1 U690 ( .A(n338), .B(n335), .Y(n121) );
  INVX1 U691 ( .A(n121), .Y(n626) );
  OR2X1 U692 ( .A(n816), .B(n820), .Y(n390) );
  INVX1 U693 ( .A(n390), .Y(n627) );
  INVX1 U694 ( .A(n132), .Y(n628) );
  AND2X1 U695 ( .A(n341), .B(n339), .Y(n124) );
  INVX1 U696 ( .A(n124), .Y(n629) );
  INVX1 U697 ( .A(n572), .Y(n630) );
  BUFX2 U698 ( .A(n125), .Y(n631) );
  INVX1 U699 ( .A(n131), .Y(n632) );
  INVX1 U700 ( .A(n379), .Y(n633) );
  BUFX2 U701 ( .A(n588), .Y(n634) );
  AND2X2 U702 ( .A(n624), .B(n138), .Y(n133) );
  OR2X2 U703 ( .A(n822), .B(n818), .Y(n377) );
  INVX1 U704 ( .A(n377), .Y(n636) );
  INVX1 U705 ( .A(n388), .Y(n637) );
  OR2X2 U706 ( .A(n816), .B(n810), .Y(n426) );
  INVX1 U707 ( .A(n355), .Y(n640) );
  INVX1 U708 ( .A(n368), .Y(n641) );
  INVX1 U709 ( .A(n391), .Y(n642) );
  INVX1 U710 ( .A(n462), .Y(n643) );
  INVX1 U711 ( .A(n385), .Y(n644) );
  INVX1 U712 ( .A(n428), .Y(n645) );
  INVX1 U713 ( .A(n435), .Y(n646) );
  INVX1 U714 ( .A(n354), .Y(n647) );
  INVX1 U715 ( .A(n400), .Y(n648) );
  INVX1 U716 ( .A(n367), .Y(n649) );
  OR2X2 U717 ( .A(n808), .B(n819), .Y(n409) );
  INVX1 U718 ( .A(n409), .Y(n650) );
  INVX1 U719 ( .A(n399), .Y(n651) );
  INVX1 U720 ( .A(n370), .Y(n652) );
  INVX1 U721 ( .A(n382), .Y(n653) );
  INVX1 U722 ( .A(n393), .Y(n654) );
  INVX1 U723 ( .A(n459), .Y(n655) );
  OR2X1 U724 ( .A(n808), .B(n810), .Y(n461) );
  INVX1 U725 ( .A(n461), .Y(n656) );
  INVX1 U726 ( .A(n397), .Y(n657) );
  INVX1 U727 ( .A(n386), .Y(n658) );
  INVX1 U728 ( .A(n392), .Y(n659) );
  OR2X2 U729 ( .A(n563), .B(n566), .Y(n402) );
  INVX1 U730 ( .A(n402), .Y(n660) );
  INVX1 U731 ( .A(n356), .Y(n661) );
  INVX1 U732 ( .A(n411), .Y(n662) );
  INVX1 U733 ( .A(n381), .Y(n663) );
  INVX1 U734 ( .A(n437), .Y(n664) );
  OR2X1 U735 ( .A(n808), .B(n814), .Y(n443) );
  INVX1 U736 ( .A(n443), .Y(n665) );
  INVX1 U737 ( .A(n421), .Y(n666) );
  OR2X1 U738 ( .A(n824), .B(n809), .Y(n358) );
  INVX1 U739 ( .A(n358), .Y(n667) );
  INVX1 U740 ( .A(n404), .Y(n668) );
  OR2X1 U741 ( .A(n808), .B(n809), .Y(n463) );
  INVX1 U742 ( .A(n463), .Y(n669) );
  INVX1 U743 ( .A(n348), .Y(n670) );
  OR2X2 U744 ( .A(n823), .B(n822), .Y(n361) );
  INVX1 U745 ( .A(n361), .Y(n671) );
  OR2X2 U746 ( .A(n548), .B(n807), .Y(n455) );
  OR2X1 U747 ( .A(n824), .B(n810), .Y(n357) );
  INVX1 U748 ( .A(n357), .Y(n674) );
  INVX1 U749 ( .A(n412), .Y(n675) );
  INVX1 U750 ( .A(n403), .Y(n676) );
  INVX1 U751 ( .A(n422), .Y(n677) );
  INVX1 U752 ( .A(n359), .Y(n678) );
  INVX1 U753 ( .A(n395), .Y(n679) );
  INVX2 U754 ( .A(b[15]), .Y(n824) );
  OR2X2 U755 ( .A(n551), .B(n809), .Y(n448) );
  INVX1 U756 ( .A(n394), .Y(n682) );
  OR2X2 U757 ( .A(n822), .B(n811), .Y(n383) );
  INVX1 U758 ( .A(n383), .Y(n683) );
  INVX1 U759 ( .A(n350), .Y(n684) );
  OR2X1 U760 ( .A(n814), .B(n809), .Y(n442) );
  INVX1 U761 ( .A(n442), .Y(n685) );
  OR2X2 U762 ( .A(n553), .B(n810), .Y(n447) );
  OR2X1 U763 ( .A(n814), .B(n807), .Y(n444) );
  INVX1 U764 ( .A(n444), .Y(n690) );
  INVX1 U765 ( .A(n414), .Y(n692) );
  INVX1 U766 ( .A(n372), .Y(n693) );
  INVX1 U767 ( .A(n384), .Y(n694) );
  INVX1 U768 ( .A(n432), .Y(n695) );
  INVX1 U769 ( .A(n349), .Y(n696) );
  OR2X2 U770 ( .A(n823), .B(n820), .Y(n362) );
  INVX1 U771 ( .A(n362), .Y(n697) );
  INVX1 U772 ( .A(n351), .Y(n698) );
  INVX1 U773 ( .A(n376), .Y(n699) );
  INVX1 U774 ( .A(n364), .Y(n700) );
  INVX1 U775 ( .A(n441), .Y(n701) );
  OR2X2 U776 ( .A(n553), .B(n811), .Y(n446) );
  INVX1 U777 ( .A(n418), .Y(n704) );
  AND2X1 U778 ( .A(n182), .B(n177), .Y(n41) );
  INVX1 U779 ( .A(n41), .Y(n705) );
  AND2X1 U780 ( .A(n189), .B(n196), .Y(n49) );
  INVX1 U781 ( .A(n49), .Y(n706) );
  AND2X1 U782 ( .A(n214), .B(n205), .Y(n57) );
  INVX1 U783 ( .A(n57), .Y(n707) );
  INVX1 U784 ( .A(n431), .Y(n708) );
  INVX1 U785 ( .A(n407), .Y(n709) );
  OR2X2 U786 ( .A(n816), .B(n809), .Y(n427) );
  INVX1 U787 ( .A(n427), .Y(n710) );
  INVX1 U788 ( .A(n440), .Y(n711) );
  INVX1 U789 ( .A(n424), .Y(n712) );
  INVX1 U790 ( .A(n416), .Y(n714) );
  OR2X1 U791 ( .A(n810), .B(n809), .Y(n460) );
  INVX1 U792 ( .A(n460), .Y(n715) );
  INVX1 U793 ( .A(n451), .Y(n716) );
  OR2X1 U794 ( .A(n810), .B(n562), .Y(n434) );
  INVX1 U795 ( .A(n434), .Y(n717) );
  INVX1 U796 ( .A(n81), .Y(n718) );
  AND2X1 U797 ( .A(n236), .B(n225), .Y(n65) );
  INVX1 U798 ( .A(n65), .Y(n719) );
  INVX1 U799 ( .A(n73), .Y(n720) );
  AND2X1 U800 ( .A(n173), .B(n176), .Y(n36) );
  INVX1 U801 ( .A(n36), .Y(n721) );
  AND2X1 U802 ( .A(n197), .B(n204), .Y(n52) );
  INVX1 U803 ( .A(n52), .Y(n722) );
  AND2X2 U804 ( .A(n314), .B(n307), .Y(n99) );
  INVX1 U805 ( .A(n99), .Y(n723) );
  INVX1 U806 ( .A(n353), .Y(n724) );
  INVX1 U807 ( .A(n378), .Y(n725) );
  INVX1 U808 ( .A(n389), .Y(n726) );
  INVX1 U809 ( .A(n445), .Y(n727) );
  INVX1 U810 ( .A(n2), .Y(n729) );
  INVX1 U811 ( .A(n110), .Y(n730) );
  AND2X2 U812 ( .A(n296), .B(n575), .Y(n88) );
  INVX1 U813 ( .A(n88), .Y(n731) );
  AND2X1 U814 ( .A(n183), .B(n188), .Y(n44) );
  INVX1 U815 ( .A(n44), .Y(n732) );
  INVX1 U816 ( .A(n60), .Y(n733) );
  INVX1 U817 ( .A(n76), .Y(n734) );
  INVX1 U818 ( .A(n465), .Y(n735) );
  OR2X2 U819 ( .A(n735), .B(a[1]), .Y(n796) );
  INVX1 U820 ( .A(n363), .Y(n736) );
  OR2X2 U821 ( .A(n822), .B(n820), .Y(n375) );
  INVX1 U822 ( .A(n375), .Y(n737) );
  INVX2 U823 ( .A(b[13]), .Y(n822) );
  OR2X2 U824 ( .A(n824), .B(n566), .Y(n352) );
  INVX1 U825 ( .A(n352), .Y(n738) );
  INVX1 U826 ( .A(n365), .Y(n739) );
  INVX1 U827 ( .A(n450), .Y(n740) );
  INVX1 U828 ( .A(n369), .Y(n741) );
  INVX1 U829 ( .A(n425), .Y(n742) );
  INVX1 U830 ( .A(n417), .Y(n743) );
  INVX1 U831 ( .A(n408), .Y(n744) );
  OR2X2 U832 ( .A(n307), .B(n314), .Y(n98) );
  INVX1 U833 ( .A(n98), .Y(n745) );
  INVX1 U834 ( .A(n98), .Y(n746) );
  AND2X1 U835 ( .A(n334), .B(n329), .Y(n115) );
  INVX1 U836 ( .A(n115), .Y(n747) );
  INVX1 U837 ( .A(n68), .Y(n748) );
  OR2X1 U838 ( .A(n176), .B(n173), .Y(n35) );
  INVX1 U839 ( .A(n35), .Y(n749) );
  INVX1 U840 ( .A(n346), .Y(n750) );
  INVX1 U841 ( .A(n401), .Y(n751) );
  INVX1 U842 ( .A(n380), .Y(n752) );
  INVX1 U843 ( .A(n430), .Y(n753) );
  INVX1 U844 ( .A(n423), .Y(n754) );
  INVX1 U845 ( .A(n415), .Y(n755) );
  INVX1 U846 ( .A(n406), .Y(n756) );
  INVX1 U847 ( .A(n360), .Y(n757) );
  OR2X1 U848 ( .A(n820), .B(n810), .Y(n396) );
  INVX1 U849 ( .A(n396), .Y(n759) );
  BUFX2 U850 ( .A(n77), .Y(n760) );
  BUFX2 U851 ( .A(n53), .Y(n761) );
  INVX1 U852 ( .A(n102), .Y(n762) );
  INVX1 U853 ( .A(n3), .Y(n763) );
  INVX1 U854 ( .A(n13), .Y(n764) );
  OR2X2 U855 ( .A(n275), .B(n286), .Y(n792) );
  AND2X1 U856 ( .A(n169), .B(n172), .Y(n33) );
  INVX1 U857 ( .A(n33), .Y(n765) );
  INVX1 U858 ( .A(n93), .Y(n766) );
  OR2X1 U859 ( .A(n188), .B(n183), .Y(n43) );
  INVX1 U860 ( .A(n43), .Y(n767) );
  OR2X1 U861 ( .A(n204), .B(n197), .Y(n51) );
  INVX1 U862 ( .A(n51), .Y(n768) );
  OR2X1 U863 ( .A(n215), .B(n224), .Y(n59) );
  INVX1 U864 ( .A(n59), .Y(n769) );
  INVX1 U865 ( .A(n347), .Y(n772) );
  INVX1 U866 ( .A(n366), .Y(n773) );
  INVX1 U867 ( .A(n413), .Y(n774) );
  INVX1 U868 ( .A(n371), .Y(n775) );
  INVX1 U869 ( .A(n438), .Y(n776) );
  OR2X1 U870 ( .A(n808), .B(n820), .Y(n398) );
  INVX1 U871 ( .A(n398), .Y(n777) );
  OR2X2 U872 ( .A(n822), .B(n807), .Y(n387) );
  INVX1 U873 ( .A(n405), .Y(n779) );
  INVX1 U874 ( .A(n453), .Y(n780) );
  INVX1 U875 ( .A(n101), .Y(n781) );
  BUFX2 U876 ( .A(n82), .Y(n782) );
  INVX1 U877 ( .A(n587), .Y(n116) );
  INVX1 U878 ( .A(n731), .Y(n86) );
  OR2X1 U879 ( .A(n196), .B(n189), .Y(n783) );
  OR2X1 U880 ( .A(n249), .B(n262), .Y(n784) );
  OR2X1 U881 ( .A(n205), .B(n214), .Y(n785) );
  OR2X1 U882 ( .A(n225), .B(n236), .Y(n786) );
  INVX1 U883 ( .A(n781), .Y(n156) );
  OR2X1 U884 ( .A(n335), .B(n338), .Y(n787) );
  OR2X1 U885 ( .A(n343), .B(n344), .Y(n788) );
  OR2X1 U886 ( .A(n172), .B(n169), .Y(n791) );
  OR2X1 U887 ( .A(n177), .B(n182), .Y(n793) );
  INVX1 U888 ( .A(n632), .Y(n162) );
  XNOR2X1 U889 ( .A(n603), .B(n798), .Y(product[6]) );
  INVX1 U890 ( .A(n631), .Y(n798) );
  INVX1 U891 ( .A(b[8]), .Y(n815) );
  INVX1 U892 ( .A(n745), .Y(n155) );
  INVX1 U893 ( .A(n585), .Y(n136) );
  INVX1 U894 ( .A(n591), .Y(n94) );
  XOR2X1 U895 ( .A(n167), .B(n168), .Y(n799) );
  XOR2X1 U896 ( .A(n556), .B(n799), .Y(product[27]) );
  XOR2X1 U897 ( .A(a[4]), .B(n780), .Y(n333) );
  INVX1 U898 ( .A(n29), .Y(n139) );
  INVX1 U899 ( .A(n104), .Y(n103) );
  INVX1 U900 ( .A(n592), .Y(n804) );
  INVX1 U901 ( .A(n804), .Y(n805) );
endmodule


module alu_DW_mult_uns_26 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n26, n27, n28, n29, n33, n34, n35,
         n36, n37, n41, n42, n43, n44, n45, n49, n50, n51, n52, n53, n57, n58,
         n59, n60, n61, n65, n66, n67, n68, n69, n73, n74, n75, n76, n77, n81,
         n82, n83, n84, n87, n88, n89, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n110, n111, n115, n116, n117,
         n121, n122, n123, n124, n125, n129, n130, n131, n132, n133, n134,
         n138, n139, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n457, n458, n459, n460, n461,
         n462, n463, n465, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802;
  assign product[0] = b[0];

  FAX1 U2 ( .A(a[15]), .B(n647), .C(n26), .YC(product[31]), .YS(product[30])
         );
  FAX1 U3 ( .A(n749), .B(n164), .C(n27), .YC(n26), .YS(product[29]) );
  FAX1 U4 ( .A(n165), .B(n166), .C(n28), .YC(n27), .YS(product[28]) );
  FAX1 U5 ( .A(n167), .B(n168), .C(n139), .YC(n28), .YS(product[27]) );
  XNOR2X1 U7 ( .A(n759), .B(n724), .Y(product[26]) );
  AOI21X1 U8 ( .A(n34), .B(n765), .C(n33), .Y(n29) );
  XOR2X1 U15 ( .A(n616), .B(n697), .Y(product[25]) );
  OAI21X1 U16 ( .A(n728), .B(n617), .C(n713), .Y(n34) );
  XNOR2X1 U21 ( .A(n758), .B(n738), .Y(product[24]) );
  AOI21X1 U22 ( .A(n42), .B(n768), .C(n41), .Y(n37) );
  XOR2X1 U29 ( .A(n613), .B(n586), .Y(product[23]) );
  OAI21X1 U30 ( .A(n744), .B(n614), .C(n725), .Y(n42) );
  XNOR2X1 U35 ( .A(n549), .B(n578), .Y(product[22]) );
  AOI21X1 U36 ( .A(n50), .B(n766), .C(n49), .Y(n45) );
  XOR2X1 U43 ( .A(n611), .B(n585), .Y(product[21]) );
  OAI21X1 U44 ( .A(n554), .B(n743), .C(n714), .Y(n50) );
  XNOR2X1 U49 ( .A(n757), .B(n577), .Y(product[20]) );
  AOI21X1 U50 ( .A(n58), .B(n769), .C(n57), .Y(n53) );
  XOR2X1 U57 ( .A(n609), .B(n584), .Y(product[19]) );
  OAI21X1 U58 ( .A(n746), .B(n610), .C(n727), .Y(n58) );
  XNOR2X1 U63 ( .A(n66), .B(n576), .Y(product[18]) );
  AOI21X1 U64 ( .A(n66), .B(n761), .C(n65), .Y(n61) );
  XOR2X1 U71 ( .A(n606), .B(n583), .Y(product[17]) );
  OAI21X1 U72 ( .A(n745), .B(n607), .C(n726), .Y(n66) );
  XNOR2X1 U77 ( .A(n548), .B(n575), .Y(product[16]) );
  AOI21X1 U78 ( .A(n74), .B(n760), .C(n73), .Y(n69) );
  XOR2X1 U85 ( .A(n735), .B(n582), .Y(product[15]) );
  OAI21X1 U86 ( .A(n747), .B(n735), .C(n715), .Y(n74) );
  XNOR2X1 U91 ( .A(n550), .B(n574), .Y(product[14]) );
  AOI21X1 U92 ( .A(n82), .B(n767), .C(n81), .Y(n77) );
  XOR2X1 U99 ( .A(n567), .B(n581), .Y(product[13]) );
  OAI21X1 U100 ( .A(n556), .B(n553), .C(n552), .Y(n82) );
  AOI21X1 U102 ( .A(n87), .B(n93), .C(n88), .Y(n84) );
  XNOR2X1 U109 ( .A(n94), .B(n573), .Y(product[12]) );
  AOI21X1 U110 ( .A(n94), .B(n763), .C(n93), .Y(n89) );
  XNOR2X1 U117 ( .A(n100), .B(n686), .Y(product[11]) );
  AOI21X1 U119 ( .A(n559), .B(n104), .C(n97), .Y(n95) );
  OAI21X1 U121 ( .A(n755), .B(n722), .C(n703), .Y(n97) );
  XOR2X1 U126 ( .A(n103), .B(n580), .Y(product[10]) );
  OAI21X1 U127 ( .A(n736), .B(n103), .C(n755), .Y(n100) );
  XOR2X1 U132 ( .A(n566), .B(n579), .Y(product[9]) );
  OAI21X1 U134 ( .A(n555), .B(n562), .C(n557), .Y(n104) );
  AOI21X1 U136 ( .A(n762), .B(n115), .C(n110), .Y(n106) );
  XNOR2X1 U143 ( .A(n116), .B(n572), .Y(product[8]) );
  AOI21X1 U144 ( .A(n116), .B(n764), .C(n115), .Y(n111) );
  XNOR2X1 U151 ( .A(n122), .B(n571), .Y(product[7]) );
  AOI21X1 U153 ( .A(n122), .B(n770), .C(n121), .Y(n117) );
  XOR2X1 U160 ( .A(n569), .B(n618), .Y(product[6]) );
  OAI21X1 U161 ( .A(n598), .B(n618), .C(n595), .Y(n122) );
  XNOR2X1 U166 ( .A(n130), .B(n570), .Y(product[5]) );
  AOI21X1 U167 ( .A(n130), .B(n771), .C(n129), .Y(n125) );
  XOR2X1 U174 ( .A(n568), .B(n551), .Y(product[4]) );
  OAI21X1 U175 ( .A(n551), .B(n599), .C(n594), .Y(n130) );
  XNOR2X1 U180 ( .A(n134), .B(n138), .Y(product[3]) );
  FAX1 U190 ( .A(a[14]), .B(n604), .C(n593), .YC(n164), .YS(n165) );
  FAX1 U191 ( .A(n676), .B(n677), .C(n170), .YC(n166), .YS(n167) );
  FAX1 U192 ( .A(n657), .B(n174), .C(n171), .YC(n168), .YS(n169) );
  FAX1 U193 ( .A(a[13]), .B(n603), .C(n592), .YC(n170), .YS(n171) );
  FAX1 U194 ( .A(n180), .B(n175), .C(n178), .YC(n172), .YS(n173) );
  FAX1 U195 ( .A(n633), .B(n631), .C(n632), .YC(n174), .YS(n175) );
  FAX1 U196 ( .A(n181), .B(n184), .C(n179), .YC(n176), .YS(n177) );
  FAX1 U197 ( .A(n670), .B(n671), .C(n186), .YC(n178), .YS(n179) );
  FAX1 U198 ( .A(a[12]), .B(n601), .C(n591), .YC(n180), .YS(n181) );
  FAX1 U199 ( .A(n187), .B(n185), .C(n190), .YC(n182), .YS(n183) );
  FAX1 U200 ( .A(n750), .B(n194), .C(n192), .YC(n184), .YS(n185) );
  FAX1 U201 ( .A(n638), .B(n637), .C(n639), .YC(n186), .YS(n187) );
  FAX1 U202 ( .A(n200), .B(n191), .C(n198), .YC(n188), .YS(n189) );
  FAX1 U203 ( .A(n202), .B(n195), .C(n193), .YC(n190), .YS(n191) );
  FAX1 U204 ( .A(n628), .B(n626), .C(n627), .YC(n192), .YS(n193) );
  FAX1 U205 ( .A(a[11]), .B(n602), .C(n590), .YC(n194), .YS(n195) );
  FAX1 U206 ( .A(n208), .B(n199), .C(n206), .YC(n196), .YS(n197) );
  FAX1 U207 ( .A(n210), .B(n203), .C(n201), .YC(n198), .YS(n199) );
  FAX1 U208 ( .A(n652), .B(n653), .C(n212), .YC(n200), .YS(n201) );
  FAX1 U209 ( .A(n621), .B(n619), .C(n620), .YC(n202), .YS(n203) );
  FAX1 U210 ( .A(n209), .B(n216), .C(n207), .YC(n204), .YS(n205) );
  FAX1 U211 ( .A(n213), .B(n211), .C(n218), .YC(n206), .YS(n207) );
  FAX1 U212 ( .A(n729), .B(n222), .C(n220), .YC(n208), .YS(n209) );
  FAX1 U213 ( .A(n646), .B(n644), .C(n645), .YC(n210), .YS(n211) );
  FAX1 U214 ( .A(a[10]), .B(n643), .C(n642), .YC(n212), .YS(n213) );
  FAX1 U215 ( .A(n219), .B(n226), .C(n217), .YC(n214), .YS(n215) );
  FAX1 U216 ( .A(n223), .B(n230), .C(n228), .YC(n216), .YS(n217) );
  FAX1 U217 ( .A(n234), .B(n232), .C(n221), .YC(n218), .YS(n219) );
  FAX1 U218 ( .A(n658), .B(n659), .C(n660), .YC(n220), .YS(n221) );
  FAX1 U219 ( .A(n667), .B(n665), .C(n666), .YC(n222), .YS(n223) );
  FAX1 U220 ( .A(n229), .B(n238), .C(n227), .YC(n224), .YS(n225) );
  FAX1 U221 ( .A(n242), .B(n231), .C(n240), .YC(n226), .YS(n227) );
  FAX1 U222 ( .A(n244), .B(n235), .C(n233), .YC(n228), .YS(n229) );
  FAX1 U223 ( .A(n719), .B(n718), .C(n246), .YC(n230), .YS(n231) );
  FAX1 U224 ( .A(n707), .B(n705), .C(n706), .YC(n232), .YS(n233) );
  FAX1 U225 ( .A(a[9]), .B(n625), .C(n624), .YC(n234), .YS(n235) );
  FAX1 U226 ( .A(n241), .B(n250), .C(n239), .YC(n236), .YS(n237) );
  FAX1 U227 ( .A(n254), .B(n243), .C(n252), .YC(n238), .YS(n239) );
  FAX1 U228 ( .A(n256), .B(n247), .C(n245), .YC(n240), .YS(n241) );
  FAX1 U229 ( .A(n751), .B(n260), .C(n258), .YC(n242), .YS(n243) );
  FAX1 U230 ( .A(n682), .B(n684), .C(n683), .YC(n244), .YS(n245) );
  FAX1 U231 ( .A(n662), .B(n664), .C(n663), .YC(n246), .YS(n247) );
  FAX1 U232 ( .A(n253), .B(n264), .C(n251), .YC(n248), .YS(n249) );
  FAX1 U233 ( .A(n268), .B(n255), .C(n266), .YC(n250), .YS(n251) );
  FAX1 U234 ( .A(n270), .B(n259), .C(n257), .YC(n252), .YS(n253) );
  FAX1 U235 ( .A(n721), .B(n272), .C(n261), .YC(n254), .YS(n255) );
  FAX1 U236 ( .A(n688), .B(n690), .C(n689), .YC(n256), .YS(n257) );
  FAX1 U237 ( .A(n692), .B(n693), .C(n694), .YC(n258), .YS(n259) );
  HAX1 U238 ( .A(a[8]), .B(n696), .YC(n260), .YS(n261) );
  FAX1 U239 ( .A(n267), .B(n276), .C(n265), .YC(n262), .YS(n263) );
  FAX1 U240 ( .A(n271), .B(n269), .C(n278), .YC(n264), .YS(n265) );
  FAX1 U241 ( .A(n273), .B(n282), .C(n280), .YC(n266), .YS(n267) );
  FAX1 U242 ( .A(n733), .B(n734), .C(n284), .YC(n268), .YS(n269) );
  FAX1 U243 ( .A(n710), .B(n709), .C(n708), .YC(n270), .YS(n271) );
  HAX1 U244 ( .A(n668), .B(n669), .YC(n272), .YS(n273) );
  FAX1 U245 ( .A(n279), .B(n288), .C(n277), .YC(n274), .YS(n275) );
  FAX1 U246 ( .A(n283), .B(n281), .C(n290), .YC(n276), .YS(n277) );
  FAX1 U247 ( .A(n294), .B(n285), .C(n292), .YC(n278), .YS(n279) );
  FAX1 U248 ( .A(n731), .B(n730), .C(n732), .YC(n280), .YS(n281) );
  FAX1 U249 ( .A(n754), .B(n753), .C(n752), .YC(n282), .YS(n283) );
  HAX1 U250 ( .A(a[7]), .B(n685), .YC(n284), .YS(n285) );
  FAX1 U251 ( .A(n291), .B(n298), .C(n289), .YC(n286), .YS(n287) );
  FAX1 U252 ( .A(n774), .B(n293), .C(n300), .YC(n288), .YS(n289) );
  FAX1 U253 ( .A(n720), .B(n304), .C(n295), .YC(n290), .YS(n291) );
  FAX1 U254 ( .A(n785), .B(n600), .C(n589), .YC(n292), .YS(n293) );
  HAX1 U255 ( .A(n636), .B(n635), .YC(n294), .YS(n295) );
  FAX1 U257 ( .A(n305), .B(n310), .C(n303), .YC(n298), .YS(n299) );
  FAX1 U258 ( .A(n679), .B(n678), .C(n312), .YC(n300), .YS(n301) );
  HAX1 U260 ( .A(a[6]), .B(n675), .YC(n304), .YS(n305) );
  FAX1 U261 ( .A(n311), .B(n316), .C(n309), .YC(n306), .YS(n307) );
  FAX1 U262 ( .A(n313), .B(n320), .C(n318), .YC(n308), .YS(n309) );
  FAX1 U263 ( .A(n674), .B(n673), .C(n672), .YC(n310), .YS(n311) );
  HAX1 U264 ( .A(n622), .B(n623), .YC(n312), .YS(n313) );
  FAX1 U265 ( .A(n319), .B(n324), .C(n317), .YC(n314), .YS(n315) );
  FAX1 U266 ( .A(n691), .B(n326), .C(n321), .YC(n316), .YS(n317) );
  FAX1 U267 ( .A(n680), .B(n442), .C(n681), .YC(n318), .YS(n319) );
  HAX1 U268 ( .A(a[5]), .B(n634), .YC(n320), .YS(n321) );
  FAX1 U269 ( .A(n327), .B(n330), .C(n325), .YC(n322), .YS(n323) );
  FAX1 U270 ( .A(n651), .B(n650), .C(n332), .YC(n324), .YS(n325) );
  HAX1 U271 ( .A(n630), .B(n629), .YC(n326), .YS(n327) );
  FAX1 U272 ( .A(n336), .B(n333), .C(n331), .YC(n328), .YS(n329) );
  FAX1 U273 ( .A(n777), .B(n656), .C(n655), .YC(n330), .YS(n331) );
  HAX1 U274 ( .A(a[4]), .B(n641), .YC(n332), .YS(n333) );
  FAX1 U275 ( .A(n717), .B(n340), .C(n337), .YC(n334), .YS(n335) );
  HAX1 U276 ( .A(n565), .B(n564), .YC(n336), .YS(n337) );
  FAX1 U277 ( .A(n648), .B(n649), .C(n342), .YC(n338), .YS(n339) );
  HAX1 U278 ( .A(a[3]), .B(n654), .YC(n340), .YS(n341) );
  HAX1 U279 ( .A(n459), .B(n640), .YC(n342), .YS(n343) );
  HAX1 U280 ( .A(a[2]), .B(n462), .YC(n344), .YS(n345) );
  INVX8 U434 ( .A(b[2]), .Y(n788) );
  OR2X1 U435 ( .A(n793), .B(n789), .Y(n441) );
  OR2X1 U436 ( .A(n787), .B(n786), .Y(n465) );
  OR2X1 U437 ( .A(n797), .B(n796), .Y(n400) );
  OR2X1 U438 ( .A(n795), .B(n796), .Y(n411) );
  OR2X1 U439 ( .A(n802), .B(n789), .Y(n357) );
  OR2X1 U440 ( .A(n793), .B(n797), .Y(n403) );
  OR2X1 U441 ( .A(n796), .B(n794), .Y(n412) );
  OR2X1 U442 ( .A(n792), .B(n797), .Y(n404) );
  OR2X1 U443 ( .A(n800), .B(n789), .Y(n384) );
  OR2X1 U444 ( .A(n792), .B(n796), .Y(n414) );
  OR2X1 U445 ( .A(n797), .B(n790), .Y(n406) );
  OR2X1 U446 ( .A(n796), .B(n791), .Y(n415) );
  OR2X1 U447 ( .A(n796), .B(n790), .Y(n416) );
  OR2X1 U448 ( .A(n797), .B(n789), .Y(n407) );
  OR2X1 U449 ( .A(n796), .B(n789), .Y(n417) );
  OR2X1 U450 ( .A(n797), .B(n788), .Y(n408) );
  OR2X1 U451 ( .A(n793), .B(n796), .Y(n413) );
  INVX1 U452 ( .A(n385), .Y(n692) );
  OR2X1 U453 ( .A(n787), .B(n796), .Y(n419) );
  OR2X1 U454 ( .A(n797), .B(n786), .Y(n410) );
  OR2X1 U455 ( .A(n787), .B(n795), .Y(n428) );
  OR2X1 U456 ( .A(n801), .B(n796), .Y(n364) );
  OR2X1 U457 ( .A(n801), .B(n797), .Y(n363) );
  OR2X1 U458 ( .A(n800), .B(n796), .Y(n377) );
  OR2X1 U459 ( .A(n795), .B(n797), .Y(n401) );
  OR2X1 U460 ( .A(n796), .B(n788), .Y(n418) );
  INVX1 U461 ( .A(n441), .Y(n672) );
  INVX1 U462 ( .A(n446), .Y(n673) );
  AND2X1 U463 ( .A(b[7]), .B(b[2]), .Y(n442) );
  INVX1 U464 ( .A(n452), .Y(n651) );
  OR2X1 U465 ( .A(n787), .B(n788), .Y(n463) );
  INVX1 U466 ( .A(b[13]), .Y(n800) );
  OR2X1 U467 ( .A(n802), .B(n796), .Y(n350) );
  OR2X1 U468 ( .A(n802), .B(n797), .Y(n349) );
  AND2X1 U469 ( .A(n698), .B(n768), .Y(n3) );
  AND2X1 U470 ( .A(n687), .B(n87), .Y(n14) );
  AND2X1 U471 ( .A(n587), .B(n138), .Y(n133) );
  AND2X1 U472 ( .A(n661), .B(n773), .Y(product[2]) );
  OR2X1 U473 ( .A(n597), .B(n287), .Y(n87) );
  INVX2 U474 ( .A(b[10]), .Y(n796) );
  INVX1 U475 ( .A(b[0]), .Y(n786) );
  INVX2 U476 ( .A(b[9]), .Y(n795) );
  INVX1 U477 ( .A(b[7]), .Y(n793) );
  INVX2 U478 ( .A(b[6]), .Y(n792) );
  INVX2 U479 ( .A(b[11]), .Y(n797) );
  AND2X1 U480 ( .A(n597), .B(n287), .Y(n88) );
  INVX1 U481 ( .A(b[1]), .Y(n787) );
  INVX1 U482 ( .A(b[3]), .Y(n789) );
  INVX1 U483 ( .A(b[4]), .Y(n790) );
  AND2X1 U484 ( .A(b[3]), .B(b[4]), .Y(n777) );
  INVX1 U485 ( .A(b[5]), .Y(n791) );
  BUFX2 U486 ( .A(n299), .Y(n547) );
  OAI21X1 U487 ( .A(n747), .B(n735), .C(n715), .Y(n548) );
  OAI21X1 U488 ( .A(n554), .B(n743), .C(n714), .Y(n549) );
  BUFX2 U489 ( .A(n82), .Y(n550) );
  OR2X2 U490 ( .A(n797), .B(n798), .Y(n388) );
  OR2X2 U491 ( .A(n797), .B(n794), .Y(n402) );
  OR2X2 U492 ( .A(n797), .B(n791), .Y(n405) );
  XNOR2X1 U493 ( .A(n410), .B(n419), .Y(n775) );
  INVX1 U494 ( .A(n419), .Y(n737) );
  OR2X1 U495 ( .A(n787), .B(n789), .Y(n461) );
  INVX8 U496 ( .A(b[8]), .Y(n794) );
  AND2X2 U497 ( .A(a[1]), .B(n716), .Y(n138) );
  AND2X2 U498 ( .A(n308), .B(n299), .Y(n779) );
  OR2X2 U499 ( .A(n787), .B(n797), .Y(n409) );
  INVX1 U500 ( .A(n133), .Y(n551) );
  BUFX2 U501 ( .A(n84), .Y(n552) );
  AND2X2 U502 ( .A(n763), .B(n87), .Y(n83) );
  INVX1 U503 ( .A(n83), .Y(n553) );
  BUFX2 U504 ( .A(n53), .Y(n554) );
  BUFX2 U505 ( .A(n117), .Y(n555) );
  BUFX2 U506 ( .A(n95), .Y(n556) );
  AND2X1 U507 ( .A(b[4]), .B(b[8]), .Y(n785) );
  BUFX2 U508 ( .A(n106), .Y(n557) );
  AND2X1 U509 ( .A(n756), .B(n723), .Y(n782) );
  INVX1 U510 ( .A(n782), .Y(n558) );
  OR2X1 U511 ( .A(n722), .B(n736), .Y(n96) );
  INVX1 U512 ( .A(n96), .Y(n559) );
  AND2X2 U513 ( .A(n301), .B(n299), .Y(n780) );
  INVX1 U514 ( .A(n780), .Y(n560) );
  AND2X1 U515 ( .A(n737), .B(n723), .Y(n783) );
  INVX1 U516 ( .A(n783), .Y(n561) );
  AND2X1 U517 ( .A(n764), .B(n762), .Y(n105) );
  INVX1 U518 ( .A(n105), .Y(n562) );
  AND2X1 U519 ( .A(n737), .B(n756), .Y(n784) );
  INVX1 U520 ( .A(n784), .Y(n563) );
  OR2X1 U521 ( .A(n787), .B(n791), .Y(n454) );
  INVX1 U522 ( .A(n454), .Y(n564) );
  OR2X1 U523 ( .A(n790), .B(n788), .Y(n457) );
  INVX1 U524 ( .A(n457), .Y(n565) );
  BUFX2 U525 ( .A(n111), .Y(n566) );
  BUFX2 U526 ( .A(n89), .Y(n567) );
  AND2X1 U527 ( .A(n594), .B(n131), .Y(n23) );
  INVX1 U528 ( .A(n23), .Y(n568) );
  AND2X1 U529 ( .A(n595), .B(n123), .Y(n21) );
  INVX1 U530 ( .A(n21), .Y(n569) );
  AND2X1 U531 ( .A(n740), .B(n771), .Y(n22) );
  INVX1 U532 ( .A(n22), .Y(n570) );
  AND2X1 U533 ( .A(n588), .B(n770), .Y(n20) );
  INVX1 U534 ( .A(n20), .Y(n571) );
  AND2X1 U535 ( .A(n741), .B(n764), .Y(n19) );
  INVX1 U536 ( .A(n19), .Y(n572) );
  AND2X1 U537 ( .A(n742), .B(n763), .Y(n15) );
  INVX1 U538 ( .A(n15), .Y(n573) );
  AND2X1 U539 ( .A(n701), .B(n767), .Y(n13) );
  INVX1 U540 ( .A(n13), .Y(n574) );
  AND2X1 U541 ( .A(n702), .B(n760), .Y(n11) );
  INVX1 U542 ( .A(n11), .Y(n575) );
  AND2X1 U543 ( .A(n712), .B(n761), .Y(n9) );
  INVX1 U544 ( .A(n9), .Y(n576) );
  AND2X1 U545 ( .A(n700), .B(n769), .Y(n7) );
  INVX1 U546 ( .A(n7), .Y(n577) );
  AND2X1 U547 ( .A(n699), .B(n766), .Y(n5) );
  INVX1 U548 ( .A(n5), .Y(n578) );
  AND2X1 U549 ( .A(n711), .B(n762), .Y(n18) );
  INVX1 U550 ( .A(n18), .Y(n579) );
  AND2X1 U551 ( .A(n755), .B(n101), .Y(n17) );
  INVX1 U552 ( .A(n17), .Y(n580) );
  INVX1 U553 ( .A(n14), .Y(n581) );
  AND2X1 U554 ( .A(n715), .B(n75), .Y(n12) );
  INVX1 U555 ( .A(n12), .Y(n582) );
  AND2X1 U556 ( .A(n726), .B(n67), .Y(n10) );
  INVX1 U557 ( .A(n10), .Y(n583) );
  AND2X1 U558 ( .A(n727), .B(n59), .Y(n8) );
  INVX1 U559 ( .A(n8), .Y(n584) );
  AND2X1 U560 ( .A(n714), .B(n51), .Y(n6) );
  INVX1 U561 ( .A(n6), .Y(n585) );
  AND2X1 U562 ( .A(n725), .B(n43), .Y(n4) );
  INVX1 U563 ( .A(n4), .Y(n586) );
  OR2X1 U564 ( .A(n788), .B(n786), .Y(n134) );
  INVX1 U565 ( .A(n134), .Y(n587) );
  AND2X1 U566 ( .A(n338), .B(n335), .Y(n121) );
  INVX1 U567 ( .A(n121), .Y(n588) );
  OR2X1 U568 ( .A(n793), .B(n791), .Y(n439) );
  INVX1 U569 ( .A(n439), .Y(n589) );
  OR2X1 U570 ( .A(n795), .B(n798), .Y(n390) );
  INVX1 U571 ( .A(n390), .Y(n590) );
  INVX1 U572 ( .A(n377), .Y(n591) );
  INVX1 U573 ( .A(n363), .Y(n592) );
  OR2X1 U574 ( .A(n802), .B(n798), .Y(n348) );
  INVX1 U575 ( .A(n348), .Y(n593) );
  AND2X1 U576 ( .A(n704), .B(n345), .Y(n132) );
  INVX1 U577 ( .A(n132), .Y(n594) );
  AND2X1 U578 ( .A(n341), .B(n339), .Y(n124) );
  INVX1 U579 ( .A(n124), .Y(n595) );
  INVX1 U580 ( .A(n776), .Y(n596) );
  INVX1 U581 ( .A(n596), .Y(n597) );
  OR2X1 U582 ( .A(n339), .B(n341), .Y(n123) );
  INVX1 U583 ( .A(n123), .Y(n598) );
  OR2X1 U584 ( .A(n345), .B(n704), .Y(n131) );
  INVX1 U585 ( .A(n131), .Y(n599) );
  OR2X1 U586 ( .A(n795), .B(n789), .Y(n426) );
  INVX1 U587 ( .A(n426), .Y(n600) );
  INVX1 U588 ( .A(n388), .Y(n601) );
  OR2X1 U589 ( .A(n800), .B(n794), .Y(n379) );
  INVX1 U590 ( .A(n379), .Y(n602) );
  OR2X1 U591 ( .A(n800), .B(n798), .Y(n375) );
  INVX1 U592 ( .A(n375), .Y(n603) );
  OR2X1 U593 ( .A(n801), .B(n800), .Y(n361) );
  INVX1 U594 ( .A(n361), .Y(n604) );
  INVX1 U595 ( .A(n69), .Y(n605) );
  INVX1 U596 ( .A(n605), .Y(n606) );
  INVX1 U597 ( .A(n605), .Y(n607) );
  INVX1 U598 ( .A(n61), .Y(n608) );
  INVX1 U599 ( .A(n608), .Y(n609) );
  INVX1 U600 ( .A(n608), .Y(n610) );
  BUFX2 U601 ( .A(n554), .Y(n611) );
  INVX1 U602 ( .A(n45), .Y(n612) );
  INVX1 U603 ( .A(n612), .Y(n613) );
  INVX1 U604 ( .A(n612), .Y(n614) );
  INVX1 U605 ( .A(n37), .Y(n615) );
  INVX1 U606 ( .A(n615), .Y(n616) );
  INVX1 U607 ( .A(n615), .Y(n617) );
  BUFX2 U608 ( .A(n125), .Y(n618) );
  OR2X1 U609 ( .A(n801), .B(n792), .Y(n368) );
  INVX1 U610 ( .A(n368), .Y(n619) );
  OR2X1 U611 ( .A(n802), .B(n791), .Y(n355) );
  INVX1 U612 ( .A(n355), .Y(n620) );
  OR2X1 U613 ( .A(n798), .B(n794), .Y(n391) );
  INVX1 U614 ( .A(n391), .Y(n621) );
  OR2X1 U615 ( .A(n794), .B(n788), .Y(n435) );
  INVX1 U616 ( .A(n435), .Y(n622) );
  INVX1 U617 ( .A(n428), .Y(n623) );
  OR2X1 U618 ( .A(n791), .B(n798), .Y(n394) );
  INVX1 U619 ( .A(n394), .Y(n624) );
  OR2X1 U620 ( .A(n800), .B(n790), .Y(n383) );
  INVX1 U621 ( .A(n383), .Y(n625) );
  OR2X1 U622 ( .A(n801), .B(n793), .Y(n367) );
  INVX1 U623 ( .A(n367), .Y(n626) );
  OR2X1 U624 ( .A(n802), .B(n792), .Y(n354) );
  INVX1 U625 ( .A(n354), .Y(n627) );
  INVX1 U626 ( .A(n400), .Y(n628) );
  OR2X1 U627 ( .A(n787), .B(n793), .Y(n443) );
  INVX1 U628 ( .A(n443), .Y(n629) );
  OR2X1 U629 ( .A(n794), .B(n786), .Y(n437) );
  INVX1 U630 ( .A(n437), .Y(n630) );
  OR2X1 U631 ( .A(n797), .B(n800), .Y(n376) );
  INVX1 U632 ( .A(n376), .Y(n631) );
  OR2X1 U633 ( .A(n802), .B(n795), .Y(n351) );
  INVX1 U634 ( .A(n351), .Y(n632) );
  INVX1 U635 ( .A(n364), .Y(n633) );
  OR2X1 U636 ( .A(n791), .B(n790), .Y(n451) );
  INVX1 U637 ( .A(n451), .Y(n634) );
  INVX1 U638 ( .A(n409), .Y(n635) );
  OR2X1 U639 ( .A(n799), .B(n786), .Y(n399) );
  INVX1 U640 ( .A(n399), .Y(n636) );
  OR2X1 U641 ( .A(n795), .B(n800), .Y(n378) );
  INVX1 U642 ( .A(n378), .Y(n637) );
  OR2X1 U643 ( .A(n796), .B(n798), .Y(n389) );
  INVX1 U644 ( .A(n389), .Y(n638) );
  OR2X1 U645 ( .A(n802), .B(n793), .Y(n353) );
  INVX1 U646 ( .A(n353), .Y(n639) );
  INVX1 U647 ( .A(n461), .Y(n640) );
  OR2X1 U648 ( .A(n791), .B(n788), .Y(n453) );
  INVX1 U649 ( .A(n453), .Y(n641) );
  OR2X1 U650 ( .A(n793), .B(n798), .Y(n392) );
  INVX1 U651 ( .A(n392), .Y(n642) );
  INVX1 U652 ( .A(n402), .Y(n643) );
  OR2X1 U653 ( .A(n792), .B(n800), .Y(n381) );
  INVX1 U654 ( .A(n381), .Y(n644) );
  OR2X1 U655 ( .A(n802), .B(n790), .Y(n356) );
  INVX1 U656 ( .A(n356), .Y(n645) );
  INVX1 U657 ( .A(n411), .Y(n646) );
  OR2X1 U658 ( .A(n802), .B(n801), .Y(n346) );
  INVX1 U659 ( .A(n346), .Y(n647) );
  OR2X1 U660 ( .A(n791), .B(n786), .Y(n455) );
  INVX1 U661 ( .A(n455), .Y(n648) );
  OR2X1 U662 ( .A(n787), .B(n790), .Y(n458) );
  INVX1 U663 ( .A(n458), .Y(n649) );
  OR2X1 U664 ( .A(n792), .B(n788), .Y(n448) );
  INVX1 U665 ( .A(n448), .Y(n650) );
  OR2X1 U666 ( .A(n791), .B(n789), .Y(n452) );
  OR2X1 U667 ( .A(n793), .B(n800), .Y(n380) );
  INVX1 U668 ( .A(n380), .Y(n652) );
  INVX1 U669 ( .A(n401), .Y(n653) );
  OR2X1 U670 ( .A(n789), .B(n788), .Y(n460) );
  INVX1 U671 ( .A(n460), .Y(n654) );
  OR2X1 U672 ( .A(n787), .B(n792), .Y(n449) );
  INVX1 U673 ( .A(n449), .Y(n655) );
  OR2X1 U674 ( .A(n793), .B(n786), .Y(n444) );
  INVX1 U675 ( .A(n444), .Y(n656) );
  INVX1 U676 ( .A(n350), .Y(n657) );
  OR2X1 U677 ( .A(n792), .B(n798), .Y(n393) );
  INVX1 U678 ( .A(n393), .Y(n658) );
  OR2X1 U679 ( .A(n800), .B(n791), .Y(n382) );
  INVX1 U680 ( .A(n382), .Y(n659) );
  OR2X1 U681 ( .A(n801), .B(n790), .Y(n370) );
  INVX1 U682 ( .A(n370), .Y(n660) );
  INVX1 U683 ( .A(n138), .Y(n661) );
  OR2X1 U684 ( .A(n798), .B(n790), .Y(n395) );
  INVX1 U685 ( .A(n395), .Y(n662) );
  OR2X1 U686 ( .A(n802), .B(n787), .Y(n359) );
  INVX1 U687 ( .A(n359), .Y(n663) );
  OR2X1 U688 ( .A(n793), .B(n795), .Y(n422) );
  INVX1 U689 ( .A(n422), .Y(n664) );
  INVX1 U690 ( .A(n403), .Y(n665) );
  INVX1 U691 ( .A(n357), .Y(n666) );
  INVX1 U692 ( .A(n412), .Y(n667) );
  OR2X1 U693 ( .A(n799), .B(n788), .Y(n397) );
  INVX1 U694 ( .A(n397), .Y(n668) );
  OR2X1 U695 ( .A(n787), .B(n800), .Y(n386) );
  INVX1 U696 ( .A(n386), .Y(n669) );
  OR2X1 U697 ( .A(n801), .B(n795), .Y(n365) );
  INVX1 U698 ( .A(n365), .Y(n670) );
  OR2X1 U699 ( .A(n802), .B(n794), .Y(n352) );
  INVX1 U700 ( .A(n352), .Y(n671) );
  OR2X1 U701 ( .A(n792), .B(n790), .Y(n446) );
  OR2X1 U702 ( .A(n796), .B(n786), .Y(n420) );
  INVX1 U703 ( .A(n420), .Y(n674) );
  OR2X2 U704 ( .A(n789), .B(n794), .Y(n434) );
  INVX1 U705 ( .A(n434), .Y(n675) );
  OR2X1 U706 ( .A(n801), .B(n798), .Y(n362) );
  INVX1 U707 ( .A(n362), .Y(n676) );
  INVX1 U708 ( .A(n349), .Y(n677) );
  OR2X1 U709 ( .A(n793), .B(n790), .Y(n440) );
  INVX1 U710 ( .A(n440), .Y(n678) );
  OR2X1 U711 ( .A(n795), .B(n788), .Y(n427) );
  INVX1 U712 ( .A(n427), .Y(n679) );
  OR2X1 U713 ( .A(n795), .B(n786), .Y(n429) );
  INVX1 U714 ( .A(n429), .Y(n680) );
  OR2X1 U715 ( .A(n787), .B(n794), .Y(n436) );
  INVX1 U716 ( .A(n436), .Y(n681) );
  INVX1 U717 ( .A(n384), .Y(n682) );
  OR2X1 U718 ( .A(n801), .B(n788), .Y(n372) );
  INVX1 U719 ( .A(n372), .Y(n683) );
  INVX1 U720 ( .A(n414), .Y(n684) );
  OR2X1 U721 ( .A(n791), .B(n794), .Y(n432) );
  INVX1 U722 ( .A(n432), .Y(n685) );
  AND2X1 U723 ( .A(n703), .B(n98), .Y(n16) );
  INVX1 U724 ( .A(n16), .Y(n686) );
  INVX1 U725 ( .A(n88), .Y(n687) );
  INVX1 U726 ( .A(n406), .Y(n688) );
  OR2X1 U727 ( .A(n792), .B(n795), .Y(n423) );
  INVX1 U728 ( .A(n423), .Y(n689) );
  INVX1 U729 ( .A(n415), .Y(n690) );
  OR2X1 U730 ( .A(n792), .B(n789), .Y(n447) );
  INVX1 U731 ( .A(n447), .Y(n691) );
  OR2X1 U732 ( .A(n800), .B(n788), .Y(n385) );
  OR2X1 U733 ( .A(n787), .B(n801), .Y(n373) );
  INVX1 U734 ( .A(n373), .Y(n693) );
  OR2X1 U735 ( .A(n802), .B(n786), .Y(n360) );
  INVX1 U736 ( .A(n360), .Y(n694) );
  INVX1 U737 ( .A(n779), .Y(n695) );
  OR2X1 U738 ( .A(n798), .B(n789), .Y(n396) );
  INVX1 U739 ( .A(n396), .Y(n696) );
  AND2X1 U740 ( .A(n713), .B(n35), .Y(n2) );
  INVX1 U741 ( .A(n2), .Y(n697) );
  AND2X1 U742 ( .A(n182), .B(n177), .Y(n41) );
  INVX1 U743 ( .A(n41), .Y(n698) );
  AND2X1 U744 ( .A(n189), .B(n196), .Y(n49) );
  INVX1 U745 ( .A(n49), .Y(n699) );
  AND2X1 U746 ( .A(n214), .B(n205), .Y(n57) );
  INVX1 U747 ( .A(n57), .Y(n700) );
  AND2X1 U748 ( .A(n286), .B(n275), .Y(n81) );
  INVX1 U749 ( .A(n81), .Y(n701) );
  AND2X1 U750 ( .A(n262), .B(n249), .Y(n73) );
  INVX1 U751 ( .A(n73), .Y(n702) );
  AND2X1 U752 ( .A(n314), .B(n307), .Y(n99) );
  INVX1 U753 ( .A(n99), .Y(n703) );
  INVX1 U754 ( .A(n463), .Y(n704) );
  INVX1 U755 ( .A(n404), .Y(n705) );
  OR2X1 U756 ( .A(n802), .B(n788), .Y(n358) );
  INVX1 U757 ( .A(n358), .Y(n706) );
  OR2X1 U758 ( .A(n795), .B(n794), .Y(n421) );
  INVX1 U759 ( .A(n421), .Y(n707) );
  OR2X1 U760 ( .A(n801), .B(n786), .Y(n374) );
  INVX1 U761 ( .A(n374), .Y(n708) );
  OR2X1 U762 ( .A(n795), .B(n791), .Y(n424) );
  INVX1 U763 ( .A(n424), .Y(n709) );
  INVX1 U764 ( .A(n416), .Y(n710) );
  AND2X1 U765 ( .A(n328), .B(n323), .Y(n110) );
  INVX1 U766 ( .A(n110), .Y(n711) );
  AND2X1 U767 ( .A(n236), .B(n225), .Y(n65) );
  INVX1 U768 ( .A(n65), .Y(n712) );
  AND2X1 U769 ( .A(n173), .B(n176), .Y(n36) );
  INVX1 U770 ( .A(n36), .Y(n713) );
  AND2X1 U771 ( .A(n197), .B(n204), .Y(n52) );
  INVX1 U772 ( .A(n52), .Y(n714) );
  AND2X1 U773 ( .A(n274), .B(n263), .Y(n76) );
  INVX1 U774 ( .A(n76), .Y(n715) );
  INVX1 U775 ( .A(n465), .Y(n716) );
  OR2X2 U776 ( .A(n716), .B(a[1]), .Y(n773) );
  OR2X1 U777 ( .A(n792), .B(n786), .Y(n450) );
  INVX1 U778 ( .A(n450), .Y(n717) );
  OR2X1 U779 ( .A(n801), .B(n789), .Y(n371) );
  INVX1 U780 ( .A(n371), .Y(n718) );
  INVX1 U781 ( .A(n413), .Y(n719) );
  INVX1 U782 ( .A(n418), .Y(n720) );
  OR2X1 U783 ( .A(n793), .B(n794), .Y(n430) );
  INVX1 U784 ( .A(n430), .Y(n721) );
  OR2X1 U785 ( .A(n307), .B(n314), .Y(n98) );
  INVX1 U786 ( .A(n98), .Y(n722) );
  OR2X1 U787 ( .A(n792), .B(n791), .Y(n445) );
  INVX1 U788 ( .A(n445), .Y(n723) );
  AND2X1 U789 ( .A(n739), .B(n765), .Y(n1) );
  INVX1 U790 ( .A(n1), .Y(n724) );
  AND2X1 U791 ( .A(n183), .B(n188), .Y(n44) );
  INVX1 U792 ( .A(n44), .Y(n725) );
  AND2X1 U793 ( .A(n248), .B(n237), .Y(n68) );
  INVX1 U794 ( .A(n68), .Y(n726) );
  AND2X1 U795 ( .A(n224), .B(n215), .Y(n60) );
  INVX1 U796 ( .A(n60), .Y(n727) );
  OR2X1 U797 ( .A(n176), .B(n173), .Y(n35) );
  INVX1 U798 ( .A(n35), .Y(n728) );
  OR2X1 U799 ( .A(n801), .B(n791), .Y(n369) );
  INVX1 U800 ( .A(n369), .Y(n729) );
  INVX1 U801 ( .A(n408), .Y(n730) );
  OR2X1 U802 ( .A(n800), .B(n786), .Y(n387) );
  INVX1 U803 ( .A(n387), .Y(n731) );
  OR2X1 U804 ( .A(n795), .B(n790), .Y(n425) );
  INVX1 U805 ( .A(n425), .Y(n732) );
  INVX1 U806 ( .A(n407), .Y(n733) );
  OR2X1 U807 ( .A(n792), .B(n794), .Y(n431) );
  INVX1 U808 ( .A(n431), .Y(n734) );
  BUFX2 U809 ( .A(n77), .Y(n735) );
  OR2X1 U810 ( .A(n315), .B(n322), .Y(n101) );
  INVX1 U811 ( .A(n101), .Y(n736) );
  INVX1 U812 ( .A(n3), .Y(n738) );
  AND2X1 U813 ( .A(n169), .B(n172), .Y(n33) );
  INVX1 U814 ( .A(n33), .Y(n739) );
  AND2X1 U815 ( .A(n344), .B(n343), .Y(n129) );
  INVX1 U816 ( .A(n129), .Y(n740) );
  AND2X1 U817 ( .A(n334), .B(n329), .Y(n115) );
  INVX1 U818 ( .A(n115), .Y(n741) );
  AND2X1 U819 ( .A(n306), .B(n297), .Y(n93) );
  INVX1 U820 ( .A(n93), .Y(n742) );
  OR2X1 U821 ( .A(n204), .B(n197), .Y(n51) );
  INVX1 U822 ( .A(n51), .Y(n743) );
  OR2X1 U823 ( .A(n188), .B(n183), .Y(n43) );
  INVX1 U824 ( .A(n43), .Y(n744) );
  OR2X1 U825 ( .A(n237), .B(n248), .Y(n67) );
  INVX1 U826 ( .A(n67), .Y(n745) );
  OR2X1 U827 ( .A(n215), .B(n224), .Y(n59) );
  INVX1 U828 ( .A(n59), .Y(n746) );
  OR2X1 U829 ( .A(n263), .B(n274), .Y(n75) );
  INVX1 U830 ( .A(n75), .Y(n747) );
  AND2X1 U831 ( .A(n301), .B(n308), .Y(n781) );
  INVX1 U832 ( .A(n781), .Y(n748) );
  OR2X1 U833 ( .A(n802), .B(n800), .Y(n347) );
  INVX1 U834 ( .A(n347), .Y(n749) );
  OR2X1 U835 ( .A(n801), .B(n794), .Y(n366) );
  INVX1 U836 ( .A(n366), .Y(n750) );
  INVX1 U837 ( .A(n405), .Y(n751) );
  OR2X1 U838 ( .A(n793), .B(n792), .Y(n438) );
  INVX1 U839 ( .A(n438), .Y(n752) );
  OR2X1 U840 ( .A(n787), .B(n798), .Y(n398) );
  INVX1 U841 ( .A(n398), .Y(n753) );
  INVX1 U842 ( .A(n417), .Y(n754) );
  AND2X1 U843 ( .A(n322), .B(n315), .Y(n102) );
  INVX1 U844 ( .A(n102), .Y(n755) );
  INVX1 U845 ( .A(n410), .Y(n756) );
  BUFX2 U846 ( .A(n58), .Y(n757) );
  BUFX2 U847 ( .A(n42), .Y(n758) );
  BUFX2 U848 ( .A(n34), .Y(n759) );
  OR2X1 U849 ( .A(n249), .B(n262), .Y(n760) );
  OR2X1 U850 ( .A(n225), .B(n236), .Y(n761) );
  INVX1 U851 ( .A(n29), .Y(n139) );
  OR2X1 U852 ( .A(n323), .B(n328), .Y(n762) );
  OR2X1 U853 ( .A(n297), .B(n306), .Y(n763) );
  OR2X1 U854 ( .A(n329), .B(n334), .Y(n764) );
  OR2X1 U855 ( .A(n172), .B(n169), .Y(n765) );
  OR2X1 U856 ( .A(n196), .B(n189), .Y(n766) );
  OR2X1 U857 ( .A(n275), .B(n286), .Y(n767) );
  OR2X1 U858 ( .A(n177), .B(n182), .Y(n768) );
  OR2X1 U859 ( .A(n205), .B(n214), .Y(n769) );
  BUFX2 U860 ( .A(n302), .Y(n774) );
  OR2X1 U861 ( .A(n335), .B(n338), .Y(n770) );
  INVX1 U862 ( .A(b[15]), .Y(n802) );
  OR2X1 U863 ( .A(n343), .B(n344), .Y(n771) );
  AND2X1 U864 ( .A(b[4]), .B(b[0]), .Y(n459) );
  AND2X1 U865 ( .A(b[3]), .B(b[0]), .Y(n462) );
  INVX1 U866 ( .A(b[14]), .Y(n801) );
  INVX1 U867 ( .A(b[12]), .Y(n798) );
  INVX1 U868 ( .A(b[12]), .Y(n799) );
  XNOR2X1 U869 ( .A(n723), .B(n775), .Y(n303) );
  NAND3X1 U870 ( .A(n695), .B(n560), .C(n748), .Y(n776) );
  INVX1 U871 ( .A(n555), .Y(n116) );
  XOR2X1 U872 ( .A(n308), .B(n301), .Y(n778) );
  XOR2X1 U873 ( .A(n547), .B(n778), .Y(n297) );
  NAND3X1 U874 ( .A(n558), .B(n561), .C(n563), .Y(n302) );
  INVX1 U875 ( .A(n556), .Y(n94) );
  INVX1 U876 ( .A(n104), .Y(n103) );
endmodule


module alu_DW01_add_20 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n19, n75, n76;

  XOR2X1 U1 ( .A(n3), .B(n1), .Y(SUM[15]) );
  XOR2X1 U2 ( .A(A[15]), .B(B[15]), .Y(n1) );
  FAX1 U3 ( .A(B[14]), .B(A[14]), .C(n4), .YC(n3), .YS(SUM[14]) );
  FAX1 U4 ( .A(B[13]), .B(A[13]), .C(n5), .YC(n4), .YS(SUM[13]) );
  FAX1 U5 ( .A(B[12]), .B(A[12]), .C(n6), .YC(n5), .YS(SUM[12]) );
  FAX1 U6 ( .A(B[11]), .B(A[11]), .C(n7), .YC(n6), .YS(SUM[11]) );
  FAX1 U7 ( .A(B[10]), .B(A[10]), .C(n8), .YC(n7), .YS(SUM[10]) );
  FAX1 U8 ( .A(B[9]), .B(A[9]), .C(n9), .YC(n8), .YS(SUM[9]) );
  FAX1 U9 ( .A(B[8]), .B(A[8]), .C(n10), .YC(n9), .YS(SUM[8]) );
  FAX1 U10 ( .A(B[7]), .B(A[7]), .C(n11), .YC(n10), .YS(SUM[7]) );
  FAX1 U11 ( .A(B[6]), .B(A[6]), .C(n12), .YC(n11), .YS(SUM[6]) );
  FAX1 U12 ( .A(B[5]), .B(A[5]), .C(n13), .YC(n12), .YS(SUM[5]) );
  FAX1 U13 ( .A(A[4]), .B(B[4]), .C(n14), .YC(n13), .YS(SUM[4]) );
  FAX1 U14 ( .A(A[3]), .B(B[3]), .C(n15), .YC(n14), .YS(SUM[3]) );
  FAX1 U15 ( .A(A[2]), .B(B[2]), .C(n16), .YC(n15), .YS(SUM[2]) );
  FAX1 U16 ( .A(A[1]), .B(B[1]), .C(n19), .YC(n16), .YS(SUM[1]) );
  AND2X1 U26 ( .A(A[0]), .B(B[0]), .Y(n19) );
  AND2X1 U27 ( .A(n75), .B(n76), .Y(SUM[0]) );
  INVX1 U28 ( .A(n19), .Y(n75) );
  OR2X1 U29 ( .A(B[0]), .B(A[0]), .Y(n76) );
endmodule


module alu_DW01_add_18 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n19, n75, n76;

  XOR2X1 U1 ( .A(n3), .B(n1), .Y(SUM[15]) );
  XOR2X1 U2 ( .A(A[15]), .B(B[15]), .Y(n1) );
  FAX1 U3 ( .A(B[14]), .B(A[14]), .C(n4), .YC(n3), .YS(SUM[14]) );
  FAX1 U4 ( .A(B[13]), .B(A[13]), .C(n5), .YC(n4), .YS(SUM[13]) );
  FAX1 U5 ( .A(B[12]), .B(A[12]), .C(n6), .YC(n5), .YS(SUM[12]) );
  FAX1 U6 ( .A(B[11]), .B(A[11]), .C(n7), .YC(n6), .YS(SUM[11]) );
  FAX1 U7 ( .A(B[10]), .B(A[10]), .C(n8), .YC(n7), .YS(SUM[10]) );
  FAX1 U8 ( .A(B[9]), .B(A[9]), .C(n9), .YC(n8), .YS(SUM[9]) );
  FAX1 U9 ( .A(B[8]), .B(A[8]), .C(n10), .YC(n9), .YS(SUM[8]) );
  FAX1 U10 ( .A(B[7]), .B(A[7]), .C(n11), .YC(n10), .YS(SUM[7]) );
  FAX1 U11 ( .A(B[6]), .B(A[6]), .C(n12), .YC(n11), .YS(SUM[6]) );
  FAX1 U12 ( .A(A[5]), .B(B[5]), .C(n13), .YC(n12), .YS(SUM[5]) );
  FAX1 U13 ( .A(A[4]), .B(B[4]), .C(n14), .YC(n13), .YS(SUM[4]) );
  FAX1 U14 ( .A(A[3]), .B(B[3]), .C(n15), .YC(n14), .YS(SUM[3]) );
  FAX1 U15 ( .A(A[2]), .B(B[2]), .C(n16), .YC(n15), .YS(SUM[2]) );
  FAX1 U16 ( .A(A[1]), .B(B[1]), .C(n19), .YC(n16), .YS(SUM[1]) );
  AND2X1 U26 ( .A(n75), .B(n76), .Y(SUM[0]) );
  AND2X1 U27 ( .A(A[0]), .B(B[0]), .Y(n19) );
  INVX1 U28 ( .A(n19), .Y(n75) );
  OR2X1 U29 ( .A(B[0]), .B(A[0]), .Y(n76) );
endmodule


module alu_DW01_sub_19 ( A, B, CI, DIFF, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103;

  XOR2X1 U1 ( .A(n2), .B(n1), .Y(DIFF[15]) );
  FAX1 U3 ( .A(n103), .B(A[14]), .C(n3), .YC(n2), .YS(DIFF[14]) );
  FAX1 U4 ( .A(n102), .B(A[13]), .C(n4), .YC(n3), .YS(DIFF[13]) );
  FAX1 U5 ( .A(n101), .B(A[12]), .C(n5), .YC(n4), .YS(DIFF[12]) );
  FAX1 U6 ( .A(n100), .B(A[11]), .C(n6), .YC(n5), .YS(DIFF[11]) );
  FAX1 U7 ( .A(n99), .B(A[10]), .C(n7), .YC(n6), .YS(DIFF[10]) );
  FAX1 U8 ( .A(n98), .B(A[9]), .C(n8), .YC(n7), .YS(DIFF[9]) );
  FAX1 U9 ( .A(n97), .B(A[8]), .C(n9), .YC(n8), .YS(DIFF[8]) );
  FAX1 U10 ( .A(n96), .B(A[7]), .C(n10), .YC(n9), .YS(DIFF[7]) );
  FAX1 U11 ( .A(n95), .B(A[6]), .C(n11), .YC(n10), .YS(DIFF[6]) );
  FAX1 U12 ( .A(n94), .B(A[5]), .C(n12), .YC(n11), .YS(DIFF[5]) );
  FAX1 U13 ( .A(n93), .B(A[4]), .C(n13), .YC(n12), .YS(DIFF[4]) );
  FAX1 U14 ( .A(n92), .B(A[3]), .C(n14), .YC(n13), .YS(DIFF[3]) );
  FAX1 U15 ( .A(A[2]), .B(n91), .C(n15), .YC(n14), .YS(DIFF[2]) );
  FAX1 U16 ( .A(n90), .B(A[1]), .C(n88), .YC(n15), .YS(DIFF[1]) );
  XNOR2X1 U18 ( .A(A[0]), .B(n89), .Y(DIFF[0]) );
  INVX1 U39 ( .A(B[0]), .Y(n89) );
  INVX1 U40 ( .A(B[2]), .Y(n91) );
  OR2X1 U41 ( .A(A[0]), .B(n89), .Y(n88) );
  INVX1 U42 ( .A(B[3]), .Y(n92) );
  INVX1 U43 ( .A(B[8]), .Y(n97) );
  INVX1 U44 ( .A(B[10]), .Y(n99) );
  INVX1 U45 ( .A(B[9]), .Y(n98) );
  INVX1 U46 ( .A(B[11]), .Y(n100) );
  INVX1 U47 ( .A(B[7]), .Y(n96) );
  INVX1 U48 ( .A(B[12]), .Y(n101) );
  INVX1 U49 ( .A(B[5]), .Y(n94) );
  INVX1 U50 ( .A(B[6]), .Y(n95) );
  XNOR2X1 U51 ( .A(A[15]), .B(B[15]), .Y(n1) );
  INVX1 U52 ( .A(B[14]), .Y(n103) );
  INVX1 U53 ( .A(B[13]), .Y(n102) );
  INVX1 U54 ( .A(B[1]), .Y(n90) );
  INVX1 U55 ( .A(B[4]), .Y(n93) );
endmodule


module alu_DW01_sub_18 ( A, B, CI, DIFF, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102;

  XOR2X1 U1 ( .A(n2), .B(n1), .Y(DIFF[15]) );
  FAX1 U3 ( .A(n102), .B(A[14]), .C(n3), .YC(n2), .YS(DIFF[14]) );
  FAX1 U4 ( .A(n101), .B(A[13]), .C(n4), .YC(n3), .YS(DIFF[13]) );
  FAX1 U5 ( .A(n100), .B(A[12]), .C(n5), .YC(n4), .YS(DIFF[12]) );
  FAX1 U6 ( .A(n99), .B(A[11]), .C(n6), .YC(n5), .YS(DIFF[11]) );
  FAX1 U7 ( .A(n98), .B(A[10]), .C(n7), .YC(n6), .YS(DIFF[10]) );
  FAX1 U8 ( .A(n97), .B(A[9]), .C(n8), .YC(n7), .YS(DIFF[9]) );
  FAX1 U9 ( .A(n96), .B(A[8]), .C(n9), .YC(n8), .YS(DIFF[8]) );
  FAX1 U10 ( .A(n95), .B(A[7]), .C(n10), .YC(n9), .YS(DIFF[7]) );
  FAX1 U11 ( .A(n94), .B(A[6]), .C(n11), .YC(n10), .YS(DIFF[6]) );
  FAX1 U12 ( .A(A[5]), .B(n93), .C(n12), .YC(n11), .YS(DIFF[5]) );
  FAX1 U13 ( .A(A[4]), .B(n92), .C(n13), .YC(n12), .YS(DIFF[4]) );
  FAX1 U14 ( .A(A[3]), .B(n91), .C(n14), .YC(n13), .YS(DIFF[3]) );
  FAX1 U15 ( .A(A[2]), .B(n90), .C(n15), .YC(n14), .YS(DIFF[2]) );
  FAX1 U16 ( .A(A[1]), .B(n89), .C(n16), .YC(n15), .YS(DIFF[1]) );
  XNOR2X1 U18 ( .A(n88), .B(A[0]), .Y(DIFF[0]) );
  OR2X1 U39 ( .A(n88), .B(A[0]), .Y(n16) );
  INVX1 U40 ( .A(B[2]), .Y(n90) );
  INVX1 U41 ( .A(B[1]), .Y(n89) );
  INVX1 U42 ( .A(B[3]), .Y(n91) );
  INVX1 U43 ( .A(B[4]), .Y(n92) );
  INVX1 U44 ( .A(B[9]), .Y(n97) );
  INVX1 U45 ( .A(B[6]), .Y(n94) );
  INVX1 U46 ( .A(B[7]), .Y(n95) );
  INVX1 U47 ( .A(B[11]), .Y(n99) );
  INVX1 U48 ( .A(B[12]), .Y(n100) );
  XNOR2X1 U49 ( .A(A[15]), .B(B[15]), .Y(n1) );
  INVX1 U50 ( .A(B[14]), .Y(n102) );
  INVX1 U51 ( .A(B[13]), .Y(n101) );
  INVX1 U52 ( .A(B[5]), .Y(n93) );
  INVX1 U53 ( .A(B[0]), .Y(n88) );
  INVX1 U54 ( .A(B[10]), .Y(n98) );
  INVX1 U55 ( .A(B[8]), .Y(n96) );
endmodule


module alu_DW01_sub_21 ( A, B, CI, DIFF, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103;

  FAX1 U3 ( .A(n103), .B(A[14]), .C(n3), .YC(n2), .YS(DIFF[14]) );
  FAX1 U4 ( .A(n102), .B(A[13]), .C(n4), .YC(n3), .YS(DIFF[13]) );
  FAX1 U5 ( .A(n101), .B(A[12]), .C(n5), .YC(n4), .YS(DIFF[12]) );
  FAX1 U6 ( .A(n100), .B(A[11]), .C(n6), .YC(n5), .YS(DIFF[11]) );
  FAX1 U7 ( .A(n99), .B(A[10]), .C(n7), .YC(n6), .YS(DIFF[10]) );
  FAX1 U8 ( .A(n98), .B(A[9]), .C(n8), .YC(n7), .YS(DIFF[9]) );
  FAX1 U9 ( .A(n97), .B(A[8]), .C(n9), .YC(n8), .YS(DIFF[8]) );
  FAX1 U10 ( .A(n96), .B(A[7]), .C(n10), .YC(n9), .YS(DIFF[7]) );
  FAX1 U11 ( .A(n95), .B(A[6]), .C(n11), .YC(n10), .YS(DIFF[6]) );
  FAX1 U12 ( .A(n94), .B(A[5]), .C(n12), .YC(n11), .YS(DIFF[5]) );
  FAX1 U13 ( .A(n93), .B(A[4]), .C(n13), .YC(n12), .YS(DIFF[4]) );
  FAX1 U14 ( .A(n92), .B(A[3]), .C(n14), .YC(n13), .YS(DIFF[3]) );
  FAX1 U15 ( .A(A[2]), .B(n91), .C(n15), .YC(n14), .YS(DIFF[2]) );
  FAX1 U16 ( .A(n90), .B(A[1]), .C(n16), .YC(n15), .YS(DIFF[1]) );
  XNOR2X1 U18 ( .A(n89), .B(A[0]), .Y(DIFF[0]) );
  OR2X1 U39 ( .A(n89), .B(A[0]), .Y(n16) );
  INVX2 U40 ( .A(B[1]), .Y(n90) );
  INVX1 U41 ( .A(B[0]), .Y(n89) );
  XOR2X1 U42 ( .A(A[15]), .B(B[15]), .Y(n88) );
  XNOR2X1 U43 ( .A(n2), .B(n88), .Y(DIFF[15]) );
  INVX1 U44 ( .A(B[2]), .Y(n91) );
  INVX1 U45 ( .A(B[3]), .Y(n92) );
  INVX1 U46 ( .A(B[8]), .Y(n97) );
  INVX1 U47 ( .A(B[9]), .Y(n98) );
  INVX1 U48 ( .A(B[10]), .Y(n99) );
  INVX1 U49 ( .A(B[12]), .Y(n101) );
  INVX1 U50 ( .A(B[11]), .Y(n100) );
  INVX1 U51 ( .A(B[4]), .Y(n93) );
  INVX1 U52 ( .A(B[5]), .Y(n94) );
  INVX1 U53 ( .A(B[6]), .Y(n95) );
  INVX1 U54 ( .A(B[7]), .Y(n96) );
  INVX1 U55 ( .A(B[14]), .Y(n103) );
  INVX1 U56 ( .A(B[13]), .Y(n102) );
endmodule


module alu_DW01_sub_20 ( A, B, CI, DIFF, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102;

  XOR2X1 U1 ( .A(n2), .B(n1), .Y(DIFF[15]) );
  FAX1 U3 ( .A(n102), .B(A[14]), .C(n3), .YC(n2), .YS(DIFF[14]) );
  FAX1 U4 ( .A(n101), .B(A[13]), .C(n4), .YC(n3), .YS(DIFF[13]) );
  FAX1 U5 ( .A(n100), .B(A[12]), .C(n5), .YC(n4), .YS(DIFF[12]) );
  FAX1 U6 ( .A(n99), .B(A[11]), .C(n6), .YC(n5), .YS(DIFF[11]) );
  FAX1 U7 ( .A(n98), .B(A[10]), .C(n7), .YC(n6), .YS(DIFF[10]) );
  FAX1 U8 ( .A(n97), .B(A[9]), .C(n8), .YC(n7), .YS(DIFF[9]) );
  FAX1 U9 ( .A(n96), .B(A[8]), .C(n9), .YC(n8), .YS(DIFF[8]) );
  FAX1 U10 ( .A(n95), .B(A[7]), .C(n10), .YC(n9), .YS(DIFF[7]) );
  FAX1 U11 ( .A(n94), .B(A[6]), .C(n11), .YC(n10), .YS(DIFF[6]) );
  FAX1 U12 ( .A(n93), .B(A[5]), .C(n12), .YC(n11), .YS(DIFF[5]) );
  FAX1 U13 ( .A(A[4]), .B(n92), .C(n13), .YC(n12), .YS(DIFF[4]) );
  FAX1 U14 ( .A(A[3]), .B(n91), .C(n14), .YC(n13), .YS(DIFF[3]) );
  FAX1 U15 ( .A(A[2]), .B(n90), .C(n15), .YC(n14), .YS(DIFF[2]) );
  FAX1 U16 ( .A(A[1]), .B(n89), .C(n16), .YC(n15), .YS(DIFF[1]) );
  XNOR2X1 U18 ( .A(n88), .B(A[0]), .Y(DIFF[0]) );
  OR2X1 U39 ( .A(n88), .B(A[0]), .Y(n16) );
  INVX1 U40 ( .A(B[2]), .Y(n90) );
  INVX1 U41 ( .A(B[1]), .Y(n89) );
  INVX1 U42 ( .A(B[4]), .Y(n92) );
  INVX1 U43 ( .A(B[3]), .Y(n91) );
  INVX1 U44 ( .A(B[8]), .Y(n96) );
  INVX1 U45 ( .A(B[9]), .Y(n97) );
  INVX1 U46 ( .A(B[10]), .Y(n98) );
  INVX1 U47 ( .A(B[6]), .Y(n94) );
  INVX1 U48 ( .A(B[14]), .Y(n102) );
  INVX1 U49 ( .A(B[12]), .Y(n100) );
  INVX1 U50 ( .A(B[11]), .Y(n99) );
  INVX1 U51 ( .A(B[5]), .Y(n93) );
  INVX1 U52 ( .A(B[7]), .Y(n95) );
  INVX1 U53 ( .A(B[0]), .Y(n88) );
  XNOR2X1 U54 ( .A(A[15]), .B(B[15]), .Y(n1) );
  INVX1 U55 ( .A(B[13]), .Y(n101) );
endmodule


module alu_DW_mult_uns_29 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n16, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n147, n148, n149, n150, n151,
         n152, n153, n154, n155;
  assign product[0] = b[0];

  FAX1 U2 ( .A(a[7]), .B(n125), .C(n3), .YC(product[15]), .YS(product[14]) );
  FAX1 U3 ( .A(n138), .B(n18), .C(n4), .YC(n3), .YS(product[13]) );
  FAX1 U4 ( .A(n19), .B(n20), .C(n5), .YC(n4), .YS(product[12]) );
  FAX1 U5 ( .A(n21), .B(n22), .C(n6), .YC(n5), .YS(product[11]) );
  FAX1 U6 ( .A(n26), .B(n23), .C(n7), .YC(n6), .YS(product[10]) );
  FAX1 U7 ( .A(n30), .B(n27), .C(n8), .YC(n7), .YS(product[9]) );
  FAX1 U8 ( .A(n36), .B(n31), .C(n9), .YC(n8), .YS(product[8]) );
  FAX1 U9 ( .A(n40), .B(n37), .C(n10), .YC(n9), .YS(product[7]) );
  FAX1 U10 ( .A(n43), .B(n41), .C(n11), .YC(n10), .YS(product[6]) );
  FAX1 U11 ( .A(n46), .B(n45), .C(n12), .YC(n11), .YS(product[5]) );
  FAX1 U12 ( .A(n143), .B(n47), .C(n13), .YC(n12), .YS(product[4]) );
  HAX1 U13 ( .A(n126), .B(n16), .YC(n13), .YS(product[3]) );
  FAX1 U20 ( .A(a[6]), .B(n127), .C(n128), .YC(n18), .YS(n19) );
  FAX1 U21 ( .A(n144), .B(n145), .C(n24), .YC(n20), .YS(n21) );
  FAX1 U22 ( .A(n140), .B(n28), .C(n25), .YC(n22), .YS(n23) );
  FAX1 U23 ( .A(a[5]), .B(n131), .C(n130), .YC(n24), .YS(n25) );
  FAX1 U24 ( .A(n34), .B(n32), .C(n29), .YC(n26), .YS(n27) );
  FAX1 U25 ( .A(n134), .B(n133), .C(n132), .YC(n28), .YS(n29) );
  FAX1 U26 ( .A(n38), .B(n35), .C(n33), .YC(n30), .YS(n31) );
  FAX1 U27 ( .A(n137), .B(n136), .C(n135), .YC(n32), .YS(n33) );
  HAX1 U28 ( .A(a[4]), .B(n122), .YC(n34), .YS(n35) );
  FAX1 U29 ( .A(n139), .B(n42), .C(n39), .YC(n36), .YS(n37) );
  HAX1 U30 ( .A(n120), .B(n121), .YC(n38), .YS(n39) );
  FAX1 U31 ( .A(n142), .B(n141), .C(n44), .YC(n40), .YS(n41) );
  HAX1 U32 ( .A(a[3]), .B(n118), .YC(n42), .YS(n43) );
  HAX1 U33 ( .A(n124), .B(n123), .YC(n44), .YS(n45) );
  HAX1 U34 ( .A(a[2]), .B(n119), .YC(n46), .YS(n47) );
  INVX1 U80 ( .A(b[1]), .Y(n149) );
  OR2X1 U81 ( .A(n129), .B(a[1]), .Y(n147) );
  AND2X1 U82 ( .A(a[1]), .B(n129), .Y(n16) );
  INVX1 U83 ( .A(n16), .Y(n117) );
  OR2X1 U84 ( .A(n151), .B(n150), .Y(n70) );
  INVX1 U85 ( .A(n70), .Y(n118) );
  OR2X1 U86 ( .A(n151), .B(n148), .Y(n72) );
  INVX1 U87 ( .A(n72), .Y(n119) );
  OR2X1 U88 ( .A(n152), .B(n150), .Y(n67) );
  INVX1 U89 ( .A(n67), .Y(n120) );
  OR2X1 U90 ( .A(n149), .B(n153), .Y(n64) );
  INVX1 U91 ( .A(n64), .Y(n121) );
  OR2X1 U92 ( .A(n153), .B(n150), .Y(n63) );
  INVX1 U93 ( .A(n63), .Y(n122) );
  OR2X1 U94 ( .A(n149), .B(n151), .Y(n71) );
  INVX1 U95 ( .A(n71), .Y(n123) );
  OR2X1 U96 ( .A(n152), .B(n148), .Y(n69) );
  INVX1 U97 ( .A(n69), .Y(n124) );
  OR2X1 U98 ( .A(n155), .B(n154), .Y(n48) );
  INVX1 U99 ( .A(n48), .Y(n125) );
  OR2X1 U100 ( .A(n150), .B(n148), .Y(n74) );
  INVX1 U101 ( .A(n74), .Y(n126) );
  OR2X1 U102 ( .A(n155), .B(n152), .Y(n50) );
  INVX1 U103 ( .A(n50), .Y(n127) );
  OR2X1 U104 ( .A(n154), .B(n153), .Y(n55) );
  INVX1 U105 ( .A(n55), .Y(n128) );
  OR2X1 U106 ( .A(n149), .B(n148), .Y(n75) );
  INVX1 U107 ( .A(n75), .Y(n129) );
  OR2X1 U108 ( .A(n155), .B(n150), .Y(n52) );
  INVX1 U109 ( .A(n52), .Y(n130) );
  OR2X1 U110 ( .A(n153), .B(n152), .Y(n61) );
  INVX1 U111 ( .A(n61), .Y(n131) );
  OR2X1 U112 ( .A(n149), .B(n155), .Y(n53) );
  INVX1 U113 ( .A(n53), .Y(n132) );
  OR2X1 U114 ( .A(n154), .B(n150), .Y(n58) );
  INVX1 U115 ( .A(n58), .Y(n133) );
  OR2X1 U116 ( .A(n153), .B(n151), .Y(n62) );
  INVX1 U117 ( .A(n62), .Y(n134) );
  OR2X1 U118 ( .A(n149), .B(n154), .Y(n59) );
  INVX1 U119 ( .A(n59), .Y(n135) );
  OR2X1 U120 ( .A(n155), .B(n148), .Y(n54) );
  INVX1 U121 ( .A(n54), .Y(n136) );
  OR2X1 U122 ( .A(n151), .B(n152), .Y(n66) );
  INVX1 U123 ( .A(n66), .Y(n137) );
  OR2X1 U124 ( .A(n155), .B(n153), .Y(n49) );
  INVX1 U125 ( .A(n49), .Y(n138) );
  OR2X1 U126 ( .A(n154), .B(n148), .Y(n60) );
  INVX1 U127 ( .A(n60), .Y(n139) );
  OR2X1 U128 ( .A(n154), .B(n151), .Y(n57) );
  INVX1 U129 ( .A(n57), .Y(n140) );
  OR2X1 U130 ( .A(n149), .B(n152), .Y(n68) );
  INVX1 U131 ( .A(n68), .Y(n141) );
  OR2X1 U132 ( .A(n153), .B(n148), .Y(n65) );
  INVX1 U133 ( .A(n65), .Y(n142) );
  OR2X1 U134 ( .A(n149), .B(n150), .Y(n73) );
  INVX1 U135 ( .A(n73), .Y(n143) );
  OR2X1 U136 ( .A(n154), .B(n152), .Y(n56) );
  INVX1 U137 ( .A(n56), .Y(n144) );
  OR2X1 U138 ( .A(n155), .B(n151), .Y(n51) );
  INVX1 U139 ( .A(n51), .Y(n145) );
  AND2X1 U140 ( .A(n117), .B(n147), .Y(product[2]) );
  INVX1 U141 ( .A(a[5]), .Y(n153) );
  INVX1 U142 ( .A(b[2]), .Y(n150) );
  INVX1 U143 ( .A(b[7]), .Y(n155) );
  INVX1 U144 ( .A(b[3]), .Y(n151) );
  INVX1 U145 ( .A(b[4]), .Y(n152) );
  INVX1 U146 ( .A(b[6]), .Y(n154) );
  INVX1 U147 ( .A(b[0]), .Y(n148) );
endmodule


module alu_DW_mult_uns_31 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n16, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n147, n148, n149, n150, n151,
         n152, n153, n154, n155;
  assign product[0] = b[0];

  FAX1 U2 ( .A(a[7]), .B(n140), .C(n3), .YC(product[15]), .YS(product[14]) );
  FAX1 U3 ( .A(n145), .B(n18), .C(n4), .YC(n3), .YS(product[13]) );
  FAX1 U4 ( .A(n19), .B(n20), .C(n5), .YC(n4), .YS(product[12]) );
  FAX1 U5 ( .A(n21), .B(n22), .C(n6), .YC(n5), .YS(product[11]) );
  FAX1 U6 ( .A(n26), .B(n23), .C(n7), .YC(n6), .YS(product[10]) );
  FAX1 U7 ( .A(n30), .B(n27), .C(n8), .YC(n7), .YS(product[9]) );
  FAX1 U8 ( .A(n36), .B(n31), .C(n9), .YC(n8), .YS(product[8]) );
  FAX1 U9 ( .A(n40), .B(n37), .C(n10), .YC(n9), .YS(product[7]) );
  FAX1 U10 ( .A(n43), .B(n41), .C(n11), .YC(n10), .YS(product[6]) );
  FAX1 U11 ( .A(n46), .B(n45), .C(n12), .YC(n11), .YS(product[5]) );
  FAX1 U12 ( .A(n143), .B(n47), .C(n13), .YC(n12), .YS(product[4]) );
  HAX1 U13 ( .A(n123), .B(n16), .YC(n13), .YS(product[3]) );
  FAX1 U20 ( .A(a[6]), .B(n125), .C(n124), .YC(n18), .YS(n19) );
  FAX1 U21 ( .A(n132), .B(n131), .C(n24), .YC(n20), .YS(n21) );
  FAX1 U22 ( .A(n144), .B(n28), .C(n25), .YC(n22), .YS(n23) );
  FAX1 U23 ( .A(a[5]), .B(n134), .C(n133), .YC(n24), .YS(n25) );
  FAX1 U24 ( .A(n34), .B(n32), .C(n29), .YC(n26), .YS(n27) );
  FAX1 U25 ( .A(n128), .B(n127), .C(n126), .YC(n28), .YS(n29) );
  FAX1 U26 ( .A(n38), .B(n35), .C(n33), .YC(n30), .YS(n31) );
  FAX1 U27 ( .A(n137), .B(n138), .C(n136), .YC(n32), .YS(n33) );
  HAX1 U28 ( .A(a[4]), .B(n129), .YC(n34), .YS(n35) );
  FAX1 U29 ( .A(n135), .B(n42), .C(n39), .YC(n36), .YS(n37) );
  HAX1 U30 ( .A(n120), .B(n119), .YC(n38), .YS(n39) );
  FAX1 U31 ( .A(n142), .B(n141), .C(n44), .YC(n40), .YS(n41) );
  HAX1 U32 ( .A(a[3]), .B(n139), .YC(n42), .YS(n43) );
  HAX1 U33 ( .A(n122), .B(n121), .YC(n44), .YS(n45) );
  HAX1 U34 ( .A(a[2]), .B(n118), .YC(n46), .YS(n47) );
  OR2X1 U80 ( .A(n151), .B(n148), .Y(n72) );
  OR2X1 U81 ( .A(n155), .B(n150), .Y(n52) );
  OR2X1 U82 ( .A(n154), .B(n150), .Y(n58) );
  INVX2 U83 ( .A(b[3]), .Y(n151) );
  OR2X1 U84 ( .A(n153), .B(n150), .Y(n63) );
  OR2X1 U85 ( .A(n149), .B(n150), .Y(n73) );
  INVX1 U86 ( .A(b[1]), .Y(n149) );
  INVX1 U87 ( .A(b[2]), .Y(n150) );
  OR2X1 U88 ( .A(n130), .B(a[1]), .Y(n147) );
  AND2X1 U89 ( .A(a[1]), .B(n130), .Y(n16) );
  INVX1 U90 ( .A(n16), .Y(n117) );
  INVX1 U91 ( .A(n72), .Y(n118) );
  OR2X1 U92 ( .A(n149), .B(n153), .Y(n64) );
  INVX1 U93 ( .A(n64), .Y(n119) );
  OR2X1 U94 ( .A(n152), .B(n150), .Y(n67) );
  INVX1 U95 ( .A(n67), .Y(n120) );
  OR2X1 U96 ( .A(n149), .B(n151), .Y(n71) );
  INVX1 U97 ( .A(n71), .Y(n121) );
  OR2X1 U98 ( .A(n152), .B(n148), .Y(n69) );
  INVX1 U99 ( .A(n69), .Y(n122) );
  OR2X1 U100 ( .A(n150), .B(n148), .Y(n74) );
  INVX1 U101 ( .A(n74), .Y(n123) );
  OR2X1 U102 ( .A(n154), .B(n153), .Y(n55) );
  INVX1 U103 ( .A(n55), .Y(n124) );
  OR2X1 U104 ( .A(n155), .B(n152), .Y(n50) );
  INVX1 U105 ( .A(n50), .Y(n125) );
  OR2X1 U106 ( .A(n149), .B(n155), .Y(n53) );
  INVX1 U107 ( .A(n53), .Y(n126) );
  INVX1 U108 ( .A(n58), .Y(n127) );
  OR2X1 U109 ( .A(n153), .B(n151), .Y(n62) );
  INVX1 U110 ( .A(n62), .Y(n128) );
  INVX1 U111 ( .A(n63), .Y(n129) );
  OR2X1 U112 ( .A(n149), .B(n148), .Y(n75) );
  INVX1 U113 ( .A(n75), .Y(n130) );
  OR2X1 U114 ( .A(n155), .B(n151), .Y(n51) );
  INVX1 U115 ( .A(n51), .Y(n131) );
  OR2X1 U116 ( .A(n154), .B(n152), .Y(n56) );
  INVX1 U117 ( .A(n56), .Y(n132) );
  INVX1 U118 ( .A(n52), .Y(n133) );
  OR2X1 U119 ( .A(n153), .B(n152), .Y(n61) );
  INVX1 U120 ( .A(n61), .Y(n134) );
  OR2X1 U121 ( .A(n154), .B(n148), .Y(n60) );
  INVX1 U122 ( .A(n60), .Y(n135) );
  OR2X1 U123 ( .A(n149), .B(n154), .Y(n59) );
  INVX1 U124 ( .A(n59), .Y(n136) );
  OR2X1 U125 ( .A(n151), .B(n152), .Y(n66) );
  INVX1 U126 ( .A(n66), .Y(n137) );
  OR2X1 U127 ( .A(n155), .B(n148), .Y(n54) );
  INVX1 U128 ( .A(n54), .Y(n138) );
  OR2X1 U129 ( .A(n151), .B(n150), .Y(n70) );
  INVX1 U130 ( .A(n70), .Y(n139) );
  OR2X1 U131 ( .A(n155), .B(n154), .Y(n48) );
  INVX1 U132 ( .A(n48), .Y(n140) );
  OR2X1 U133 ( .A(n149), .B(n152), .Y(n68) );
  INVX1 U134 ( .A(n68), .Y(n141) );
  OR2X1 U135 ( .A(n153), .B(n148), .Y(n65) );
  INVX1 U136 ( .A(n65), .Y(n142) );
  INVX1 U137 ( .A(n73), .Y(n143) );
  OR2X1 U138 ( .A(n154), .B(n151), .Y(n57) );
  INVX1 U139 ( .A(n57), .Y(n144) );
  OR2X1 U140 ( .A(n155), .B(n153), .Y(n49) );
  INVX1 U141 ( .A(n49), .Y(n145) );
  INVX1 U142 ( .A(b[5]), .Y(n153) );
  INVX1 U143 ( .A(b[6]), .Y(n154) );
  INVX1 U144 ( .A(b[7]), .Y(n155) );
  AND2X1 U145 ( .A(n117), .B(n147), .Y(product[2]) );
  INVX1 U146 ( .A(b[4]), .Y(n152) );
  INVX1 U147 ( .A(b[0]), .Y(n148) );
endmodule


module alu_DW_mult_uns_30 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n16, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154;
  assign product[0] = b[0];

  FAX1 U2 ( .A(a[7]), .B(n128), .C(n3), .YC(product[15]), .YS(product[14]) );
  FAX1 U3 ( .A(n145), .B(n18), .C(n4), .YC(n3), .YS(product[13]) );
  FAX1 U4 ( .A(n19), .B(n20), .C(n5), .YC(n4), .YS(product[12]) );
  FAX1 U5 ( .A(n21), .B(n22), .C(n6), .YC(n5), .YS(product[11]) );
  FAX1 U6 ( .A(n26), .B(n23), .C(n7), .YC(n6), .YS(product[10]) );
  FAX1 U7 ( .A(n30), .B(n27), .C(n8), .YC(n7), .YS(product[9]) );
  FAX1 U8 ( .A(n36), .B(n31), .C(n9), .YC(n8), .YS(product[8]) );
  FAX1 U9 ( .A(n40), .B(n37), .C(n10), .YC(n9), .YS(product[7]) );
  FAX1 U10 ( .A(n43), .B(n41), .C(n11), .YC(n10), .YS(product[6]) );
  FAX1 U11 ( .A(n46), .B(n45), .C(n12), .YC(n11), .YS(product[5]) );
  FAX1 U12 ( .A(n143), .B(n47), .C(n13), .YC(n12), .YS(product[4]) );
  HAX1 U13 ( .A(n120), .B(n16), .YC(n13), .YS(product[3]) );
  FAX1 U20 ( .A(a[6]), .B(n122), .C(n121), .YC(n18), .YS(n19) );
  FAX1 U21 ( .A(n142), .B(n141), .C(n24), .YC(n20), .YS(n21) );
  FAX1 U22 ( .A(n136), .B(n28), .C(n25), .YC(n22), .YS(n23) );
  FAX1 U23 ( .A(a[5]), .B(n124), .C(n123), .YC(n24), .YS(n25) );
  FAX1 U24 ( .A(n34), .B(n32), .C(n29), .YC(n26), .YS(n27) );
  FAX1 U25 ( .A(n135), .B(n134), .C(n133), .YC(n28), .YS(n29) );
  FAX1 U26 ( .A(n38), .B(n35), .C(n33), .YC(n30), .YS(n31) );
  FAX1 U27 ( .A(n131), .B(n130), .C(n129), .YC(n32), .YS(n33) );
  HAX1 U28 ( .A(a[4]), .B(n139), .YC(n34), .YS(n35) );
  FAX1 U29 ( .A(n144), .B(n42), .C(n39), .YC(n36), .YS(n37) );
  HAX1 U30 ( .A(n127), .B(n126), .YC(n38), .YS(n39) );
  FAX1 U31 ( .A(n137), .B(n138), .C(n44), .YC(n40), .YS(n41) );
  HAX1 U32 ( .A(a[3]), .B(n117), .YC(n42), .YS(n43) );
  HAX1 U33 ( .A(n119), .B(n118), .YC(n44), .YS(n45) );
  HAX1 U34 ( .A(a[2]), .B(n125), .YC(n46), .YS(n47) );
  OR2X1 U80 ( .A(n150), .B(n151), .Y(n66) );
  OR2X1 U81 ( .A(n140), .B(a[1]), .Y(n146) );
  AND2X1 U82 ( .A(a[1]), .B(n140), .Y(n16) );
  AND2X1 U83 ( .A(n132), .B(n146), .Y(product[2]) );
  INVX2 U84 ( .A(b[3]), .Y(n150) );
  OR2X1 U85 ( .A(n150), .B(n149), .Y(n70) );
  INVX1 U86 ( .A(n70), .Y(n117) );
  OR2X1 U87 ( .A(n148), .B(n150), .Y(n71) );
  INVX1 U88 ( .A(n71), .Y(n118) );
  OR2X1 U89 ( .A(n151), .B(n147), .Y(n69) );
  INVX1 U90 ( .A(n69), .Y(n119) );
  OR2X1 U91 ( .A(n149), .B(n147), .Y(n74) );
  INVX1 U92 ( .A(n74), .Y(n120) );
  OR2X1 U93 ( .A(n153), .B(n152), .Y(n55) );
  INVX1 U94 ( .A(n55), .Y(n121) );
  OR2X1 U95 ( .A(n154), .B(n151), .Y(n50) );
  INVX1 U96 ( .A(n50), .Y(n122) );
  OR2X1 U97 ( .A(n154), .B(n149), .Y(n52) );
  INVX1 U98 ( .A(n52), .Y(n123) );
  OR2X1 U99 ( .A(n152), .B(n151), .Y(n61) );
  INVX1 U100 ( .A(n61), .Y(n124) );
  OR2X1 U101 ( .A(n150), .B(n147), .Y(n72) );
  INVX1 U102 ( .A(n72), .Y(n125) );
  OR2X1 U103 ( .A(n148), .B(n152), .Y(n64) );
  INVX1 U104 ( .A(n64), .Y(n126) );
  OR2X1 U105 ( .A(n151), .B(n149), .Y(n67) );
  INVX1 U106 ( .A(n67), .Y(n127) );
  OR2X1 U107 ( .A(n154), .B(n153), .Y(n48) );
  INVX1 U108 ( .A(n48), .Y(n128) );
  OR2X1 U109 ( .A(n148), .B(n153), .Y(n59) );
  INVX1 U110 ( .A(n59), .Y(n129) );
  OR2X1 U111 ( .A(n154), .B(n147), .Y(n54) );
  INVX1 U112 ( .A(n54), .Y(n130) );
  INVX1 U113 ( .A(n66), .Y(n131) );
  INVX1 U114 ( .A(n16), .Y(n132) );
  OR2X1 U115 ( .A(n148), .B(n154), .Y(n53) );
  INVX1 U116 ( .A(n53), .Y(n133) );
  OR2X1 U117 ( .A(n153), .B(n149), .Y(n58) );
  INVX1 U118 ( .A(n58), .Y(n134) );
  OR2X1 U119 ( .A(n152), .B(n150), .Y(n62) );
  INVX1 U120 ( .A(n62), .Y(n135) );
  OR2X1 U121 ( .A(n153), .B(n150), .Y(n57) );
  INVX1 U122 ( .A(n57), .Y(n136) );
  OR2X1 U123 ( .A(n152), .B(n147), .Y(n65) );
  INVX1 U124 ( .A(n65), .Y(n137) );
  OR2X1 U125 ( .A(n148), .B(n151), .Y(n68) );
  INVX1 U126 ( .A(n68), .Y(n138) );
  OR2X1 U127 ( .A(n152), .B(n149), .Y(n63) );
  INVX1 U128 ( .A(n63), .Y(n139) );
  OR2X1 U129 ( .A(n148), .B(n147), .Y(n75) );
  INVX1 U130 ( .A(n75), .Y(n140) );
  OR2X1 U131 ( .A(n154), .B(n150), .Y(n51) );
  INVX1 U132 ( .A(n51), .Y(n141) );
  OR2X1 U133 ( .A(n153), .B(n151), .Y(n56) );
  INVX1 U134 ( .A(n56), .Y(n142) );
  OR2X1 U135 ( .A(n148), .B(n149), .Y(n73) );
  INVX1 U136 ( .A(n73), .Y(n143) );
  OR2X1 U137 ( .A(n153), .B(n147), .Y(n60) );
  INVX1 U138 ( .A(n60), .Y(n144) );
  OR2X1 U139 ( .A(n154), .B(n152), .Y(n49) );
  INVX1 U140 ( .A(n49), .Y(n145) );
  INVX1 U141 ( .A(b[2]), .Y(n149) );
  INVX1 U142 ( .A(b[6]), .Y(n153) );
  INVX1 U143 ( .A(b[1]), .Y(n148) );
  INVX1 U144 ( .A(b[7]), .Y(n154) );
  INVX1 U145 ( .A(b[5]), .Y(n152) );
  INVX1 U146 ( .A(b[0]), .Y(n147) );
  INVX1 U147 ( .A(b[4]), .Y(n151) );
endmodule


module alu_DW_mult_uns_28 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n16, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n147, n148, n149, n150, n151,
         n152, n153, n154, n155;
  assign product[0] = b[0];

  FAX1 U2 ( .A(a[7]), .B(n128), .C(n3), .YC(product[15]), .YS(product[14]) );
  FAX1 U3 ( .A(n145), .B(n18), .C(n4), .YC(n3), .YS(product[13]) );
  FAX1 U4 ( .A(n19), .B(n20), .C(n5), .YC(n4), .YS(product[12]) );
  FAX1 U5 ( .A(n21), .B(n22), .C(n6), .YC(n5), .YS(product[11]) );
  FAX1 U6 ( .A(n26), .B(n23), .C(n7), .YC(n6), .YS(product[10]) );
  FAX1 U7 ( .A(n30), .B(n27), .C(n8), .YC(n7), .YS(product[9]) );
  FAX1 U8 ( .A(n36), .B(n31), .C(n9), .YC(n8), .YS(product[8]) );
  FAX1 U9 ( .A(n40), .B(n37), .C(n10), .YC(n9), .YS(product[7]) );
  FAX1 U10 ( .A(n43), .B(n41), .C(n11), .YC(n10), .YS(product[6]) );
  FAX1 U11 ( .A(n46), .B(n45), .C(n12), .YC(n11), .YS(product[5]) );
  FAX1 U12 ( .A(n143), .B(n47), .C(n13), .YC(n12), .YS(product[4]) );
  HAX1 U13 ( .A(n120), .B(n16), .YC(n13), .YS(product[3]) );
  FAX1 U20 ( .A(a[6]), .B(n122), .C(n121), .YC(n18), .YS(n19) );
  FAX1 U21 ( .A(n139), .B(n138), .C(n24), .YC(n20), .YS(n21) );
  FAX1 U22 ( .A(n140), .B(n28), .C(n25), .YC(n22), .YS(n23) );
  FAX1 U23 ( .A(a[5]), .B(n124), .C(n123), .YC(n24), .YS(n25) );
  FAX1 U24 ( .A(n34), .B(n32), .C(n29), .YC(n26), .YS(n27) );
  FAX1 U25 ( .A(n131), .B(n130), .C(n129), .YC(n28), .YS(n29) );
  FAX1 U26 ( .A(n38), .B(n35), .C(n33), .YC(n30), .YS(n31) );
  FAX1 U27 ( .A(n135), .B(n134), .C(n133), .YC(n32), .YS(n33) );
  HAX1 U28 ( .A(a[4]), .B(n136), .YC(n34), .YS(n35) );
  FAX1 U29 ( .A(n144), .B(n42), .C(n39), .YC(n36), .YS(n37) );
  HAX1 U30 ( .A(n127), .B(n126), .YC(n38), .YS(n39) );
  FAX1 U31 ( .A(n141), .B(n142), .C(n44), .YC(n40), .YS(n41) );
  HAX1 U32 ( .A(a[3]), .B(n117), .YC(n42), .YS(n43) );
  HAX1 U33 ( .A(n119), .B(n118), .YC(n44), .YS(n45) );
  HAX1 U34 ( .A(a[2]), .B(n125), .YC(n46), .YS(n47) );
  OR2X1 U80 ( .A(n149), .B(n148), .Y(n75) );
  INVX1 U81 ( .A(b[1]), .Y(n149) );
  AND2X1 U82 ( .A(n132), .B(n147), .Y(product[2]) );
  OR2X1 U83 ( .A(n137), .B(a[1]), .Y(n147) );
  OR2X1 U84 ( .A(n151), .B(n150), .Y(n70) );
  INVX1 U85 ( .A(n70), .Y(n117) );
  OR2X1 U86 ( .A(n149), .B(n151), .Y(n71) );
  INVX1 U87 ( .A(n71), .Y(n118) );
  OR2X1 U88 ( .A(n152), .B(n148), .Y(n69) );
  INVX1 U89 ( .A(n69), .Y(n119) );
  OR2X1 U90 ( .A(n150), .B(n148), .Y(n74) );
  INVX1 U91 ( .A(n74), .Y(n120) );
  OR2X1 U92 ( .A(n154), .B(n153), .Y(n55) );
  INVX1 U93 ( .A(n55), .Y(n121) );
  OR2X1 U94 ( .A(n155), .B(n152), .Y(n50) );
  INVX1 U95 ( .A(n50), .Y(n122) );
  OR2X1 U96 ( .A(n155), .B(n150), .Y(n52) );
  INVX1 U97 ( .A(n52), .Y(n123) );
  OR2X1 U98 ( .A(n153), .B(n152), .Y(n61) );
  INVX1 U99 ( .A(n61), .Y(n124) );
  OR2X1 U100 ( .A(n151), .B(n148), .Y(n72) );
  INVX1 U101 ( .A(n72), .Y(n125) );
  OR2X1 U102 ( .A(n149), .B(n153), .Y(n64) );
  INVX1 U103 ( .A(n64), .Y(n126) );
  OR2X1 U104 ( .A(n152), .B(n150), .Y(n67) );
  INVX1 U105 ( .A(n67), .Y(n127) );
  OR2X1 U106 ( .A(n155), .B(n154), .Y(n48) );
  INVX1 U107 ( .A(n48), .Y(n128) );
  OR2X1 U108 ( .A(n149), .B(n155), .Y(n53) );
  INVX1 U109 ( .A(n53), .Y(n129) );
  OR2X1 U110 ( .A(n154), .B(n150), .Y(n58) );
  INVX1 U111 ( .A(n58), .Y(n130) );
  OR2X1 U112 ( .A(n153), .B(n151), .Y(n62) );
  INVX1 U113 ( .A(n62), .Y(n131) );
  AND2X1 U114 ( .A(a[1]), .B(n137), .Y(n16) );
  INVX1 U115 ( .A(n16), .Y(n132) );
  OR2X1 U116 ( .A(n149), .B(n154), .Y(n59) );
  INVX1 U117 ( .A(n59), .Y(n133) );
  OR2X1 U118 ( .A(n155), .B(n148), .Y(n54) );
  INVX1 U119 ( .A(n54), .Y(n134) );
  OR2X1 U120 ( .A(n151), .B(n152), .Y(n66) );
  INVX1 U121 ( .A(n66), .Y(n135) );
  OR2X1 U122 ( .A(n153), .B(n150), .Y(n63) );
  INVX1 U123 ( .A(n63), .Y(n136) );
  INVX1 U124 ( .A(n75), .Y(n137) );
  OR2X1 U125 ( .A(n155), .B(n151), .Y(n51) );
  INVX1 U126 ( .A(n51), .Y(n138) );
  OR2X1 U127 ( .A(n154), .B(n152), .Y(n56) );
  INVX1 U128 ( .A(n56), .Y(n139) );
  OR2X1 U129 ( .A(n154), .B(n151), .Y(n57) );
  INVX1 U130 ( .A(n57), .Y(n140) );
  OR2X1 U131 ( .A(n153), .B(n148), .Y(n65) );
  INVX1 U132 ( .A(n65), .Y(n141) );
  OR2X1 U133 ( .A(n149), .B(n152), .Y(n68) );
  INVX1 U134 ( .A(n68), .Y(n142) );
  OR2X1 U135 ( .A(n149), .B(n150), .Y(n73) );
  INVX1 U136 ( .A(n73), .Y(n143) );
  OR2X1 U137 ( .A(n154), .B(n148), .Y(n60) );
  INVX1 U138 ( .A(n60), .Y(n144) );
  OR2X1 U139 ( .A(n155), .B(n153), .Y(n49) );
  INVX1 U140 ( .A(n49), .Y(n145) );
  INVX1 U141 ( .A(b[2]), .Y(n150) );
  INVX1 U142 ( .A(b[5]), .Y(n153) );
  INVX1 U143 ( .A(b[6]), .Y(n154) );
  INVX1 U144 ( .A(b[7]), .Y(n155) );
  INVX1 U145 ( .A(b[0]), .Y(n148) );
  INVX1 U146 ( .A(b[4]), .Y(n152) );
  INVX1 U147 ( .A(b[3]), .Y(n151) );
endmodule


module alu_DW01_add_25 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n19, n75, n77;

  XOR2X1 U1 ( .A(n3), .B(n1), .Y(SUM[15]) );
  XOR2X1 U2 ( .A(A[15]), .B(B[15]), .Y(n1) );
  FAX1 U3 ( .A(B[14]), .B(A[14]), .C(n4), .YC(n3), .YS(SUM[14]) );
  FAX1 U4 ( .A(B[13]), .B(A[13]), .C(n5), .YC(n4), .YS(SUM[13]) );
  FAX1 U5 ( .A(B[12]), .B(A[12]), .C(n6), .YC(n5), .YS(SUM[12]) );
  FAX1 U6 ( .A(B[11]), .B(A[11]), .C(n7), .YC(n6), .YS(SUM[11]) );
  FAX1 U7 ( .A(B[10]), .B(A[10]), .C(n8), .YC(n7), .YS(SUM[10]) );
  FAX1 U8 ( .A(B[9]), .B(A[9]), .C(n9), .YC(n8), .YS(SUM[9]) );
  FAX1 U9 ( .A(A[8]), .B(B[8]), .C(n10), .YC(n9), .YS(SUM[8]) );
  FAX1 U10 ( .A(A[7]), .B(B[7]), .C(n11), .YC(n10), .YS(SUM[7]) );
  FAX1 U11 ( .A(A[6]), .B(B[6]), .C(n12), .YC(n11), .YS(SUM[6]) );
  FAX1 U12 ( .A(A[5]), .B(B[5]), .C(n13), .YC(n12), .YS(SUM[5]) );
  FAX1 U13 ( .A(A[4]), .B(B[4]), .C(n14), .YC(n13), .YS(SUM[4]) );
  FAX1 U14 ( .A(A[3]), .B(B[3]), .C(n15), .YC(n14), .YS(SUM[3]) );
  FAX1 U15 ( .A(A[2]), .B(B[2]), .C(n16), .YC(n15), .YS(SUM[2]) );
  FAX1 U16 ( .A(A[1]), .B(B[1]), .C(n19), .YC(n16), .YS(SUM[1]) );
  AND2X1 U26 ( .A(n75), .B(n77), .Y(SUM[0]) );
  AND2X1 U27 ( .A(A[0]), .B(B[0]), .Y(n19) );
  OR2X2 U28 ( .A(B[0]), .B(A[0]), .Y(n77) );
  INVX1 U29 ( .A(n19), .Y(n75) );
endmodule


module alu_DW01_add_26 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n19, n75, n77;

  XOR2X1 U1 ( .A(n3), .B(n1), .Y(SUM[15]) );
  XOR2X1 U2 ( .A(A[15]), .B(B[15]), .Y(n1) );
  FAX1 U3 ( .A(B[14]), .B(A[14]), .C(n4), .YC(n3), .YS(SUM[14]) );
  FAX1 U4 ( .A(B[13]), .B(A[13]), .C(n5), .YC(n4), .YS(SUM[13]) );
  FAX1 U5 ( .A(B[12]), .B(A[12]), .C(n6), .YC(n5), .YS(SUM[12]) );
  FAX1 U6 ( .A(B[11]), .B(A[11]), .C(n7), .YC(n6), .YS(SUM[11]) );
  FAX1 U7 ( .A(B[10]), .B(A[10]), .C(n8), .YC(n7), .YS(SUM[10]) );
  FAX1 U8 ( .A(B[9]), .B(A[9]), .C(n9), .YC(n8), .YS(SUM[9]) );
  FAX1 U9 ( .A(B[8]), .B(A[8]), .C(n10), .YC(n9), .YS(SUM[8]) );
  FAX1 U10 ( .A(A[7]), .B(B[7]), .C(n11), .YC(n10), .YS(SUM[7]) );
  FAX1 U11 ( .A(A[6]), .B(B[6]), .C(n12), .YC(n11), .YS(SUM[6]) );
  FAX1 U12 ( .A(A[5]), .B(B[5]), .C(n13), .YC(n12), .YS(SUM[5]) );
  FAX1 U13 ( .A(A[4]), .B(B[4]), .C(n14), .YC(n13), .YS(SUM[4]) );
  FAX1 U14 ( .A(A[3]), .B(B[3]), .C(n15), .YC(n14), .YS(SUM[3]) );
  FAX1 U15 ( .A(A[2]), .B(B[2]), .C(n16), .YC(n15), .YS(SUM[2]) );
  FAX1 U16 ( .A(A[1]), .B(B[1]), .C(n19), .YC(n16), .YS(SUM[1]) );
  OR2X2 U26 ( .A(B[0]), .B(A[0]), .Y(n77) );
  AND2X2 U27 ( .A(A[0]), .B(B[0]), .Y(n19) );
  AND2X1 U28 ( .A(n75), .B(n77), .Y(SUM[0]) );
  INVX1 U29 ( .A(n19), .Y(n75) );
endmodule


module alu_DW_mult_uns_105 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n2, n8, n9, n12, n14, n18, n20, n24, n26, n30, n32, n38, n42, n44,
         n46, n48, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n114, n115, n119, n120, n121, n125, n126, n127,
         n128, n129, n133, n134, n135, n136, n137, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n156, n157, n158,
         n159, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n201, n202, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n223, n224, n228, n229, n230, n234,
         n235, n236, n237, n238, n242, n243, n244, n245, n246, n250, n251,
         n252, n254, n255, n256, n268, n269, n275, n285, n286, n287, n288,
         n289, n291, n292, n293, n294, n295, n296, n297, n298, n299, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n411, n412, n413, n414, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n587, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n606, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n625, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n644, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n663, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n682, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n701, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n720, n721,
         n723, n725, n727, n729, n731, n733, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265;

  FAX1 U87 ( .A(n288), .B(n291), .C(n255), .YC(n114), .YS(product[30]) );
  XNOR2X1 U89 ( .A(n120), .B(n1114), .Y(product[29]) );
  AOI21X1 U90 ( .A(n120), .B(n1166), .C(n119), .Y(n115) );
  FAX1 U97 ( .A(n296), .B(n301), .C(n256), .YC(n120), .YS(product[28]) );
  XNOR2X1 U99 ( .A(n1156), .B(n1135), .Y(product[27]) );
  AOI21X1 U100 ( .A(n126), .B(n1162), .C(n125), .Y(n121) );
  XOR2X1 U107 ( .A(n1032), .B(n1072), .Y(product[26]) );
  OAI21X1 U108 ( .A(n1033), .B(n1144), .C(n1118), .Y(n126) );
  XNOR2X1 U113 ( .A(n1157), .B(n1137), .Y(product[25]) );
  AOI21X1 U114 ( .A(n134), .B(n1163), .C(n133), .Y(n129) );
  XOR2X1 U121 ( .A(n1029), .B(n1090), .Y(product[24]) );
  OAI21X1 U122 ( .A(n1145), .B(n1030), .C(n1119), .Y(n134) );
  XNOR2X1 U127 ( .A(n1154), .B(n1136), .Y(product[23]) );
  AOI21X1 U128 ( .A(n142), .B(n1161), .C(n141), .Y(n137) );
  XOR2X1 U135 ( .A(n1027), .B(n1060), .Y(product[22]) );
  OAI21X1 U136 ( .A(n1120), .B(n1012), .C(n1098), .Y(n142) );
  XNOR2X1 U141 ( .A(n150), .B(n1115), .Y(product[21]) );
  AOI21X1 U142 ( .A(n165), .B(n1006), .C(n147), .Y(n145) );
  OAI21X1 U144 ( .A(n1148), .B(n1025), .C(n1076), .Y(n147) );
  XNOR2X1 U149 ( .A(n157), .B(n1067), .Y(product[20]) );
  OAI21X1 U150 ( .A(n1026), .B(n164), .C(n1025), .Y(n150) );
  AOI21X1 U152 ( .A(n1158), .B(n159), .C(n156), .Y(n152) );
  XOR2X1 U159 ( .A(n164), .B(n1089), .Y(product[19]) );
  OAI21X1 U160 ( .A(n1121), .B(n164), .C(n1146), .Y(n157) );
  XNOR2X1 U169 ( .A(n172), .B(n1046), .Y(product[18]) );
  OAI21X1 U171 ( .A(n1011), .B(n1008), .C(n1016), .Y(n165) );
  AOI21X1 U173 ( .A(n991), .B(n177), .C(n169), .Y(n167) );
  OAI21X1 U175 ( .A(n1151), .B(n1106), .C(n1053), .Y(n169) );
  XOR2X1 U180 ( .A(n1080), .B(n1052), .Y(product[17]) );
  OAI21X1 U181 ( .A(n1125), .B(n1080), .C(n1151), .Y(n172) );
  XOR2X1 U186 ( .A(n1051), .B(n1050), .Y(product[16]) );
  AOI21X1 U187 ( .A(n185), .B(n1063), .C(n177), .Y(n175) );
  OAI21X1 U189 ( .A(n1147), .B(n1103), .C(n1062), .Y(n177) );
  XNOR2X1 U194 ( .A(n185), .B(n1087), .Y(product[15]) );
  AOI21X1 U195 ( .A(n185), .B(n183), .C(n184), .Y(n180) );
  XNOR2X1 U202 ( .A(n191), .B(n1021), .Y(product[14]) );
  AOI21X1 U204 ( .A(n195), .B(n1017), .C(n188), .Y(n186) );
  OAI21X1 U206 ( .A(n1150), .B(n1102), .C(n1078), .Y(n188) );
  XOR2X1 U211 ( .A(n194), .B(n1088), .Y(product[13]) );
  OAI21X1 U212 ( .A(n1124), .B(n194), .C(n1150), .Y(n191) );
  XOR2X1 U217 ( .A(n1071), .B(n1070), .Y(product[12]) );
  OAI21X1 U219 ( .A(n1019), .B(n1024), .C(n1014), .Y(n195) );
  AOI21X1 U221 ( .A(n1160), .B(n206), .C(n201), .Y(n197) );
  XNOR2X1 U228 ( .A(n207), .B(n1113), .Y(product[11]) );
  AOI21X1 U229 ( .A(n207), .B(n1164), .C(n206), .Y(n202) );
  XNOR2X1 U236 ( .A(n213), .B(n1059), .Y(product[10]) );
  AOI21X1 U238 ( .A(n1018), .B(n217), .C(n210), .Y(n208) );
  OAI21X1 U240 ( .A(n1149), .B(n1101), .C(n1077), .Y(n210) );
  XOR2X1 U245 ( .A(n1086), .B(n216), .Y(product[9]) );
  OAI21X1 U246 ( .A(n1123), .B(n216), .C(n1149), .Y(n213) );
  XOR2X1 U251 ( .A(n1069), .B(n1068), .Y(product[8]) );
  OAI21X1 U253 ( .A(n1010), .B(n1020), .C(n1013), .Y(n217) );
  AOI21X1 U255 ( .A(n1165), .B(n228), .C(n223), .Y(n219) );
  XNOR2X1 U262 ( .A(n229), .B(n1112), .Y(product[7]) );
  AOI21X1 U263 ( .A(n229), .B(n1159), .C(n228), .Y(n224) );
  XNOR2X1 U270 ( .A(n1066), .B(n235), .Y(product[6]) );
  AOI21X1 U272 ( .A(n235), .B(n1167), .C(n234), .Y(n230) );
  XOR2X1 U279 ( .A(n1009), .B(n1085), .Y(product[5]) );
  OAI21X1 U280 ( .A(n1009), .B(n1143), .C(n1117), .Y(n235) );
  XNOR2X1 U285 ( .A(n1056), .B(n243), .Y(product[4]) );
  AOI21X1 U286 ( .A(n243), .B(n1168), .C(n242), .Y(n238) );
  XOR2X1 U293 ( .A(n1058), .B(n1122), .Y(product[3]) );
  OAI21X1 U294 ( .A(n1142), .B(n1122), .C(n1097), .Y(n243) );
  XNOR2X1 U299 ( .A(n1057), .B(n1099), .Y(product[2]) );
  AOI21X1 U300 ( .A(n1169), .B(n1099), .C(n250), .Y(n246) );
  XOR2X1 U307 ( .A(n1153), .B(n252), .Y(product[1]) );
  XOR2X1 U315 ( .A(n1054), .B(n285), .Y(n286) );
  FAX1 U317 ( .A(n289), .B(n754), .C(n293), .YC(n287), .YS(n288) );
  FAX1 U319 ( .A(n755), .B(n294), .C(n297), .YC(n291), .YS(n292) );
  FAX1 U320 ( .A(n1126), .B(n1041), .C(n996), .YC(n293), .YS(n294) );
  FAX1 U321 ( .A(n756), .B(n298), .C(n303), .YC(n295), .YS(n296) );
  FAX1 U322 ( .A(n299), .B(n772), .C(n305), .YC(n297), .YS(n298) );
  FAX1 U324 ( .A(n311), .B(n304), .C(n309), .YC(n301), .YS(n302) );
  FAX1 U325 ( .A(n773), .B(n757), .C(n306), .YC(n303), .YS(n304) );
  FAX1 U326 ( .A(n1152), .B(n1042), .C(n1035), .YC(n305), .YS(n306) );
  FAX1 U327 ( .A(n319), .B(n310), .C(n317), .YC(n307), .YS(n308) );
  FAX1 U328 ( .A(n774), .B(n758), .C(n312), .YC(n309), .YS(n310) );
  FAX1 U329 ( .A(n313), .B(n790), .C(n321), .YC(n311), .YS(n312) );
  FAX1 U331 ( .A(n327), .B(n318), .C(n325), .YC(n315), .YS(n316) );
  FAX1 U332 ( .A(n775), .B(n329), .C(n320), .YC(n317), .YS(n318) );
  FAX1 U333 ( .A(n791), .B(n322), .C(n759), .YC(n319), .YS(n320) );
  FAX1 U334 ( .A(n807), .B(n1043), .C(n1064), .YC(n321), .YS(n322) );
  FAX1 U335 ( .A(n337), .B(n326), .C(n335), .YC(n323), .YS(n324) );
  FAX1 U336 ( .A(n330), .B(n339), .C(n328), .YC(n325), .YS(n326) );
  FAX1 U337 ( .A(n341), .B(n776), .C(n760), .YC(n327), .YS(n328) );
  FAX1 U338 ( .A(n331), .B(n808), .C(n792), .YC(n329), .YS(n330) );
  FAX1 U340 ( .A(n347), .B(n336), .C(n345), .YC(n333), .YS(n334) );
  FAX1 U341 ( .A(n349), .B(n340), .C(n338), .YC(n335), .YS(n336) );
  FAX1 U342 ( .A(n777), .B(n761), .C(n351), .YC(n337), .YS(n338) );
  FAX1 U343 ( .A(n809), .B(n793), .C(n342), .YC(n339), .YS(n340) );
  FAX1 U344 ( .A(n825), .B(n1081), .C(n1038), .YC(n341), .YS(n342) );
  FAX1 U345 ( .A(n348), .B(n357), .C(n346), .YC(n343), .YS(n344) );
  FAX1 U346 ( .A(n350), .B(n361), .C(n359), .YC(n345), .YS(n346) );
  FAX1 U347 ( .A(n778), .B(n352), .C(n363), .YC(n347), .YS(n348) );
  FAX1 U348 ( .A(n794), .B(n365), .C(n762), .YC(n349), .YS(n350) );
  FAX1 U349 ( .A(n353), .B(n826), .C(n810), .YC(n351), .YS(n352) );
  FAX1 U351 ( .A(n371), .B(n358), .C(n369), .YC(n355), .YS(n356) );
  FAX1 U352 ( .A(n362), .B(n373), .C(n360), .YC(n357), .YS(n358) );
  FAX1 U353 ( .A(n377), .B(n375), .C(n364), .YC(n359), .YS(n360) );
  FAX1 U354 ( .A(n811), .B(n779), .C(n763), .YC(n361), .YS(n362) );
  FAX1 U355 ( .A(n827), .B(n795), .C(n366), .YC(n363), .YS(n364) );
  FAX1 U356 ( .A(n843), .B(n1107), .C(n1040), .YC(n365), .YS(n366) );
  FAX1 U357 ( .A(n372), .B(n383), .C(n370), .YC(n367), .YS(n368) );
  FAX1 U358 ( .A(n374), .B(n387), .C(n385), .YC(n369), .YS(n370) );
  FAX1 U359 ( .A(n391), .B(n389), .C(n376), .YC(n371), .YS(n372) );
  FAX1 U360 ( .A(n780), .B(n764), .C(n378), .YC(n373), .YS(n374) );
  FAX1 U361 ( .A(n393), .B(n812), .C(n796), .YC(n375), .YS(n376) );
  FAX1 U362 ( .A(n379), .B(n844), .C(n828), .YC(n377), .YS(n378) );
  FAX1 U364 ( .A(n386), .B(n397), .C(n384), .YC(n381), .YS(n382) );
  FAX1 U365 ( .A(n401), .B(n388), .C(n399), .YC(n383), .YS(n384) );
  FAX1 U366 ( .A(n392), .B(n390), .C(n403), .YC(n385), .YS(n386) );
  FAX1 U367 ( .A(n765), .B(n407), .C(n405), .YC(n387), .YS(n388) );
  FAX1 U368 ( .A(n813), .B(n797), .C(n781), .YC(n389), .YS(n390) );
  FAX1 U369 ( .A(n829), .B(n394), .C(n845), .YC(n391), .YS(n392) );
  FAX1 U370 ( .A(n1248), .B(n9), .C(n1039), .YC(n393), .YS(n394) );
  FAX1 U371 ( .A(n400), .B(n413), .C(n398), .YC(n395), .YS(n396) );
  FAX1 U372 ( .A(n417), .B(n402), .C(n1096), .YC(n397), .YS(n398) );
  FAX1 U373 ( .A(n406), .B(n419), .C(n404), .YC(n399), .YS(n400) );
  FAX1 U374 ( .A(n408), .B(n423), .C(n421), .YC(n401), .YS(n402) );
  FAX1 U375 ( .A(n814), .B(n782), .C(n766), .YC(n403), .YS(n404) );
  FAX1 U376 ( .A(n830), .B(n798), .C(n846), .YC(n405), .YS(n406) );
  FAX1 U377 ( .A(a[1]), .B(n1079), .C(n862), .YC(n407), .YS(n408) );
  FAX1 U379 ( .A(n416), .B(n428), .C(n414), .YC(n411), .YS(n412) );
  FAX1 U380 ( .A(n432), .B(n418), .C(n430), .YC(n413), .YS(n414) );
  FAX1 U382 ( .A(n438), .B(n424), .C(n436), .YC(n417), .YS(n418) );
  FAX1 U383 ( .A(n1184), .B(n783), .C(n767), .YC(n419), .YS(n420) );
  FAX1 U384 ( .A(n863), .B(n815), .C(n847), .YC(n421), .YS(n422) );
  FAX1 U385 ( .A(a[1]), .B(n1047), .C(n831), .YC(n423), .YS(n424) );
  FAX1 U387 ( .A(n431), .B(n442), .C(n429), .YC(n426), .YS(n427) );
  FAX1 U388 ( .A(n446), .B(n433), .C(n444), .YC(n428), .YS(n429) );
  FAX1 U389 ( .A(n448), .B(n437), .C(n435), .YC(n430), .YS(n431) );
  FAX1 U390 ( .A(n452), .B(n439), .C(n1002), .YC(n432), .YS(n433) );
  FAX1 U391 ( .A(n800), .B(n784), .C(n768), .YC(n434), .YS(n435) );
  FAX1 U392 ( .A(n1193), .B(n864), .C(n848), .YC(n436), .YS(n437) );
  FAX1 U393 ( .A(n879), .B(n1044), .C(n832), .YC(n438), .YS(n439) );
  FAX1 U394 ( .A(n445), .B(n456), .C(n443), .YC(n440), .YS(n441) );
  FAX1 U395 ( .A(n460), .B(n447), .C(n458), .YC(n442), .YS(n443) );
  FAX1 U396 ( .A(n462), .B(n451), .C(n449), .YC(n444), .YS(n445) );
  FAX1 U397 ( .A(n466), .B(n453), .C(n464), .YC(n446), .YS(n447) );
  FAX1 U398 ( .A(n801), .B(n785), .C(n769), .YC(n448), .YS(n449) );
  HAX1 U400 ( .A(n880), .B(n833), .YC(n452), .YS(n453) );
  FAX1 U401 ( .A(n459), .B(n470), .C(n457), .YC(n454), .YS(n455) );
  FAX1 U402 ( .A(n463), .B(n461), .C(n472), .YC(n456), .YS(n457) );
  FAX1 U403 ( .A(n476), .B(n465), .C(n474), .YC(n458), .YS(n459) );
  FAX1 U404 ( .A(n786), .B(n478), .C(n467), .YC(n460), .YS(n461) );
  FAX1 U405 ( .A(n818), .B(n802), .C(n866), .YC(n462), .YS(n463) );
  FAX1 U406 ( .A(n735), .B(n850), .C(n770), .YC(n464), .YS(n465) );
  HAX1 U407 ( .A(n881), .B(n834), .YC(n466), .YS(n467) );
  FAX1 U408 ( .A(n473), .B(n482), .C(n471), .YC(n468), .YS(n469) );
  FAX1 U409 ( .A(n477), .B(n475), .C(n484), .YC(n470), .YS(n471) );
  FAX1 U410 ( .A(n479), .B(n488), .C(n486), .YC(n472), .YS(n473) );
  FAX1 U411 ( .A(n803), .B(n787), .C(n490), .YC(n474), .YS(n475) );
  FAX1 U412 ( .A(n819), .B(n867), .C(n851), .YC(n476), .YS(n477) );
  HAX1 U413 ( .A(n882), .B(n835), .YC(n478), .YS(n479) );
  FAX1 U414 ( .A(n485), .B(n494), .C(n483), .YC(n480), .YS(n481) );
  FAX1 U415 ( .A(n489), .B(n487), .C(n496), .YC(n482), .YS(n483) );
  FAX1 U416 ( .A(n500), .B(n491), .C(n498), .YC(n484), .YS(n485) );
  FAX1 U417 ( .A(n820), .B(n804), .C(n868), .YC(n486), .YS(n487) );
  FAX1 U418 ( .A(n736), .B(n852), .C(n788), .YC(n488), .YS(n489) );
  HAX1 U419 ( .A(n883), .B(n836), .YC(n490), .YS(n491) );
  FAX1 U420 ( .A(n497), .B(n504), .C(n495), .YC(n492), .YS(n493) );
  FAX1 U421 ( .A(n508), .B(n499), .C(n506), .YC(n494), .YS(n495) );
  FAX1 U422 ( .A(n805), .B(n510), .C(n501), .YC(n496), .YS(n497) );
  FAX1 U423 ( .A(n821), .B(n869), .C(n853), .YC(n498), .YS(n499) );
  HAX1 U424 ( .A(n884), .B(n837), .YC(n500), .YS(n501) );
  FAX1 U425 ( .A(n507), .B(n514), .C(n505), .YC(n502), .YS(n503) );
  FAX1 U426 ( .A(n511), .B(n516), .C(n509), .YC(n504), .YS(n505) );
  FAX1 U427 ( .A(n737), .B(n822), .C(n518), .YC(n506), .YS(n507) );
  FAX1 U428 ( .A(n838), .B(n870), .C(n854), .YC(n508), .YS(n509) );
  HAX1 U429 ( .A(n885), .B(n806), .YC(n510), .YS(n511) );
  FAX1 U430 ( .A(n517), .B(n522), .C(n515), .YC(n512), .YS(n513) );
  FAX1 U431 ( .A(n871), .B(n519), .C(n524), .YC(n514), .YS(n515) );
  FAX1 U432 ( .A(n823), .B(n855), .C(n526), .YC(n516), .YS(n517) );
  HAX1 U433 ( .A(n886), .B(n839), .YC(n518), .YS(n519) );
  FAX1 U434 ( .A(n525), .B(n530), .C(n523), .YC(n520), .YS(n521) );
  FAX1 U435 ( .A(n872), .B(n527), .C(n532), .YC(n522), .YS(n523) );
  FAX1 U436 ( .A(n824), .B(n840), .C(n856), .YC(n524), .YS(n525) );
  HAX1 U437 ( .A(n887), .B(n738), .YC(n526), .YS(n527) );
  FAX1 U438 ( .A(n533), .B(n536), .C(n531), .YC(n528), .YS(n529) );
  FAX1 U439 ( .A(n873), .B(n857), .C(n538), .YC(n530), .YS(n531) );
  HAX1 U440 ( .A(n888), .B(n841), .YC(n532), .YS(n533) );
  FAX1 U441 ( .A(n539), .B(n542), .C(n537), .YC(n534), .YS(n535) );
  FAX1 U442 ( .A(n842), .B(n874), .C(n858), .YC(n536), .YS(n537) );
  HAX1 U443 ( .A(n889), .B(n739), .YC(n538), .YS(n539) );
  FAX1 U444 ( .A(n859), .B(n546), .C(n543), .YC(n540), .YS(n541) );
  HAX1 U445 ( .A(n890), .B(n875), .YC(n542), .YS(n543) );
  FAX1 U446 ( .A(n860), .B(n876), .C(n547), .YC(n544), .YS(n545) );
  HAX1 U447 ( .A(n891), .B(n740), .YC(n546), .YS(n547) );
  HAX1 U448 ( .A(n892), .B(n877), .YC(n548), .YS(n549) );
  HAX1 U449 ( .A(n893), .B(n741), .YC(n550), .YS(n551) );
  MUX2X1 U451 ( .B(b[15]), .A(b[14]), .S(n1257), .Y(n552) );
  MUX2X1 U453 ( .B(b[14]), .A(b[13]), .S(n1257), .Y(n553) );
  MUX2X1 U455 ( .B(b[13]), .A(n1242), .S(n1258), .Y(n554) );
  MUX2X1 U457 ( .B(n1242), .A(b[11]), .S(n1258), .Y(n555) );
  MUX2X1 U459 ( .B(b[11]), .A(n1240), .S(n1258), .Y(n556) );
  MUX2X1 U461 ( .B(n1240), .A(n1238), .S(n1258), .Y(n557) );
  MUX2X1 U463 ( .B(n1238), .A(b[8]), .S(n1258), .Y(n558) );
  MUX2X1 U465 ( .B(b[8]), .A(n1235), .S(n1258), .Y(n559) );
  MUX2X1 U467 ( .B(n1235), .A(n1233), .S(n1258), .Y(n560) );
  MUX2X1 U469 ( .B(n1233), .A(n1231), .S(n1257), .Y(n561) );
  MUX2X1 U471 ( .B(n1231), .A(n1229), .S(n1257), .Y(n562) );
  MUX2X1 U473 ( .B(n1229), .A(n1227), .S(n1258), .Y(n563) );
  MUX2X1 U475 ( .B(n1227), .A(n1225), .S(n1258), .Y(n564) );
  MUX2X1 U477 ( .B(n1225), .A(n1222), .S(n1258), .Y(n565) );
  MUX2X1 U479 ( .B(n1222), .A(n1220), .S(n1258), .Y(n566) );
  MUX2X1 U486 ( .B(n1219), .A(n46), .S(n1065), .Y(n754) );
  MUX2X1 U488 ( .B(n1219), .A(n46), .S(n571), .Y(n755) );
  MUX2X1 U489 ( .B(b[15]), .A(b[14]), .S(n1217), .Y(n571) );
  MUX2X1 U490 ( .B(n1219), .A(n46), .S(n572), .Y(n756) );
  MUX2X1 U491 ( .B(b[14]), .A(b[13]), .S(n1217), .Y(n572) );
  MUX2X1 U492 ( .B(n1219), .A(n46), .S(n573), .Y(n757) );
  MUX2X1 U493 ( .B(b[13]), .A(n1242), .S(n1217), .Y(n573) );
  MUX2X1 U494 ( .B(n1219), .A(n46), .S(n574), .Y(n758) );
  MUX2X1 U495 ( .B(n1242), .A(b[11]), .S(n1217), .Y(n574) );
  MUX2X1 U496 ( .B(n1219), .A(n46), .S(n575), .Y(n759) );
  MUX2X1 U497 ( .B(b[11]), .A(n1240), .S(n1217), .Y(n575) );
  MUX2X1 U498 ( .B(n1219), .A(n46), .S(n576), .Y(n760) );
  MUX2X1 U499 ( .B(n1240), .A(n1238), .S(n1217), .Y(n576) );
  MUX2X1 U500 ( .B(n1219), .A(n46), .S(n577), .Y(n761) );
  MUX2X1 U501 ( .B(n1238), .A(b[8]), .S(n1217), .Y(n577) );
  MUX2X1 U502 ( .B(n1218), .A(n46), .S(n578), .Y(n762) );
  MUX2X1 U503 ( .B(b[8]), .A(n1235), .S(n1217), .Y(n578) );
  MUX2X1 U504 ( .B(n1218), .A(n46), .S(n579), .Y(n763) );
  MUX2X1 U505 ( .B(n1235), .A(n1233), .S(n1217), .Y(n579) );
  MUX2X1 U506 ( .B(n1218), .A(n46), .S(n580), .Y(n764) );
  MUX2X1 U507 ( .B(n1233), .A(n1231), .S(n1217), .Y(n580) );
  MUX2X1 U508 ( .B(n1218), .A(n46), .S(n581), .Y(n765) );
  MUX2X1 U509 ( .B(n1231), .A(n1229), .S(n1217), .Y(n581) );
  MUX2X1 U510 ( .B(n1218), .A(n46), .S(n582), .Y(n766) );
  MUX2X1 U511 ( .B(n1229), .A(n1227), .S(n48), .Y(n582) );
  MUX2X1 U512 ( .B(n1218), .A(n46), .S(n583), .Y(n767) );
  MUX2X1 U514 ( .B(n1218), .A(n46), .S(n584), .Y(n768) );
  MUX2X1 U515 ( .B(n1225), .A(n1222), .S(n48), .Y(n584) );
  MUX2X1 U516 ( .B(n1218), .A(n46), .S(n585), .Y(n769) );
  MUX2X1 U517 ( .B(n1222), .A(n1220), .S(n48), .Y(n585) );
  MUX2X1 U518 ( .B(n1218), .A(n46), .S(n587), .Y(n770) );
  MUX2X1 U524 ( .B(n1216), .A(n996), .S(n1084), .Y(n772) );
  MUX2X1 U526 ( .B(n1216), .A(n996), .S(n590), .Y(n773) );
  MUX2X1 U527 ( .B(b[15]), .A(b[14]), .S(n1173), .Y(n590) );
  MUX2X1 U528 ( .B(n1216), .A(n996), .S(n591), .Y(n774) );
  MUX2X1 U529 ( .B(n1244), .A(b[13]), .S(n1173), .Y(n591) );
  MUX2X1 U530 ( .B(n1216), .A(n996), .S(n592), .Y(n775) );
  MUX2X1 U531 ( .B(b[13]), .A(n1242), .S(n1173), .Y(n592) );
  MUX2X1 U532 ( .B(n1216), .A(n996), .S(n593), .Y(n776) );
  MUX2X1 U533 ( .B(b[12]), .A(b[11]), .S(n1173), .Y(n593) );
  MUX2X1 U534 ( .B(n1216), .A(n996), .S(n594), .Y(n777) );
  MUX2X1 U535 ( .B(b[11]), .A(n1240), .S(n1173), .Y(n594) );
  MUX2X1 U536 ( .B(n1216), .A(n996), .S(n595), .Y(n778) );
  MUX2X1 U537 ( .B(b[10]), .A(n1238), .S(n1173), .Y(n595) );
  MUX2X1 U538 ( .B(n1216), .A(n996), .S(n596), .Y(n779) );
  MUX2X1 U539 ( .B(b[9]), .A(b[8]), .S(n1173), .Y(n596) );
  MUX2X1 U540 ( .B(n1215), .A(n996), .S(n597), .Y(n780) );
  MUX2X1 U541 ( .B(b[8]), .A(n1235), .S(n1214), .Y(n597) );
  MUX2X1 U542 ( .B(n1215), .A(n996), .S(n598), .Y(n781) );
  MUX2X1 U543 ( .B(n1236), .A(n1233), .S(n1214), .Y(n598) );
  MUX2X1 U544 ( .B(n1215), .A(n996), .S(n599), .Y(n782) );
  MUX2X1 U545 ( .B(b[6]), .A(n1231), .S(n1214), .Y(n599) );
  MUX2X1 U546 ( .B(n1215), .A(n995), .S(n600), .Y(n783) );
  MUX2X1 U547 ( .B(b[5]), .A(n1229), .S(n42), .Y(n600) );
  MUX2X1 U548 ( .B(n1215), .A(n995), .S(n601), .Y(n784) );
  MUX2X1 U549 ( .B(b[4]), .A(n1227), .S(n42), .Y(n601) );
  MUX2X1 U550 ( .B(n1215), .A(n996), .S(n602), .Y(n785) );
  MUX2X1 U551 ( .B(b[3]), .A(n1225), .S(n42), .Y(n602) );
  MUX2X1 U552 ( .B(n1215), .A(n996), .S(n603), .Y(n786) );
  MUX2X1 U553 ( .B(b[2]), .A(n1222), .S(n1214), .Y(n603) );
  MUX2X1 U554 ( .B(n1215), .A(n996), .S(n604), .Y(n787) );
  MUX2X1 U555 ( .B(n1223), .A(n1220), .S(n1214), .Y(n604) );
  MUX2X1 U556 ( .B(n1215), .A(n996), .S(n606), .Y(n788) );
  OR2X1 U557 ( .A(n42), .B(n1221), .Y(n606) );
  MUX2X1 U562 ( .B(n1213), .A(n1034), .S(n1049), .Y(n790) );
  MUX2X1 U564 ( .B(n1213), .A(n1034), .S(n609), .Y(n791) );
  MUX2X1 U565 ( .B(b[15]), .A(b[14]), .S(n1155), .Y(n609) );
  MUX2X1 U566 ( .B(n1213), .A(n1034), .S(n610), .Y(n792) );
  MUX2X1 U567 ( .B(n1244), .A(b[13]), .S(n1155), .Y(n610) );
  MUX2X1 U568 ( .B(n1213), .A(n1035), .S(n611), .Y(n793) );
  MUX2X1 U569 ( .B(b[13]), .A(n1242), .S(n1155), .Y(n611) );
  MUX2X1 U570 ( .B(n1213), .A(n1034), .S(n612), .Y(n794) );
  MUX2X1 U571 ( .B(n1242), .A(b[11]), .S(n1155), .Y(n612) );
  MUX2X1 U572 ( .B(n1213), .A(n1035), .S(n613), .Y(n795) );
  MUX2X1 U573 ( .B(b[11]), .A(n1240), .S(n1155), .Y(n613) );
  MUX2X1 U574 ( .B(n1213), .A(n1035), .S(n614), .Y(n796) );
  MUX2X1 U575 ( .B(b[10]), .A(n1238), .S(n1155), .Y(n614) );
  MUX2X1 U576 ( .B(n1213), .A(n1034), .S(n615), .Y(n797) );
  MUX2X1 U577 ( .B(b[9]), .A(b[8]), .S(n1155), .Y(n615) );
  MUX2X1 U578 ( .B(n1212), .A(n1034), .S(n616), .Y(n798) );
  MUX2X1 U579 ( .B(b[8]), .A(n1235), .S(n1155), .Y(n616) );
  MUX2X1 U581 ( .B(n1236), .A(n1233), .S(n1171), .Y(n617) );
  MUX2X1 U582 ( .B(n1212), .A(n1035), .S(n618), .Y(n800) );
  MUX2X1 U583 ( .B(n1233), .A(n1231), .S(n1155), .Y(n618) );
  MUX2X1 U584 ( .B(n1212), .A(n1034), .S(n619), .Y(n801) );
  MUX2X1 U585 ( .B(b[5]), .A(n1229), .S(n1155), .Y(n619) );
  MUX2X1 U586 ( .B(n1212), .A(n1035), .S(n620), .Y(n802) );
  MUX2X1 U587 ( .B(b[4]), .A(n1227), .S(n1155), .Y(n620) );
  MUX2X1 U588 ( .B(n1212), .A(n1034), .S(n621), .Y(n803) );
  MUX2X1 U589 ( .B(b[3]), .A(n1225), .S(n1155), .Y(n621) );
  MUX2X1 U590 ( .B(n1212), .A(n1035), .S(n622), .Y(n804) );
  MUX2X1 U591 ( .B(b[2]), .A(n1222), .S(n1155), .Y(n622) );
  MUX2X1 U592 ( .B(n1212), .A(n1034), .S(n623), .Y(n805) );
  MUX2X1 U593 ( .B(n1223), .A(n1220), .S(n1155), .Y(n623) );
  MUX2X1 U594 ( .B(n1212), .A(n1035), .S(n625), .Y(n806) );
  MUX2X1 U600 ( .B(n1211), .A(n807), .S(n1083), .Y(n808) );
  MUX2X1 U602 ( .B(n1211), .A(n807), .S(n628), .Y(n809) );
  MUX2X1 U603 ( .B(b[15]), .A(b[14]), .S(n1209), .Y(n628) );
  MUX2X1 U604 ( .B(n1211), .A(n807), .S(n629), .Y(n810) );
  MUX2X1 U605 ( .B(b[14]), .A(b[13]), .S(n1209), .Y(n629) );
  MUX2X1 U606 ( .B(n1211), .A(n807), .S(n630), .Y(n811) );
  MUX2X1 U607 ( .B(b[13]), .A(n1242), .S(n1209), .Y(n630) );
  MUX2X1 U608 ( .B(n1211), .A(n807), .S(n631), .Y(n812) );
  MUX2X1 U609 ( .B(n1242), .A(b[11]), .S(n1209), .Y(n631) );
  MUX2X1 U610 ( .B(n1211), .A(n807), .S(n632), .Y(n813) );
  MUX2X1 U611 ( .B(b[11]), .A(n1240), .S(n1209), .Y(n632) );
  MUX2X1 U612 ( .B(n1211), .A(n807), .S(n633), .Y(n814) );
  MUX2X1 U613 ( .B(n1240), .A(n1238), .S(n1209), .Y(n633) );
  MUX2X1 U614 ( .B(n1211), .A(n807), .S(n634), .Y(n815) );
  MUX2X1 U615 ( .B(n1238), .A(b[8]), .S(n1209), .Y(n634) );
  MUX2X1 U617 ( .B(b[8]), .A(n1235), .S(n1208), .Y(n635) );
  MUX2X1 U619 ( .B(n1235), .A(n1233), .S(n1208), .Y(n636) );
  MUX2X1 U620 ( .B(n1210), .A(n807), .S(n637), .Y(n818) );
  MUX2X1 U621 ( .B(n1233), .A(n1231), .S(n1208), .Y(n637) );
  MUX2X1 U622 ( .B(n1210), .A(n807), .S(n638), .Y(n819) );
  MUX2X1 U623 ( .B(n1231), .A(n1229), .S(n1208), .Y(n638) );
  MUX2X1 U624 ( .B(n1210), .A(n807), .S(n639), .Y(n820) );
  MUX2X1 U625 ( .B(n1229), .A(n1227), .S(n1208), .Y(n639) );
  MUX2X1 U626 ( .B(n1210), .A(n807), .S(n640), .Y(n821) );
  MUX2X1 U627 ( .B(n1227), .A(n1225), .S(n1208), .Y(n640) );
  MUX2X1 U628 ( .B(n1210), .A(n807), .S(n641), .Y(n822) );
  MUX2X1 U629 ( .B(n1225), .A(n1222), .S(n1208), .Y(n641) );
  MUX2X1 U630 ( .B(n1210), .A(n807), .S(n642), .Y(n823) );
  MUX2X1 U631 ( .B(n1222), .A(n1220), .S(n1208), .Y(n642) );
  MUX2X1 U632 ( .B(n1210), .A(n807), .S(n644), .Y(n824) );
  AND2X1 U635 ( .A(n1207), .B(n729), .Y(n739) );
  MUX2X1 U638 ( .B(n1207), .A(n825), .S(n1110), .Y(n826) );
  MUX2X1 U640 ( .B(n1207), .A(n825), .S(n647), .Y(n827) );
  MUX2X1 U641 ( .B(b[15]), .A(b[14]), .S(n1205), .Y(n647) );
  MUX2X1 U642 ( .B(n1207), .A(n825), .S(n648), .Y(n828) );
  MUX2X1 U643 ( .B(b[14]), .A(b[13]), .S(n1205), .Y(n648) );
  MUX2X1 U644 ( .B(n1207), .A(n825), .S(n649), .Y(n829) );
  MUX2X1 U645 ( .B(b[13]), .A(n1242), .S(n1205), .Y(n649) );
  MUX2X1 U646 ( .B(n1207), .A(n825), .S(n650), .Y(n830) );
  MUX2X1 U647 ( .B(n1242), .A(b[11]), .S(n1205), .Y(n650) );
  MUX2X1 U648 ( .B(n1207), .A(n825), .S(n651), .Y(n831) );
  MUX2X1 U649 ( .B(b[11]), .A(n1240), .S(n1205), .Y(n651) );
  MUX2X1 U650 ( .B(n1207), .A(n825), .S(n652), .Y(n832) );
  MUX2X1 U651 ( .B(n1240), .A(n1238), .S(n1205), .Y(n652) );
  MUX2X1 U652 ( .B(n1207), .A(n825), .S(n653), .Y(n833) );
  MUX2X1 U653 ( .B(n1238), .A(b[8]), .S(n1205), .Y(n653) );
  MUX2X1 U654 ( .B(n1206), .A(n825), .S(n654), .Y(n834) );
  MUX2X1 U655 ( .B(b[8]), .A(n1235), .S(n1204), .Y(n654) );
  MUX2X1 U656 ( .B(n1206), .A(n825), .S(n655), .Y(n835) );
  MUX2X1 U657 ( .B(n1235), .A(n1233), .S(n1204), .Y(n655) );
  MUX2X1 U658 ( .B(n1206), .A(n825), .S(n656), .Y(n836) );
  MUX2X1 U659 ( .B(n1233), .A(n1231), .S(n1204), .Y(n656) );
  MUX2X1 U660 ( .B(n1206), .A(n825), .S(n657), .Y(n837) );
  MUX2X1 U661 ( .B(n1231), .A(n1229), .S(n1204), .Y(n657) );
  MUX2X1 U662 ( .B(n1206), .A(n825), .S(n658), .Y(n838) );
  MUX2X1 U663 ( .B(n1229), .A(n1227), .S(n1204), .Y(n658) );
  MUX2X1 U664 ( .B(n1206), .A(n825), .S(n659), .Y(n839) );
  MUX2X1 U665 ( .B(n1227), .A(n1225), .S(n1204), .Y(n659) );
  MUX2X1 U666 ( .B(n1206), .A(n825), .S(n660), .Y(n840) );
  MUX2X1 U667 ( .B(n1225), .A(n1222), .S(n1204), .Y(n660) );
  MUX2X1 U668 ( .B(n1206), .A(n825), .S(n661), .Y(n841) );
  MUX2X1 U669 ( .B(n1222), .A(n1220), .S(n1204), .Y(n661) );
  MUX2X1 U670 ( .B(n1206), .A(n825), .S(n663), .Y(n842) );
  OR2X1 U671 ( .A(n1205), .B(n1221), .Y(n663) );
  AND2X1 U673 ( .A(n1203), .B(n731), .Y(n740) );
  MUX2X1 U676 ( .B(n1203), .A(n843), .S(n1133), .Y(n844) );
  MUX2X1 U678 ( .B(n1203), .A(n843), .S(n666), .Y(n845) );
  MUX2X1 U679 ( .B(b[15]), .A(b[14]), .S(n1201), .Y(n666) );
  MUX2X1 U680 ( .B(n1203), .A(n843), .S(n667), .Y(n846) );
  MUX2X1 U681 ( .B(n1244), .A(b[13]), .S(n1201), .Y(n667) );
  MUX2X1 U682 ( .B(n1203), .A(n843), .S(n668), .Y(n847) );
  MUX2X1 U683 ( .B(b[13]), .A(n1242), .S(n1201), .Y(n668) );
  MUX2X1 U684 ( .B(n1203), .A(n843), .S(n669), .Y(n848) );
  MUX2X1 U685 ( .B(n1242), .A(b[11]), .S(n1201), .Y(n669) );
  MUX2X1 U686 ( .B(n1203), .A(n843), .S(n670), .Y(n849) );
  MUX2X1 U687 ( .B(b[11]), .A(n1240), .S(n1201), .Y(n670) );
  MUX2X1 U688 ( .B(n1203), .A(n843), .S(n671), .Y(n850) );
  MUX2X1 U689 ( .B(b[10]), .A(n1238), .S(n1201), .Y(n671) );
  MUX2X1 U690 ( .B(n1203), .A(n843), .S(n672), .Y(n851) );
  MUX2X1 U691 ( .B(b[9]), .A(b[8]), .S(n1201), .Y(n672) );
  MUX2X1 U692 ( .B(n1202), .A(n843), .S(n673), .Y(n852) );
  MUX2X1 U693 ( .B(b[8]), .A(n1235), .S(n1200), .Y(n673) );
  MUX2X1 U694 ( .B(n1202), .A(n843), .S(n674), .Y(n853) );
  MUX2X1 U695 ( .B(n1236), .A(n1233), .S(n1200), .Y(n674) );
  MUX2X1 U696 ( .B(n1202), .A(n843), .S(n675), .Y(n854) );
  MUX2X1 U697 ( .B(b[6]), .A(n1231), .S(n1200), .Y(n675) );
  MUX2X1 U698 ( .B(n1202), .A(n843), .S(n676), .Y(n855) );
  MUX2X1 U699 ( .B(b[5]), .A(n1229), .S(n1200), .Y(n676) );
  MUX2X1 U700 ( .B(n1202), .A(n843), .S(n677), .Y(n856) );
  MUX2X1 U701 ( .B(b[4]), .A(n1227), .S(n1200), .Y(n677) );
  MUX2X1 U702 ( .B(n1202), .A(n843), .S(n678), .Y(n857) );
  MUX2X1 U703 ( .B(b[3]), .A(n1225), .S(n1200), .Y(n678) );
  MUX2X1 U704 ( .B(n1202), .A(n843), .S(n679), .Y(n858) );
  MUX2X1 U705 ( .B(b[2]), .A(n1222), .S(n1200), .Y(n679) );
  MUX2X1 U706 ( .B(n1202), .A(n843), .S(n680), .Y(n859) );
  MUX2X1 U707 ( .B(n1223), .A(n1220), .S(n1200), .Y(n680) );
  MUX2X1 U708 ( .B(n1202), .A(n843), .S(n682), .Y(n860) );
  OR2X1 U709 ( .A(n1201), .B(n1221), .Y(n682) );
  AND2X1 U711 ( .A(n1199), .B(n733), .Y(n741) );
  MUX2X1 U714 ( .B(n1199), .A(n9), .S(n1134), .Y(n862) );
  MUX2X1 U716 ( .B(n1199), .A(n9), .S(n685), .Y(n863) );
  MUX2X1 U717 ( .B(b[15]), .A(b[14]), .S(n1197), .Y(n685) );
  MUX2X1 U718 ( .B(n1199), .A(n9), .S(n686), .Y(n864) );
  MUX2X1 U719 ( .B(n1244), .A(b[13]), .S(n1197), .Y(n686) );
  MUX2X1 U720 ( .B(n1199), .A(n9), .S(n687), .Y(n865) );
  MUX2X1 U721 ( .B(b[13]), .A(n1242), .S(n1197), .Y(n687) );
  MUX2X1 U722 ( .B(n1199), .A(n9), .S(n688), .Y(n866) );
  MUX2X1 U723 ( .B(n1242), .A(b[11]), .S(n1197), .Y(n688) );
  MUX2X1 U724 ( .B(n1199), .A(n9), .S(n689), .Y(n867) );
  MUX2X1 U725 ( .B(b[11]), .A(n1240), .S(n1197), .Y(n689) );
  MUX2X1 U726 ( .B(n1199), .A(n9), .S(n690), .Y(n868) );
  MUX2X1 U727 ( .B(b[10]), .A(n1238), .S(n1197), .Y(n690) );
  MUX2X1 U728 ( .B(n1199), .A(n9), .S(n691), .Y(n869) );
  MUX2X1 U729 ( .B(b[9]), .A(b[8]), .S(n1197), .Y(n691) );
  MUX2X1 U730 ( .B(n1198), .A(n9), .S(n692), .Y(n870) );
  MUX2X1 U731 ( .B(b[8]), .A(n1235), .S(n1196), .Y(n692) );
  MUX2X1 U732 ( .B(n1198), .A(n9), .S(n693), .Y(n871) );
  MUX2X1 U733 ( .B(n1236), .A(n1233), .S(n1196), .Y(n693) );
  MUX2X1 U734 ( .B(n1198), .A(n9), .S(n694), .Y(n872) );
  MUX2X1 U735 ( .B(b[6]), .A(n1231), .S(n1196), .Y(n694) );
  MUX2X1 U736 ( .B(n1198), .A(n9), .S(n695), .Y(n873) );
  MUX2X1 U737 ( .B(b[5]), .A(n1229), .S(n1196), .Y(n695) );
  MUX2X1 U738 ( .B(n1198), .A(n9), .S(n696), .Y(n874) );
  MUX2X1 U739 ( .B(b[4]), .A(n1227), .S(n1196), .Y(n696) );
  MUX2X1 U740 ( .B(n1198), .A(n9), .S(n697), .Y(n875) );
  MUX2X1 U741 ( .B(b[3]), .A(n1225), .S(n1196), .Y(n697) );
  MUX2X1 U742 ( .B(n1198), .A(n9), .S(n698), .Y(n876) );
  MUX2X1 U743 ( .B(b[2]), .A(n1222), .S(n1196), .Y(n698) );
  MUX2X1 U744 ( .B(n1198), .A(n9), .S(n699), .Y(n877) );
  MUX2X1 U745 ( .B(n1223), .A(n1220), .S(n1196), .Y(n699) );
  MUX2X1 U746 ( .B(n1198), .A(n9), .S(n701), .Y(n878) );
  OR2X1 U747 ( .A(n1197), .B(n1221), .Y(n701) );
  AND2X1 U749 ( .A(n1195), .B(a[1]), .Y(n742) );
  MUX2X1 U752 ( .B(n1195), .A(n1248), .S(n1111), .Y(n879) );
  MUX2X1 U754 ( .B(n1195), .A(n1248), .S(n704), .Y(n880) );
  MUX2X1 U755 ( .B(b[15]), .A(b[14]), .S(n1246), .Y(n704) );
  MUX2X1 U756 ( .B(n1195), .A(n1248), .S(n705), .Y(n881) );
  MUX2X1 U757 ( .B(n1244), .A(b[13]), .S(n1246), .Y(n705) );
  MUX2X1 U758 ( .B(n1195), .A(n1248), .S(n706), .Y(n882) );
  MUX2X1 U759 ( .B(b[13]), .A(n1242), .S(n1246), .Y(n706) );
  MUX2X1 U760 ( .B(n1195), .A(n1248), .S(n707), .Y(n883) );
  MUX2X1 U761 ( .B(n1242), .A(b[11]), .S(n1246), .Y(n707) );
  MUX2X1 U762 ( .B(n1195), .A(n1248), .S(n708), .Y(n884) );
  MUX2X1 U763 ( .B(b[11]), .A(n1240), .S(n1246), .Y(n708) );
  MUX2X1 U764 ( .B(n1195), .A(n1248), .S(n709), .Y(n885) );
  MUX2X1 U765 ( .B(b[10]), .A(n1238), .S(n1246), .Y(n709) );
  MUX2X1 U766 ( .B(n1195), .A(n1248), .S(n710), .Y(n886) );
  MUX2X1 U767 ( .B(b[9]), .A(b[8]), .S(n1246), .Y(n710) );
  MUX2X1 U768 ( .B(n1194), .A(n1248), .S(n711), .Y(n887) );
  MUX2X1 U769 ( .B(b[8]), .A(n1235), .S(n1246), .Y(n711) );
  MUX2X1 U770 ( .B(n1194), .A(n1248), .S(n712), .Y(n888) );
  MUX2X1 U771 ( .B(n1236), .A(n1233), .S(n1246), .Y(n712) );
  MUX2X1 U772 ( .B(n1194), .A(n1248), .S(n713), .Y(n889) );
  MUX2X1 U773 ( .B(n1233), .A(n1231), .S(n1247), .Y(n713) );
  MUX2X1 U774 ( .B(n1194), .A(n1248), .S(n714), .Y(n890) );
  MUX2X1 U775 ( .B(b[5]), .A(n1229), .S(n1247), .Y(n714) );
  MUX2X1 U776 ( .B(n1194), .A(n1248), .S(n715), .Y(n891) );
  MUX2X1 U777 ( .B(b[4]), .A(n1227), .S(n1247), .Y(n715) );
  MUX2X1 U778 ( .B(n1194), .A(n1248), .S(n716), .Y(n892) );
  MUX2X1 U779 ( .B(b[3]), .A(n1225), .S(n1246), .Y(n716) );
  MUX2X1 U780 ( .B(n1194), .A(n1248), .S(n717), .Y(n893) );
  MUX2X1 U781 ( .B(b[2]), .A(n1222), .S(n1246), .Y(n717) );
  MUX2X1 U782 ( .B(n1194), .A(n1248), .S(n718), .Y(n894) );
  MUX2X1 U783 ( .B(n1223), .A(n1220), .S(n1246), .Y(n718) );
  MUX2X1 U784 ( .B(n1194), .A(n1248), .S(n720), .Y(n895) );
  OR2X1 U785 ( .A(n1247), .B(n1221), .Y(n720) );
  OAI21X1 U789 ( .A(n994), .B(a[13]), .C(n1258), .Y(n44) );
  OAI21X1 U794 ( .A(a[12]), .B(n1254), .C(n1256), .Y(n38) );
  OAI21X1 U799 ( .A(a[9]), .B(a[10]), .C(n1255), .Y(n32) );
  OAI21X1 U804 ( .A(a[8]), .B(a[7]), .C(n1253), .Y(n26) );
  XNOR2X1 U807 ( .A(a[7]), .B(a[8]), .Y(n30) );
  OAI21X1 U809 ( .A(a[6]), .B(n1250), .C(n1252), .Y(n20) );
  XNOR2X1 U812 ( .A(n1250), .B(a[6]), .Y(n24) );
  OAI21X1 U814 ( .A(a[4]), .B(a[3]), .C(n1251), .Y(n14) );
  XNOR2X1 U817 ( .A(a[3]), .B(a[4]), .Y(n18) );
  OAI21X1 U819 ( .A(a[2]), .B(a[1]), .C(n1249), .Y(n8) );
  XNOR2X1 U822 ( .A(a[1]), .B(a[2]), .Y(n12) );
  BUFX4 U829 ( .A(n48), .Y(n1217) );
  INVX2 U830 ( .A(n998), .Y(n48) );
  INVX2 U831 ( .A(n733), .Y(n9) );
  INVX1 U832 ( .A(a[11]), .Y(n1255) );
  BUFX2 U833 ( .A(n789), .Y(n1035) );
  INVX1 U834 ( .A(n751), .Y(n1047) );
  OR2X1 U835 ( .A(n566), .B(n1257), .Y(n751) );
  INVX1 U836 ( .A(n46), .Y(n569) );
  INVX1 U837 ( .A(n1237), .Y(n1235) );
  INVX1 U838 ( .A(a[5]), .Y(n1251) );
  AND2X1 U839 ( .A(n1212), .B(n1181), .Y(n1182) );
  AND2X1 U840 ( .A(n789), .B(n617), .Y(n1183) );
  AND2X1 U841 ( .A(n1254), .B(n1253), .Y(n1263) );
  OR2X1 U842 ( .A(n556), .B(n1258), .Y(n745) );
  OR2X1 U843 ( .A(n558), .B(n1258), .Y(n746) );
  AND2X1 U844 ( .A(n367), .B(n356), .Y(n149) );
  OR2X1 U845 ( .A(n481), .B(n492), .Y(n1160) );
  OR2X1 U846 ( .A(n493), .B(n502), .Y(n1164) );
  OR2X1 U847 ( .A(n521), .B(n528), .Y(n1165) );
  OR2X1 U848 ( .A(n529), .B(n534), .Y(n1159) );
  OR2X1 U849 ( .A(n565), .B(n1258), .Y(n750) );
  OR2X1 U850 ( .A(n568), .B(n1257), .Y(n752) );
  OR2X1 U851 ( .A(n1257), .B(n1221), .Y(n568) );
  AND2X1 U852 ( .A(b[15]), .B(n1209), .Y(n627) );
  OR2X1 U853 ( .A(n562), .B(n1257), .Y(n748) );
  AND2X1 U854 ( .A(b[15]), .B(n1205), .Y(n646) );
  INVX1 U855 ( .A(n749), .Y(n1039) );
  OR2X1 U856 ( .A(n564), .B(n1258), .Y(n749) );
  AND2X1 U857 ( .A(n849), .B(n865), .Y(n1177) );
  AND2X1 U858 ( .A(n865), .B(n1172), .Y(n1175) );
  OR2X1 U859 ( .A(n560), .B(n1257), .Y(n747) );
  INVX2 U860 ( .A(n1241), .Y(n1240) );
  AND2X1 U861 ( .A(n1219), .B(n569), .Y(n735) );
  AND2X1 U862 ( .A(n1216), .B(n723), .Y(n736) );
  OR2X1 U863 ( .A(n1155), .B(n1221), .Y(n625) );
  OR2X1 U864 ( .A(n1209), .B(n1221), .Y(n644) );
  AND2X1 U865 ( .A(a[7]), .B(n1251), .Y(n1261) );
  AND2X1 U866 ( .A(n1250), .B(n1249), .Y(n1260) );
  AND2X1 U867 ( .A(n434), .B(n422), .Y(n992) );
  AND2X1 U868 ( .A(n1129), .B(n1130), .Y(n1184) );
  AND2X1 U869 ( .A(n1213), .B(n725), .Y(n737) );
  INVX2 U870 ( .A(n731), .Y(n843) );
  BUFX2 U871 ( .A(n12), .Y(n1197) );
  OR2X1 U872 ( .A(n554), .B(n1258), .Y(n744) );
  AND2X1 U873 ( .A(b[15]), .B(n1173), .Y(n589) );
  AND2X1 U874 ( .A(b[15]), .B(n1155), .Y(n608) );
  AND2X1 U875 ( .A(n468), .B(n455), .Y(n190) );
  OR2X1 U876 ( .A(n503), .B(n512), .Y(n211) );
  AND2X1 U877 ( .A(a[0]), .B(n1248), .Y(n2) );
  OR2X1 U878 ( .A(n552), .B(n1257), .Y(n743) );
  AND2X1 U879 ( .A(n1158), .B(n158), .Y(n151) );
  AND2X1 U880 ( .A(n512), .B(n503), .Y(n212) );
  AND2X1 U881 ( .A(n1091), .B(n1162), .Y(n87) );
  AND2X1 U882 ( .A(n1092), .B(n1163), .Y(n89) );
  AND2X1 U883 ( .A(n1073), .B(n1161), .Y(n91) );
  AND2X1 U884 ( .A(n1076), .B(n148), .Y(n93) );
  AND2X1 U885 ( .A(n1061), .B(n1158), .Y(n94) );
  AND2X1 U886 ( .A(n1146), .B(n158), .Y(n95) );
  AND2X1 U887 ( .A(n1053), .B(n997), .Y(n96) );
  AND2X1 U888 ( .A(n1151), .B(n268), .Y(n97) );
  AND2X1 U889 ( .A(n1062), .B(n269), .Y(n98) );
  AND2X1 U890 ( .A(n1147), .B(n183), .Y(n99) );
  AND2X1 U891 ( .A(n1150), .B(n192), .Y(n101) );
  AND2X1 U892 ( .A(n1095), .B(n1160), .Y(n102) );
  AND2X1 U893 ( .A(n1141), .B(n1164), .Y(n103) );
  AND2X1 U894 ( .A(n1094), .B(n1165), .Y(n106) );
  AND2X1 U895 ( .A(n1140), .B(n1159), .Y(n107) );
  BUFX2 U896 ( .A(n165), .Y(n990) );
  BUFX2 U897 ( .A(n30), .Y(n1209) );
  INVX4 U898 ( .A(n1239), .Y(n1238) );
  INVX2 U899 ( .A(a[15]), .Y(n1258) );
  INVX2 U900 ( .A(n1243), .Y(n1242) );
  INVX1 U901 ( .A(a[7]), .Y(n1252) );
  INVX1 U902 ( .A(a[15]), .Y(n1257) );
  AND2X1 U903 ( .A(n502), .B(n493), .Y(n206) );
  INVX1 U904 ( .A(a[13]), .Y(n1256) );
  INVX1 U905 ( .A(b[14]), .Y(n1245) );
  AND2X1 U906 ( .A(n1003), .B(n1007), .Y(n1022) );
  INVX1 U907 ( .A(n725), .Y(n789) );
  INVX2 U908 ( .A(n1234), .Y(n1233) );
  AND2X1 U909 ( .A(n1109), .B(n1108), .Y(n1193) );
  OR2X1 U910 ( .A(n553), .B(n1258), .Y(n289) );
  OR2X1 U911 ( .A(n559), .B(n1258), .Y(n331) );
  OR2X1 U912 ( .A(n561), .B(n1257), .Y(n353) );
  OR2X1 U913 ( .A(n555), .B(n1257), .Y(n299) );
  OR2X1 U914 ( .A(n563), .B(n1257), .Y(n379) );
  OR2X1 U915 ( .A(n382), .B(n395), .Y(n158) );
  AND2X1 U916 ( .A(n395), .B(n382), .Y(n159) );
  AND2X1 U917 ( .A(n454), .B(n441), .Y(n184) );
  OR2X1 U918 ( .A(n513), .B(n520), .Y(n214) );
  OR2X1 U919 ( .A(n455), .B(n468), .Y(n189) );
  OR2X1 U920 ( .A(n469), .B(n480), .Y(n192) );
  AND2X1 U921 ( .A(n381), .B(n368), .Y(n156) );
  AND2X1 U922 ( .A(n528), .B(n521), .Y(n223) );
  AND2X1 U923 ( .A(n492), .B(n481), .Y(n201) );
  AND2X1 U924 ( .A(n534), .B(n529), .Y(n228) );
  OR2X1 U925 ( .A(n427), .B(n440), .Y(n178) );
  MUX2X1 U926 ( .B(n1225), .A(n1227), .S(n998), .Y(n583) );
  INVX1 U927 ( .A(n168), .Y(n991) );
  OR2X2 U928 ( .A(n992), .B(n993), .Y(n1096) );
  OR2X2 U929 ( .A(n1186), .B(n1187), .Y(n993) );
  AND2X1 U930 ( .A(a[13]), .B(n1255), .Y(n1264) );
  BUFX2 U931 ( .A(a[14]), .Y(n994) );
  INVX1 U932 ( .A(n723), .Y(n995) );
  INVX2 U933 ( .A(n723), .Y(n996) );
  INVX1 U934 ( .A(b[7]), .Y(n1237) );
  BUFX2 U935 ( .A(n170), .Y(n997) );
  INVX1 U936 ( .A(a[9]), .Y(n1253) );
  AND2X1 U937 ( .A(n807), .B(n636), .Y(n1180) );
  AND2X1 U938 ( .A(n849), .B(n1172), .Y(n1176) );
  OR2X2 U939 ( .A(n48), .B(n1221), .Y(n587) );
  XNOR2X1 U940 ( .A(n1256), .B(a[14]), .Y(n998) );
  INVX1 U941 ( .A(n173), .Y(n999) );
  AND2X2 U942 ( .A(n1210), .B(n1178), .Y(n1179) );
  INVX1 U943 ( .A(n636), .Y(n1178) );
  XNOR2X1 U944 ( .A(n1255), .B(a[12]), .Y(n1000) );
  INVX2 U945 ( .A(n1000), .Y(n42) );
  INVX1 U946 ( .A(n1255), .Y(n1254) );
  INVX8 U947 ( .A(n727), .Y(n807) );
  INVX1 U948 ( .A(b[9]), .Y(n1239) );
  INVX1 U949 ( .A(b[10]), .Y(n1241) );
  INVX8 U950 ( .A(a[1]), .Y(n1248) );
  XNOR2X1 U951 ( .A(n114), .B(n1001), .Y(product[31]) );
  XNOR2X1 U952 ( .A(n287), .B(n286), .Y(n1001) );
  BUFX4 U953 ( .A(n30), .Y(n1208) );
  AND2X2 U954 ( .A(n1004), .B(n1022), .Y(n450) );
  INVX1 U955 ( .A(n450), .Y(n1002) );
  INVX1 U956 ( .A(n1175), .Y(n1003) );
  INVX1 U957 ( .A(n1177), .Y(n1004) );
  OR2X2 U958 ( .A(n1105), .B(n999), .Y(n168) );
  INVX1 U959 ( .A(n168), .Y(n1005) );
  OR2X2 U960 ( .A(n1026), .B(n1148), .Y(n146) );
  INVX1 U961 ( .A(n146), .Y(n1006) );
  INVX1 U962 ( .A(n1176), .Y(n1007) );
  AND2X2 U963 ( .A(n1063), .B(n1005), .Y(n166) );
  INVX1 U964 ( .A(n166), .Y(n1008) );
  BUFX2 U965 ( .A(n238), .Y(n1009) );
  BUFX2 U966 ( .A(n230), .Y(n1010) );
  BUFX2 U967 ( .A(n186), .Y(n1011) );
  BUFX2 U968 ( .A(n145), .Y(n1012) );
  AND2X1 U969 ( .A(n420), .B(n422), .Y(n1186) );
  BUFX2 U970 ( .A(n219), .Y(n1013) );
  BUFX2 U971 ( .A(n197), .Y(n1014) );
  INVX1 U972 ( .A(n167), .Y(n1015) );
  INVX1 U973 ( .A(n1015), .Y(n1016) );
  INVX1 U974 ( .A(n121), .Y(n256) );
  INVX1 U975 ( .A(n115), .Y(n255) );
  OR2X1 U976 ( .A(n1102), .B(n1124), .Y(n187) );
  INVX1 U977 ( .A(n187), .Y(n1017) );
  OR2X1 U978 ( .A(n1100), .B(n1123), .Y(n209) );
  INVX1 U979 ( .A(n209), .Y(n1018) );
  AND2X1 U980 ( .A(n1164), .B(n1160), .Y(n196) );
  INVX1 U981 ( .A(n196), .Y(n1019) );
  AND2X1 U982 ( .A(n1159), .B(n1165), .Y(n218) );
  INVX1 U983 ( .A(n218), .Y(n1020) );
  AND2X1 U984 ( .A(n1078), .B(n189), .Y(n100) );
  INVX1 U985 ( .A(n100), .Y(n1021) );
  INVX1 U986 ( .A(n208), .Y(n1023) );
  INVX1 U987 ( .A(n1023), .Y(n1024) );
  BUFX2 U988 ( .A(n152), .Y(n1025) );
  INVX1 U989 ( .A(n151), .Y(n1026) );
  BUFX2 U990 ( .A(n1012), .Y(n1027) );
  INVX1 U991 ( .A(n137), .Y(n1028) );
  INVX1 U992 ( .A(n1028), .Y(n1029) );
  INVX1 U993 ( .A(n1028), .Y(n1030) );
  INVX1 U994 ( .A(n129), .Y(n1031) );
  INVX1 U995 ( .A(n1031), .Y(n1032) );
  INVX1 U996 ( .A(n1031), .Y(n1033) );
  BUFX2 U997 ( .A(n789), .Y(n1034) );
  INVX4 U998 ( .A(n721), .Y(n46) );
  AND2X2 U999 ( .A(a[15]), .B(n1256), .Y(n1265) );
  INVX1 U1000 ( .A(n1265), .Y(n1036) );
  INVX1 U1001 ( .A(n743), .Y(n1037) );
  INVX1 U1002 ( .A(n747), .Y(n1038) );
  INVX1 U1003 ( .A(n748), .Y(n1040) );
  INVX1 U1004 ( .A(n744), .Y(n1041) );
  INVX1 U1005 ( .A(n745), .Y(n1042) );
  INVX1 U1006 ( .A(n746), .Y(n1043) );
  INVX1 U1007 ( .A(n752), .Y(n1044) );
  AND2X2 U1008 ( .A(a[9]), .B(n1252), .Y(n1262) );
  INVX1 U1009 ( .A(n1262), .Y(n1045) );
  INVX1 U1010 ( .A(n96), .Y(n1046) );
  AND2X1 U1011 ( .A(a[3]), .B(n1248), .Y(n1259) );
  INVX1 U1012 ( .A(n1259), .Y(n1048) );
  INVX1 U1013 ( .A(n608), .Y(n1049) );
  BUFX4 U1014 ( .A(n1171), .Y(n1155) );
  INVX1 U1015 ( .A(n98), .Y(n1050) );
  BUFX2 U1016 ( .A(n180), .Y(n1051) );
  INVX1 U1017 ( .A(n97), .Y(n1052) );
  AND2X2 U1018 ( .A(n411), .B(n1189), .Y(n171) );
  INVX1 U1019 ( .A(n171), .Y(n1053) );
  INVX1 U1020 ( .A(n289), .Y(n1054) );
  INVX1 U1021 ( .A(n1261), .Y(n1055) );
  AND2X1 U1022 ( .A(n1075), .B(n1168), .Y(n110) );
  INVX1 U1023 ( .A(n110), .Y(n1056) );
  AND2X1 U1024 ( .A(n1074), .B(n1169), .Y(n112) );
  INVX1 U1025 ( .A(n112), .Y(n1057) );
  AND2X1 U1026 ( .A(n1097), .B(n244), .Y(n111) );
  INVX1 U1027 ( .A(n111), .Y(n1058) );
  AND2X1 U1028 ( .A(n1077), .B(n275), .Y(n104) );
  INVX1 U1029 ( .A(n104), .Y(n1059) );
  AND2X1 U1030 ( .A(n1098), .B(n143), .Y(n92) );
  INVX1 U1031 ( .A(n92), .Y(n1060) );
  INVX1 U1032 ( .A(n156), .Y(n1061) );
  AND2X2 U1033 ( .A(n440), .B(n427), .Y(n179) );
  INVX1 U1034 ( .A(n179), .Y(n1062) );
  OR2X2 U1035 ( .A(n1104), .B(n1116), .Y(n176) );
  INVX1 U1036 ( .A(n176), .Y(n1063) );
  INVX1 U1037 ( .A(n331), .Y(n1064) );
  AND2X1 U1038 ( .A(b[15]), .B(n1217), .Y(n570) );
  INVX1 U1039 ( .A(n570), .Y(n1065) );
  AND2X1 U1040 ( .A(n1093), .B(n1167), .Y(n108) );
  INVX1 U1041 ( .A(n108), .Y(n1066) );
  INVX1 U1042 ( .A(n94), .Y(n1067) );
  OR2X2 U1043 ( .A(n368), .B(n381), .Y(n1158) );
  INVX1 U1044 ( .A(n106), .Y(n1068) );
  BUFX2 U1045 ( .A(n224), .Y(n1069) );
  INVX1 U1046 ( .A(n102), .Y(n1070) );
  BUFX2 U1047 ( .A(n202), .Y(n1071) );
  AND2X1 U1048 ( .A(n1118), .B(n127), .Y(n88) );
  INVX1 U1049 ( .A(n88), .Y(n1072) );
  AND2X1 U1050 ( .A(n334), .B(n343), .Y(n141) );
  INVX1 U1051 ( .A(n141), .Y(n1073) );
  AND2X1 U1052 ( .A(n878), .B(n551), .Y(n250) );
  INVX1 U1053 ( .A(n250), .Y(n1074) );
  AND2X1 U1054 ( .A(n548), .B(n545), .Y(n242) );
  INVX1 U1055 ( .A(n242), .Y(n1075) );
  INVX1 U1056 ( .A(n149), .Y(n1076) );
  INVX1 U1057 ( .A(n212), .Y(n1077) );
  INVX1 U1058 ( .A(n190), .Y(n1078) );
  INVX1 U1059 ( .A(n750), .Y(n1079) );
  BUFX2 U1060 ( .A(n175), .Y(n1080) );
  INVX1 U1061 ( .A(n353), .Y(n1081) );
  INVX1 U1062 ( .A(n1263), .Y(n1082) );
  INVX1 U1063 ( .A(n627), .Y(n1083) );
  INVX1 U1064 ( .A(n589), .Y(n1084) );
  AND2X1 U1065 ( .A(n1117), .B(n236), .Y(n109) );
  INVX1 U1066 ( .A(n109), .Y(n1085) );
  AND2X1 U1067 ( .A(n1149), .B(n214), .Y(n105) );
  INVX1 U1068 ( .A(n105), .Y(n1086) );
  INVX1 U1069 ( .A(n99), .Y(n1087) );
  INVX1 U1070 ( .A(n101), .Y(n1088) );
  INVX1 U1071 ( .A(n95), .Y(n1089) );
  AND2X1 U1072 ( .A(n1119), .B(n135), .Y(n90) );
  INVX1 U1073 ( .A(n90), .Y(n1090) );
  AND2X1 U1074 ( .A(n302), .B(n307), .Y(n125) );
  INVX1 U1075 ( .A(n125), .Y(n1091) );
  AND2X1 U1076 ( .A(n316), .B(n323), .Y(n133) );
  INVX1 U1077 ( .A(n133), .Y(n1092) );
  AND2X1 U1078 ( .A(n540), .B(n535), .Y(n234) );
  INVX1 U1079 ( .A(n234), .Y(n1093) );
  INVX1 U1080 ( .A(n223), .Y(n1094) );
  INVX1 U1081 ( .A(n201), .Y(n1095) );
  AND2X2 U1082 ( .A(n420), .B(n434), .Y(n1187) );
  AND2X1 U1083 ( .A(n550), .B(n549), .Y(n245) );
  INVX1 U1084 ( .A(n245), .Y(n1097) );
  AND2X1 U1085 ( .A(n355), .B(n344), .Y(n144) );
  INVX1 U1086 ( .A(n144), .Y(n1098) );
  OR2X1 U1087 ( .A(n1153), .B(n252), .Y(n251) );
  INVX1 U1088 ( .A(n251), .Y(n1099) );
  INVX1 U1089 ( .A(n211), .Y(n1100) );
  INVX1 U1090 ( .A(n211), .Y(n1101) );
  INVX1 U1091 ( .A(n189), .Y(n1102) );
  INVX1 U1092 ( .A(n178), .Y(n1103) );
  INVX1 U1093 ( .A(n178), .Y(n1104) );
  OR2X2 U1094 ( .A(n411), .B(n396), .Y(n170) );
  INVX1 U1095 ( .A(n170), .Y(n1105) );
  INVX1 U1096 ( .A(n997), .Y(n1106) );
  INVX1 U1097 ( .A(n379), .Y(n1107) );
  AND2X1 U1098 ( .A(n807), .B(n635), .Y(n1192) );
  INVX1 U1099 ( .A(n1192), .Y(n1108) );
  AND2X1 U1100 ( .A(n1210), .B(n1190), .Y(n1191) );
  INVX1 U1101 ( .A(n1191), .Y(n1109) );
  AND2X1 U1102 ( .A(n1153), .B(n1170), .Y(product[0]) );
  INVX1 U1103 ( .A(n646), .Y(n1110) );
  AND2X1 U1104 ( .A(b[15]), .B(n1247), .Y(n703) );
  INVX1 U1105 ( .A(n703), .Y(n1111) );
  INVX1 U1106 ( .A(n107), .Y(n1112) );
  INVX1 U1107 ( .A(n103), .Y(n1113) );
  AND2X1 U1108 ( .A(n1139), .B(n1166), .Y(n86) );
  INVX1 U1109 ( .A(n86), .Y(n1114) );
  INVX1 U1110 ( .A(n93), .Y(n1115) );
  OR2X2 U1111 ( .A(n441), .B(n454), .Y(n183) );
  INVX1 U1112 ( .A(n183), .Y(n1116) );
  AND2X1 U1113 ( .A(n544), .B(n541), .Y(n237) );
  INVX1 U1114 ( .A(n237), .Y(n1117) );
  AND2X1 U1115 ( .A(n308), .B(n315), .Y(n128) );
  INVX1 U1116 ( .A(n128), .Y(n1118) );
  AND2X1 U1117 ( .A(n324), .B(n333), .Y(n136) );
  INVX1 U1118 ( .A(n136), .Y(n1119) );
  OR2X1 U1119 ( .A(n344), .B(n355), .Y(n143) );
  INVX1 U1120 ( .A(n143), .Y(n1120) );
  INVX1 U1121 ( .A(n158), .Y(n1121) );
  BUFX2 U1122 ( .A(n246), .Y(n1122) );
  INVX1 U1123 ( .A(n214), .Y(n1123) );
  INVX1 U1124 ( .A(n192), .Y(n1124) );
  OR2X2 U1125 ( .A(n412), .B(n426), .Y(n173) );
  INVX1 U1126 ( .A(n173), .Y(n1125) );
  INVX1 U1127 ( .A(n299), .Y(n1126) );
  INVX1 U1128 ( .A(n1264), .Y(n1127) );
  INVX1 U1129 ( .A(n1260), .Y(n1128) );
  INVX1 U1130 ( .A(n1182), .Y(n1129) );
  INVX1 U1131 ( .A(n1183), .Y(n1130) );
  INVX1 U1132 ( .A(n1180), .Y(n1131) );
  INVX1 U1133 ( .A(n1179), .Y(n1132) );
  AND2X2 U1134 ( .A(n1132), .B(n1131), .Y(n1172) );
  AND2X1 U1135 ( .A(b[15]), .B(n1201), .Y(n665) );
  INVX1 U1136 ( .A(n665), .Y(n1133) );
  AND2X1 U1137 ( .A(b[15]), .B(n1197), .Y(n684) );
  INVX1 U1138 ( .A(n684), .Y(n1134) );
  INVX1 U1139 ( .A(n87), .Y(n1135) );
  INVX1 U1140 ( .A(n91), .Y(n1136) );
  INVX1 U1141 ( .A(n89), .Y(n1137) );
  INVX1 U1142 ( .A(n2), .Y(n1138) );
  AND2X1 U1143 ( .A(n292), .B(n295), .Y(n119) );
  INVX1 U1144 ( .A(n119), .Y(n1139) );
  INVX1 U1145 ( .A(n228), .Y(n1140) );
  INVX1 U1146 ( .A(n206), .Y(n1141) );
  OR2X1 U1147 ( .A(n549), .B(n550), .Y(n244) );
  INVX1 U1148 ( .A(n244), .Y(n1142) );
  OR2X1 U1149 ( .A(n541), .B(n544), .Y(n236) );
  INVX1 U1150 ( .A(n236), .Y(n1143) );
  OR2X1 U1151 ( .A(n315), .B(n308), .Y(n127) );
  INVX1 U1152 ( .A(n127), .Y(n1144) );
  OR2X1 U1153 ( .A(n333), .B(n324), .Y(n135) );
  INVX1 U1154 ( .A(n135), .Y(n1145) );
  INVX1 U1155 ( .A(n159), .Y(n1146) );
  INVX1 U1156 ( .A(n184), .Y(n1147) );
  OR2X1 U1157 ( .A(n356), .B(n367), .Y(n148) );
  INVX1 U1158 ( .A(n148), .Y(n1148) );
  AND2X1 U1159 ( .A(n520), .B(n513), .Y(n215) );
  INVX1 U1160 ( .A(n215), .Y(n1149) );
  AND2X1 U1161 ( .A(n480), .B(n469), .Y(n193) );
  INVX1 U1162 ( .A(n193), .Y(n1150) );
  AND2X2 U1163 ( .A(n426), .B(n412), .Y(n174) );
  INVX1 U1164 ( .A(n174), .Y(n1151) );
  OR2X1 U1165 ( .A(n557), .B(n1258), .Y(n313) );
  INVX1 U1166 ( .A(n313), .Y(n1152) );
  AND2X1 U1167 ( .A(n742), .B(n895), .Y(n254) );
  INVX1 U1168 ( .A(n254), .Y(n1153) );
  BUFX2 U1169 ( .A(n142), .Y(n1154) );
  BUFX2 U1170 ( .A(n126), .Y(n1156) );
  BUFX2 U1171 ( .A(n134), .Y(n1157) );
  INVX1 U1172 ( .A(n1224), .Y(n1222) );
  INVX2 U1173 ( .A(n729), .Y(n825) );
  BUFX2 U1174 ( .A(n42), .Y(n1214) );
  INVX1 U1175 ( .A(n1221), .Y(n1220) );
  INVX1 U1176 ( .A(n217), .Y(n216) );
  INVX1 U1177 ( .A(n1024), .Y(n207) );
  INVX1 U1178 ( .A(n1010), .Y(n229) );
  INVX1 U1179 ( .A(n1101), .Y(n275) );
  OR2X1 U1180 ( .A(n343), .B(n334), .Y(n1161) );
  OR2X1 U1181 ( .A(n307), .B(n302), .Y(n1162) );
  OR2X1 U1182 ( .A(n323), .B(n316), .Y(n1163) );
  BUFX2 U1183 ( .A(n24), .Y(n1205) );
  BUFX2 U1184 ( .A(n24), .Y(n1204) );
  BUFX2 U1185 ( .A(n12), .Y(n1196) );
  BUFX2 U1186 ( .A(n1214), .Y(n1173) );
  BUFX2 U1187 ( .A(n44), .Y(n1218) );
  BUFX2 U1188 ( .A(n20), .Y(n1206) );
  BUFX2 U1189 ( .A(n8), .Y(n1198) );
  BUFX2 U1190 ( .A(n44), .Y(n1219) );
  BUFX2 U1191 ( .A(n20), .Y(n1207) );
  BUFX2 U1192 ( .A(n8), .Y(n1199) );
  INVX1 U1193 ( .A(n1228), .Y(n1227) );
  INVX1 U1194 ( .A(n1226), .Y(n1225) );
  OR2X1 U1195 ( .A(n295), .B(n292), .Y(n1166) );
  OR2X1 U1196 ( .A(n535), .B(n540), .Y(n1167) );
  OR2X1 U1197 ( .A(n545), .B(n548), .Y(n1168) );
  BUFX2 U1198 ( .A(n18), .Y(n1201) );
  BUFX2 U1199 ( .A(n18), .Y(n1200) );
  INVX1 U1200 ( .A(b[3]), .Y(n1228) );
  BUFX2 U1201 ( .A(n14), .Y(n1202) );
  BUFX2 U1202 ( .A(n38), .Y(n1215) );
  BUFX2 U1203 ( .A(n1138), .Y(n1194) );
  BUFX2 U1204 ( .A(n32), .Y(n1213) );
  BUFX2 U1205 ( .A(n14), .Y(n1203) );
  BUFX2 U1206 ( .A(n38), .Y(n1216) );
  BUFX2 U1207 ( .A(n32), .Y(n1212) );
  BUFX2 U1208 ( .A(n1138), .Y(n1195) );
  INVX1 U1209 ( .A(n1230), .Y(n1229) );
  INVX1 U1210 ( .A(n894), .Y(n252) );
  INVX1 U1211 ( .A(b[2]), .Y(n1226) );
  INVX1 U1212 ( .A(n1251), .Y(n1250) );
  OR2X1 U1213 ( .A(n551), .B(n878), .Y(n1169) );
  INVX1 U1214 ( .A(n1224), .Y(n1223) );
  INVX1 U1215 ( .A(n1245), .Y(n1244) );
  OR2X1 U1216 ( .A(n895), .B(n742), .Y(n1170) );
  XOR2X1 U1217 ( .A(n1253), .B(a[10]), .Y(n1171) );
  AND2X1 U1218 ( .A(n1211), .B(n727), .Y(n738) );
  BUFX2 U1219 ( .A(n26), .Y(n1211) );
  BUFX2 U1220 ( .A(n26), .Y(n1210) );
  INVX1 U1221 ( .A(b[1]), .Y(n1224) );
  INVX1 U1222 ( .A(b[4]), .Y(n1230) );
  INVX1 U1223 ( .A(b[6]), .Y(n1234) );
  INVX1 U1224 ( .A(a[3]), .Y(n1249) );
  INVX1 U1225 ( .A(n1232), .Y(n1231) );
  INVX1 U1226 ( .A(n1237), .Y(n1236) );
  INVX1 U1227 ( .A(b[0]), .Y(n1221) );
  INVX1 U1228 ( .A(b[12]), .Y(n1243) );
  INVX1 U1229 ( .A(b[5]), .Y(n1232) );
  INVX1 U1230 ( .A(a[0]), .Y(n1247) );
  INVX1 U1231 ( .A(a[0]), .Y(n1246) );
  INVX1 U1232 ( .A(n990), .Y(n164) );
  XOR2X1 U1233 ( .A(n865), .B(n849), .Y(n1174) );
  XOR2X1 U1234 ( .A(n1172), .B(n1174), .Y(n451) );
  INVX1 U1235 ( .A(n617), .Y(n1181) );
  XOR2X1 U1236 ( .A(n420), .B(n434), .Y(n1185) );
  XOR2X1 U1237 ( .A(n422), .B(n1185), .Y(n416) );
  INVX1 U1238 ( .A(n1103), .Y(n269) );
  INVX1 U1239 ( .A(n1011), .Y(n185) );
  INVX1 U1240 ( .A(n195), .Y(n194) );
  INVX1 U1241 ( .A(n396), .Y(n1188) );
  INVX1 U1242 ( .A(n1188), .Y(n1189) );
  INVX1 U1243 ( .A(n635), .Y(n1190) );
  INVX1 U1244 ( .A(n1125), .Y(n268) );
  OAI21X1 U1245 ( .A(a[2]), .B(n1249), .C(n1048), .Y(n733) );
  OAI21X1 U1246 ( .A(a[4]), .B(n1251), .C(n1128), .Y(n731) );
  OAI21X1 U1247 ( .A(a[6]), .B(n1252), .C(n1055), .Y(n729) );
  OAI21X1 U1248 ( .A(a[8]), .B(n1253), .C(n1045), .Y(n727) );
  OAI21X1 U1249 ( .A(a[10]), .B(n1255), .C(n1082), .Y(n725) );
  OAI21X1 U1250 ( .A(a[12]), .B(n1256), .C(n1127), .Y(n723) );
  OAI21X1 U1251 ( .A(n994), .B(n1258), .C(n1036), .Y(n721) );
  XOR2X1 U1252 ( .A(n46), .B(n1037), .Y(n285) );
endmodule


module alu ( clk, oprA, oprB, shift_amount, op, ww, result, mult32_result );
  input [0:63] oprA;
  input [0:63] oprB;
  input [0:4] shift_amount;
  input [0:5] op;
  input [0:1] ww;
  output [0:63] result;
  output [0:63] mult32_result;
  input clk;
  wire   n10612, n10613, n10614, n10615, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1516, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1741, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n7984, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n87, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1517, n1533,
         n1549, n1565, n1581, n1613, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1742, n1758, n1774, n1790, n1806, n1838, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12;
  wire   [0:31] mult32_A;
  wire   [0:31] mult32_B;

  alu_DW02_mult_2_stage_0 ALU_MUL32 ( .A({mult32_A[0:11], n5575, 
        mult32_A[13:14], n5645, mult32_A[16:26], n5028, n5049, mult32_A[29:30], 
        n5510}), .B({n175, n5306, n5453, n5658, n5591, n5454, n5659, n5401, 
        n5521, n5657, n5660, n5590, n5592, n5661, n5593, n5456, n5457, n5663, 
        n5403, n5402, n5404, n5664, n5522, n5405, n5459, n5523, n5458, n5455, 
        n5662, n5665, n5460, n174}), .TC(1'b0), .CLK(clk), .PRODUCT(
        mult32_result) );
  alu_DW_rightsh_0 sra_516 ( .A({n6061, n6058, n6057, n6054, n6051, n21, n5734, 
        n6042, n6039, n5277, n6034, n5885, n6032, n6342, n6026, n59, n5271, 
        n6022, n6018, n6016, n5269, n6332, n5270, n6328, n5274, n6322, n6319, 
        n43, n5276, n5995, n5993, n5991, n5989, n5987, n5984, n5981, n6303, 
        n6301, n5976, n5973, n5970, n6296, n5966, n5964, n5960, n5958, n5953, 
        n5952, n5949, n6290, n5944, n5942, n5940, n5938, n5934, n5932, n5929, 
        n5927, n5925, n66, n5922, n5918, n5915, n5911}), .DATA_TC(1'b1), .SH({
        shift_amount[0], n6156, n5890, shift_amount[3], n5888}), .B({n3898, 
        n3897, n3896, n3895, n3894, n3893, n3892, n3891, n3890, n3889, n3888, 
        n3887, n3886, n3885, n3884, n3883, n3882, n3881, n3880, n3879, n3878, 
        n3877, n3876, n3875, n3874, n3873, n3872, n3871, n3870, n3869, n3868, 
        n3867, n3866, n3865, n3864, n3863, n3862, n3861, n3860, n3859, n3858, 
        n3857, n3856, n3855, n3854, n3853, n3852, n3851, n3850, n3849, n3848, 
        n3847, n3846, n3845, n3844, n3843, n3842, n3841, n3840, n3839, n3838, 
        n3837, n3836, n3835}) );
  alu_DW_rightsh_1 sra_512 ( .A({n5988, n6308, n5984, n5981, n6303, n5978, 
        n5975, n5974, n5970, n6296, n45, n5965, n5961, n5958, n5953, n5952, 
        n5948, n5947, n5944, n5942, n5940, n5937, n5933, n5931, n5929, n5926, 
        n5924, n66, n17, n5918, n5916, n5912}), .DATA_TC(1'b1), .SH({
        shift_amount[0], n6156, n5889, shift_amount[3], n5887}), .B({n3834, 
        n3833, n3832, n3831, n3830, n3829, n3828, n3827, n3826, n3825, n3824, 
        n3823, n3822, n3821, n3820, n3819, n3818, n3817, n3816, n3815, n3814, 
        n3813, n3812, n3811, n3810, n3809, n3808, n3807, n3806, n3805, n3804, 
        n3803}) );
  alu_DW_rightsh_2 sra_511 ( .A({n6060, n6059, n6057, n6055, n6052, n6049, 
        n6046, n6042, n6039, n6037, n6034, n5885, n6032, n6029, n6026, n59, 
        n5272, n5282, n6018, n5286, n5269, n6008, n10, n6004, n6003, n6322, 
        n6319, n43, n5276, n6315, n5992, n5880}), .DATA_TC(1'b1), .SH({
        shift_amount[0], n6156, n5890, shift_amount[3], n5888}), .B({n3802, 
        n3801, n3800, n3799, n3798, n3797, n3796, n3795, n3794, n3793, n3792, 
        n3791, n3790, n3789, n3788, n3787, n3786, n3785, n3784, n3783, n3782, 
        n3781, n3780, n3779, n3778, n3777, n3776, n3775, n3774, n3773, n3772, 
        n3771}) );
  alu_DW_rightsh_15 sra_482 ( .A({n6061, n6058, n6057, n6054, n6052, n6049, 
        n5734, n6042, n6039, n6038, n6034, n5885, n6032, n6342, n6026, n59, 
        n5271, n6022, n6018, n6016, n5285, n6008, n6330, n6328, n5274, n6322, 
        n6319, n27, n5276, n6315, n5993, n5879, n5989, n5986, n5983, n5981, 
        n5980, n5977, n5975, n5973, n5970, n5969, n45, n5965, n5961, n5958, 
        n5955, n5952, n5948, n6290, n5945, n5942, n5941, n5938, n5934, n5932, 
        n5929, n5927, n5925, n66, n5922, n5918, n5916, n5911}), .DATA_TC(1'b1), 
        .SH({n6163, n5904, n5901, n5899, n5895, n5892}), .B({n3577, n3576, 
        n3575, n3574, n3573, n3572, n3571, n3570, n3569, n3568, n3567, n3566, 
        n3565, n3564, n3563, n3562, n3561, n3560, n3559, n3558, n3557, n3556, 
        n3555, n3554, n3553, n3552, n3551, n3550, n3549, n3548, n3547, n3546, 
        n3545, n3544, n3543, n3542, n3541, n3540, n3539, n3538, n3537, n3536, 
        n3535, n3534, n3533, n3532, n3531, n3530, n3529, n3528, n3527, n3526, 
        n3525, n3524, n3523, n3522, n3521, n3520, n3519, n3518, n3517, n3516, 
        n3515, n3514}) );
  alu_DW_rightsh_16 sra_478 ( .A({n5989, n6308, n5984, n5982, n5980, n5977, 
        n5976, n5974, n5970, n5969, n5966, n5964, n5960, n5958, n5955, n5952, 
        n5949, n6290, n5945, n6288, n5940, n5938, n5933, n5931, n5929, n5926, 
        n5924, n66, n17, n5918, n5915, n5912}), .DATA_TC(1'b1), .SH({n5906, 
        n5902, n5900, n5897, n8}), .B({n3513, n3512, n3511, n3510, n3509, 
        n3508, n3507, n3506, n3505, n3504, n3503, n3502, n3501, n3500, n3499, 
        n3498, n3497, n3496, n3495, n3494, n3493, n3492, n3491, n3490, n3489, 
        n3488, n3487, n3486, n3485, n3484, n3483, n3482}) );
  alu_DW_rightsh_17 sra_477 ( .A({n6061, n6059, n6057, n6054, n6051, n21, 
        n5734, n6043, n6039, n6037, n6034, n5885, n6032, n6029, n6026, n59, 
        n5271, n5282, n6018, n6016, n5269, n6008, n10, n6004, n6003, n5283, 
        n6000, n44, n5276, n5995, n5992, n5991}), .DATA_TC(1'b1), .SH({n6222, 
        n5882, n5908, n6217, n5267}), .B({n3481, n3480, n3479, n3478, n3477, 
        n3476, n3475, n3474, n3473, n3472, n3471, n3470, n3469, n3468, n3467, 
        n3466, n3465, n3464, n3463, n3462, n3461, n3460, n3459, n3458, n3457, 
        n3456, n3455, n3454, n3453, n3452, n3451, n3450}) );
  alu_DW_rightsh_30 srl_448 ( .A({n6060, n6058, n6057, n6054, n6052, n21, 
        n5734, n6043, n6039, n5277, n6034, n5885, n6032, n6029, n6026, n59, 
        n5271, n6022, n6018, n5286, n5285, n6008, n6007, n6328, n5274, n5283, 
        n6319, n27, n5276, n6315, n5992, n5991, n5988, n5987, n5984, n5982, 
        n5980, n5978, n5975, n5973, n6297, n5968, n5966, n5965, n5961, n5958, 
        n5953, n5952, n5949, n6290, n5944, n5942, n5941, n5937, n5933, n5931, 
        n5929, n5926, n5924, n67, n5922, n5918, n5915, n5911}), .DATA_TC(1'b0), 
        .SH({shift_amount[0], n6156, n5890, shift_amount[3], n5886}), .B({
        n3256, n3255, n3254, n3253, n3252, n3251, n3250, n3249, n3248, n3247, 
        n3246, n3245, n3244, n3243, n3242, n3241, n3240, n3239, n3238, n3237, 
        n3236, n3235, n3234, n3233, n3232, n3231, n3230, n3229, n3228, n3227, 
        n3226, n3225, n3224, n3223, n3222, n3221, n3220, n3219, n3218, n3217, 
        n3216, n3215, n3214, n3213, n3212, n3211, n3210, n3209, n3208, n3207, 
        n3206, n3205, n3204, n3203, n3202, n3201, n3200, n3199, n3198, n3197, 
        n3196, n3195, n3194, n3193}) );
  alu_DW_rightsh_31 srl_444 ( .A({n5988, n5986, n5985, n5982, n6303, n6301, 
        n5975, n5974, n6297, n5968, n5966, n5964, n5960, n5957, n5953, n5952, 
        n5948, n6290, n5945, n6288, n5941, n5937, n5934, n5932, n5929, n5927, 
        n5924, n66, n6275, n5918, n5916, n5912}), .DATA_TC(1'b0), .SH({
        shift_amount[0], n6156, n6154, shift_amount[3], n5886}), .B({n3192, 
        n3191, n3190, n3189, n3188, n3187, n3186, n3185, n3184, n3183, n3182, 
        n3181, n3180, n3179, n3178, n3177, n3176, n3175, n3174, n3173, n3172, 
        n3171, n3170, n3169, n3168, n3167, n3166, n3165, n3164, n3163, n3162, 
        n3161}) );
  alu_DW_rightsh_32 srl_443 ( .A({n6061, n6058, n6057, n6054, n6052, n21, 
        n5734, n6042, n6039, n6037, n6034, n5885, n6032, n6029, n6026, n59, 
        n5272, n5282, n6018, n5286, n5269, n6332, n10, n6004, n5274, n6322, 
        n6319, n44, n5276, n6315, n5993, n5879}), .DATA_TC(1'b0), .SH({
        shift_amount[0], n6156, n5890, shift_amount[3], n5888}), .B({n3160, 
        n3159, n3158, n3157, n3156, n3155, n3154, n3153, n3152, n3151, n3150, 
        n3149, n3148, n3147, n3146, n3145, n3144, n3143, n3142, n3141, n3140, 
        n3139, n3138, n3137, n3136, n3135, n3134, n3133, n3132, n3131, n3130, 
        n3129}) );
  alu_DW_rightsh_45 srl_414 ( .A({n6060, n6059, n6354, n6055, n6052, n6049, 
        n6046, n6043, n6039, n6038, n6034, n5885, n6032, n6342, n6026, n59, 
        n5271, n6022, n6018, n6016, n5285, n6332, n6007, n6328, n6003, n5283, 
        n5268, n44, n5276, n6315, n5993, n5879, n5988, n6308, n5984, n5981, 
        n5980, n5978, n5976, n5974, n5970, n6296, n45, n5965, n5961, n5957, 
        n5955, n5952, n5949, n5947, n5944, n5942, n5940, n5937, n5934, n5932, 
        n5929, n5926, n5925, n67, n17, n5918, n5916, n5912}), .DATA_TC(1'b0), 
        .SH({n6163, n5905, n5903, n5900, n5895, n5892}), .B({n2935, n2934, 
        n2933, n2932, n2931, n2930, n2929, n2928, n2927, n2926, n2925, n2924, 
        n2923, n2922, n2921, n2920, n2919, n2918, n2917, n2916, n2915, n2914, 
        n2913, n2912, n2911, n2910, n2909, n2908, n2907, n2906, n2905, n2904, 
        n2903, n2902, n2901, n2900, n2899, n2898, n2897, n2896, n2895, n2894, 
        n2893, n2892, n2891, n2890, n2889, n2888, n2887, n2886, n2885, n2884, 
        n2883, n2882, n2881, n2880, n2879, n2878, n2877, n2876, n2875, n2874, 
        n2873, n2872}) );
  alu_DW_rightsh_46 srl_410 ( .A({n5989, n5986, n5984, n5981, n5980, n5977, 
        n5976, n5973, n6297, n5969, n5966, n5964, n5960, n5958, n5955, n5952, 
        n5948, n6290, n5945, n6288, n5940, n5937, n5934, n5932, n5929, n5927, 
        n5924, n66, n5922, n5918, n5916, n5912}), .DATA_TC(1'b0), .SH({n5906, 
        n5901, n5899, n5896, n5892}), .B({n2871, n2870, n2869, n2868, n2867, 
        n2866, n2865, n2864, n2863, n2862, n2861, n2860, n2859, n2858, n2857, 
        n2856, n2855, n2854, n2853, n2852, n2851, n2850, n2849, n2848, n2847, 
        n2846, n2845, n2844, n2843, n2842, n2841, n2840}) );
  alu_DW_rightsh_47 srl_409 ( .A({n6061, n6058, n6057, n6055, n6052, n6049, 
        n6046, n6042, n6039, n6037, n6034, n5885, n6032, n6342, n6026, n59, 
        n5272, n5282, n6018, n5286, n5269, n6008, n10, n6004, n5274, n6322, 
        n6319, n44, n5276, n6315, n5992, n5991}), .DATA_TC(1'b0), .SH({n6222, 
        n6220, n5907, n6217, n5267}), .B({n2839, n2838, n2837, n2836, n2835, 
        n2834, n2833, n2832, n2831, n2830, n2829, n2828, n2827, n2826, n2825, 
        n2824, n2823, n2822, n2821, n2820, n2819, n2818, n2817, n2816, n2815, 
        n2814, n2813, n2812, n2811, n2810, n2809, n2808}) );
  alu_DW_leftsh_0 sll_380 ( .A({n6061, n6059, n6057, n6055, n6051, n21, n5734, 
        n6043, n6039, n6037, n6034, n5885, n6032, n6029, n6026, n59, n5271, 
        n6022, n6018, n6016, n5285, n6008, n6007, n6328, n6003, n5283, n6000, 
        n27, n5276, n5995, n5993, n5991, n5989, n5987, n5984, n5981, n5980, 
        n6301, n5976, n5974, n5970, n5968, n45, n5965, n5961, n5957, n5953, 
        n5952, n5949, n6290, n5944, n5942, n5941, n5938, n5933, n5931, n5929, 
        n5926, n5925, n67, n6275, n5918, n5915, n5912}), .SH({shift_amount[0], 
        n6156, n6154, shift_amount[3], n5887}), .B({n2614, n2613, n2612, n2611, 
        n2610, n2609, n2608, n2607, n2606, n2605, n2604, n2603, n2602, n2601, 
        n2600, n2599, n2598, n2597, n2596, n2595, n2594, n2593, n2592, n2591, 
        n2590, n2589, n2588, n2587, n2586, n2585, n2584, n2583, n2582, n2581, 
        n2580, n2579, n2578, n2577, n2576, n2575, n2574, n2573, n2572, n2571, 
        n2570, n2569, n2568, n2567, n2566, n2565, n2564, n2563, n2562, n2561, 
        n2560, n2559, n2558, n2557, n2556, n2555, n2554, n2553, n2552, n2551})
         );
  alu_DW_leftsh_1 sll_376 ( .A({n5988, n6308, n5983, n5982, n5980, n5977, 
        n5975, n5973, n5970, n5969, n45, n5964, n5960, n5957, n5955, n5951, 
        n5948, n6290, n5945, n5942, n5940, n5938, n5933, n5931, n6282, n5926, 
        n5925, n67, n17, n5918, n5915, n5911}), .SH({shift_amount[0], n6156, 
        n5889, shift_amount[3], n5886}), .B({n2550, n2549, n2548, n2547, n2546, 
        n2545, n2544, n2543, n2542, n2541, n2540, n2539, n2538, n2537, n2536, 
        n2535, n2534, n2533, n2532, n2531, n2530, n2529, n2528, n2527, n2526, 
        n2525, n2524, n2523, n2522, n2521, n2520, n2519}) );
  alu_DW_leftsh_2 sll_375 ( .A({n6060, n6059, n6354, n6054, n6051, n6049, 
        n6046, n6042, n6039, n6037, n6034, n5885, n6032, n6029, n6026, n59, 
        n5272, n5282, n6018, n5286, n5269, n6332, n10, n6004, n5274, n5283, 
        n5268, n27, n5276, n6315, n5992, n5991}), .SH({shift_amount[0], n6156, 
        n5889, shift_amount[3], n5887}), .B({n2518, n2517, n2516, n2515, n2514, 
        n2513, n2512, n2511, n2510, n2509, n2508, n2507, n2506, n2505, n2504, 
        n2503, n2502, n2501, n2500, n2499, n2498, n2497, n2496, n2495, n2494, 
        n2493, n2492, n2491, n2490, n2489, n2488, n2487}) );
  alu_DW_leftsh_15 sll_346 ( .A({n6061, n6356, n6057, n6054, n6052, n21, n5734, 
        n6042, n6039, n6037, n6034, n5885, n6032, n6029, n6026, n59, n5271, 
        n6022, n6018, n6016, n5285, n6332, n6007, n6328, n6003, n6322, n6319, 
        n27, n5276, n5995, n5992, n5880, n5988, n5987, n5983, n5981, n6303, 
        n5978, n5976, n5974, n5970, n6296, n5966, n5965, n5961, n5957, n5955, 
        n5952, n5949, n5947, n5944, n5942, n5941, n5937, n5933, n5931, n5929, 
        n5927, n5924, n66, n5922, n5918, n5916, n5912}), .SH({n6163, n5906, 
        n5902, n5899, n5897, n9}), .B({n2293, n2292, n2291, n2290, n2289, 
        n2288, n2287, n2286, n2285, n2284, n2283, n2282, n2281, n2280, n2279, 
        n2278, n2277, n2276, n2275, n2274, n2273, n2272, n2271, n2270, n2269, 
        n2268, n2267, n2266, n2265, n2264, n2263, n2262, n2261, n2260, n2259, 
        n2258, n2257, n2256, n2255, n2254, n2253, n2252, n2251, n2250, n2249, 
        n2248, n2247, n2246, n2245, n2244, n2243, n2242, n2241, n2240, n2239, 
        n2238, n2237, n2236, n2235, n2234, n2233, n2232, n2231, n2230}) );
  alu_DW_leftsh_16 sll_342 ( .A({n5989, n5986, n5983, n5981, n5980, n6301, 
        n5976, n5973, n6297, n5968, n45, n5964, n5960, n5957, n5953, n5951, 
        n5948, n5947, n5945, n6288, n5941, n5937, n5934, n5932, n5929, n5927, 
        n5925, n66, n6275, n5918, n5916, n5911}), .SH({n5906, n5901, n5899, 
        n5897, n5892}), .B({n2229, n2228, n2227, n2226, n2225, n2224, n2223, 
        n2222, n2221, n2220, n2219, n2218, n2217, n2216, n2215, n2214, n2213, 
        n2212, n2211, n2210, n2209, n2208, n2207, n2206, n2205, n2204, n2203, 
        n2202, n2201, n2200, n2199, n2198}) );
  alu_DW_leftsh_17 sll_341 ( .A({n6061, n6058, n6057, n6054, n6052, n6049, 
        n6046, n6043, n6039, n6037, n6034, n5885, n6032, n6029, n6026, n59, 
        n5271, n5282, n6018, n5286, n5269, n6332, n10, n6004, n5274, n6322, 
        n5268, n43, n5276, n6315, n5993, n5880}), .SH({n6222, n5883, n5907, 
        n6217, n5267}), .B({n2197, n2196, n2195, n2194, n2193, n2192, n2191, 
        n2190, n2189, n2188, n2187, n2186, n2185, n2184, n2183, n2182, n2181, 
        n2180, n2179, n2178, n2177, n2176, n2175, n2174, n2173, n2172, n2171, 
        n2170, n2169, n2168, n2167, n2166}) );
  alu_DW01_sub_7 sub_158 ( .A({n5929, n5926, n6277, n67, n5922, n6273, n5915, 
        n5911}), .B({n6167, n6165, n6163, n5906, n5903, n5899, n5896, n9}), 
        .CI(1'b0), .DIFF({n744, n743, n742, n741, n740, n739, n738, n737}), 
        .CO() );
  alu_DW01_sub_8 sub_157 ( .A({n5948, n6290, n5944, n5942, n5941, n5937, n5934, 
        n5932}), .B({n6183, n6181, n6179, n6177, n6175, n6173, n6171, n6169}), 
        .CI(1'b0), .DIFF({n736, n735, n734, n733, n732, n731, n730, n729}), 
        .CO() );
  alu_DW01_sub_9 sub_156 ( .A({n6297, n5968, n5966, n5963, n5960, n5958, n5953, 
        n5952}), .B({n6199, n6197, n6195, n6193, n6191, n6189, n6187, n6185}), 
        .CI(1'b0), .DIFF({n728, n727, n726, n725, n724, n723, n722, n721}), 
        .CO() );
  alu_DW01_sub_10 sub_155 ( .A({n5988, n5986, n5983, n5982, n5980, n5977, 
        n5975, n5973}), .B({n6215, n6213, n6211, n6209, n6207, n6205, n6203, 
        n6201}), .CI(1'b0), .DIFF({n720, n719, n718, n717, n716, n715, n714, 
        n713}), .CO() );
  alu_DW01_sub_11 sub_154 ( .A({n6325, n58, n5268, n5997, n5276, n6315, n5993, 
        n5991}), .B({n6228, n56, n6224, n6222, n6220, n5908, n6217, n5267}), 
        .CI(1'b0), .DIFF({n712, n711, n710, n709, n708, n707, n706, n705}), 
        .CO() );
  alu_DW01_sub_12 sub_153 ( .A({n5271, n6021, n6018, n6016, n6011, n6008, 
        n6007, n6004}), .B({n6241, n6239, n6237, n5279, n6234, n6232, n20, n46}), .CI(1'b0), .DIFF({n704, n703, n702, n701, n700, n699, n698, n697}), .CO()
         );
  alu_DW01_sub_13 sub_152 ( .A({n6039, n5277, n6034, n5885, n6032, n6029, 
        n6026, n59}), .B({n6255, n6253, n6251, n6249, n6247, n6245, n6243, n70}), .CI(1'b0), .DIFF({n696, n695, n694, n693, n692, n691, n690, n689}), .CO()
         );
  alu_DW01_sub_14 sub_151 ( .A({n6061, n6059, n6057, n6055, n6052, n21, n5734, 
        n6042}), .B({n6271, n6269, n6267, n3, n6263, n6261, n6259, n6257}), 
        .CI(1'b0), .DIFF({n688, n687, n686, n685, n684, n683, n682, n681}), 
        .CO() );
  alu_DW01_add_7 add_124 ( .A({n5929, n6279, n6277, n67, n5922, n5918, n5916, 
        n5912}), .B({n6167, n6165, n6163, n5904, n5903, n5899, n5895, n9}), 
        .CI(1'b0), .SUM({n423, n422, n421, n420, n419, n418, n417, n416}), 
        .CO() );
  alu_DW01_add_8 add_123 ( .A({n5948, n5947, n5945, n6288, n5940, n5938, n5933, 
        n5931}), .B({n6183, n6181, n6179, n6177, n6175, n6173, n6171, n6169}), 
        .CI(1'b0), .SUM({n415, n414, n413, n412, n411, n410, n409, n408}), 
        .CO() );
  alu_DW01_add_9 add_122 ( .A({n5970, n6296, n5966, n5963, n5960, n5957, n5953, 
        n5952}), .B({n6199, n6197, n6195, n6193, n6191, n6189, n6187, n6185}), 
        .CI(1'b0), .SUM({n407, n406, n405, n404, n403, n402, n401, n400}), 
        .CO() );
  alu_DW01_add_10 add_121 ( .A({n5989, n6308, n5984, n5982, n5980, n6301, 
        n5976, n5974}), .B({n6215, n6213, n6211, n6209, n6207, n6205, n6203, 
        n6201}), .CI(1'b0), .SUM({n399, n398, n397, n396, n395, n394, n393, 
        n392}), .CO() );
  alu_DW01_add_11 add_120 ( .A({n6325, n58, n5268, n5997, n5276, n5995, n5992, 
        n5879}), .B({n6228, n56, n6224, n6222, n5883, n5907, n6217, n5267}), 
        .CI(1'b0), .SUM({n391, n390, n389, n388, n387, n386, n385, n384}), 
        .CO() );
  alu_DW01_add_12 add_119 ( .A({n5272, n6021, n6018, n5278, n6334, n6008, 
        n6007, n6328}), .B({n6241, n6239, n6237, n5280, n6234, n6232, n19, n46}), .CI(1'b0), .SUM({n383, n382, n381, n380, n379, n378, n377, n376}), .CO() );
  alu_DW01_add_13 add_118 ( .A({n6039, n5277, n6034, n5885, n6032, n6029, 
        n6026, n59}), .B({n6255, n6253, n6251, n6249, n6247, n6245, n6243, n70}), .CI(1'b0), .SUM({n375, n374, n373, n372, n371, n370, n369, n368}), .CO() );
  alu_DW01_add_14 add_117 ( .A({n6060, n6058, n6057, n6055, n6051, n6049, 
        n6046, n6043}), .B({n6271, n6269, n6267, n3, n6263, n6261, n6259, 
        n6257}), .CI(1'b0), .SUM({n367, n366, n365, n364, n363, n362, n361, 
        n360}), .CO() );
  alu_DW_mult_uns_23 mult_240 ( .a({n5948, n5947, n5944, n6288, n5941, n5937, 
        n5933, n5932}), .b({n5948, n6290, n5944, n5942, n6286, n5937, n5934, 
        n5931}), .product({n1579, n1578, n1577, n1576, n1575, n1574, n1573, 
        n1572, n1571, n1570, n1569, n1568, n1567, n1566, 
        SYNOPSYS_UNCONNECTED_1, n1564}) );
  alu_DW_mult_uns_22 mult_188 ( .a({n5948, n5947, n5945, n5942, n6286, n5938, 
        n5935, n5932}), .b({n6183, n6181, n6179, n6177, n6175, n6173, n6171, 
        n6169}), .product({n1065, n1064, n1063, n1062, n1061, n1060, n1059, 
        n1058, n1057, n1056, n1055, n1054, n1053, n1052, n1051, n1050}) );
  alu_DW_mult_uns_19 mult_239 ( .a({n5988, n5986, n5984, n5981, n5980, n6301, 
        n5975, n5973}), .b({n5989, n6308, n5983, n5981, n5980, n5978, n5976, 
        n5972}), .product({n1563, n1562, n1561, n1560, n1559, n1558, n1557, 
        n1556, n1555, n1554, n1553, n1552, n1551, n1550, 
        SYNOPSYS_UNCONNECTED_2, n1548}) );
  alu_DW_mult_uns_18 mult_187 ( .a({n5988, n5987, n5984, n5982, n5980, n5977, 
        oprA[38], n5972}), .b({n6215, n6213, n6211, n6209, n6207, n6205, n6203, 
        n6201}), .product({n1049, n1048, n1047, n1046, n1045, n1044, n1043, 
        n1042, n1041, n1040, n1039, n1038, n1037, n1036, n1035, n1034}) );
  alu_DW_mult_uns_11 mult_238 ( .a({n5271, n6022, n6018, n6016, n5285, n6008, 
        n6007, n6328}), .b({n5271, n6021, n6018, n5278, n6011, n6008, n6007, 
        n6004}), .product({n1547, n1546, n1545, n1544, n1543, n1542, n1541, 
        n1540, n1539, n1538, n1537, n1536, n1535, n1534, 
        SYNOPSYS_UNCONNECTED_3, n1532}) );
  alu_DW_mult_uns_10 mult_186 ( .a({n5272, n6021, n6018, n5278, n6334, n6008, 
        n6007, n6004}), .b({n6241, n6239, n6237, n5280, n6234, n6232, n20, n46}), .product({n1033, n1032, n1031, n1030, n1029, n1028, n1027, n1026, n1025, 
        n1024, n1023, n1022, n1021, n1020, n1019, n1018}) );
  alu_DW_mult_uns_15 mult_237 ( .a({n6061, n6058, n6057, n6055, n6051, n6049, 
        n5734, n6042}), .b({n6060, n6058, n6057, n6055, n6052, n6049, n5734, 
        n6043}), .product({n1531, n1530, n1529, n1528, n1527, n1526, n1525, 
        n1524, n1523, n1522, n1521, n1520, n1519, n1518, 
        SYNOPSYS_UNCONNECTED_4, n1516}) );
  alu_DW_mult_uns_14 mult_185 ( .a({n6061, n6059, n6057, n6054, n6051, n6048, 
        n6347, n6041}), .b({n6271, n6269, n6267, n2, n6263, n6261, n6259, 
        n6257}), .product({n1017, n1016, n1015, n1014, n1013, n1012, n1011, 
        n1010, n1009, n1008, n1007, n1006, n1005, n1004, n1003, n1002}) );
  alu_DW_mult_uns_6 mult_214 ( .a({n5929, n5926, n6277, n67, n17, n5918, n5915, 
        n5910}), .b({n6167, n6165, n6163, n5904, n5901, n5899, n5895, n5892}), 
        .product({n1322, n1321, n1320, n1319, n1318, n1317, n1316, n1315, 
        n1314, n1313, n1312, n1311, n1310, n1309, n1308, n1307}) );
  alu_DW_mult_uns_4 mult_213 ( .a({n5970, n5969, n5966, n5963, n5960, n5958, 
        n5955, n5951}), .b({n6199, n6197, n6195, n6193, n6191, oprB[45], n6187, 
        n6185}), .product({n1306, n1305, n1304, n1303, n1302, n1301, n1300, 
        n1299, n1298, n1297, n1296, n1295, n1294, n1293, n1292, n1291}) );
  alu_DW_mult_uns_0 mult_212 ( .a({n6325, n58, n5268, n5997, n5276, n6314, 
        n5992, n5990}), .b({n6228, n56, n6224, n6222, n6220, n5907, n6217, 
        n5267}), .product({n1290, n1289, n1288, n1287, n1286, n1285, n1284, 
        n1283, n1282, n1281, n1280, n1279, n1278, n1277, n1276, n1275}) );
  alu_DW_mult_uns_2 mult_211 ( .a({n6345, n5277, n6034, n37, n6032, n6028, 
        n6025, n59}), .b({n6255, n6253, n6251, n6249, n6247, n15, n6243, n23}), 
        .product({n1274, n1273, n1272, n1271, n1270, n1269, n1268, n1267, 
        n1266, n1265, n1264, n1263, n1262, n1261, n1260, n1259}) );
  alu_DW01_sub_15 sub_174 ( .A({n6061, n6058, n6057, n6055, n6052, n21, n5734, 
        n6043, n6039, n6037, n6034, n5885, n6032, n6342, n6026, n59, n6024, 
        n5282, n6018, n5286, n5285, n6009, n6007, n6004, n5274, n5283, n6000, 
        n44, n5276, n6314, n5992, n5991, n5989, n5986, n5984, oprA[35], n5980, 
        n5977, oprA[38], n5973, n5970, n5969, n5966, n5965, n5961, n5956, 
        n5954, n5952, n5949, n5946, n5945, n5942, n5940, n5937, n5935, n5932, 
        n5928, n5927, n5924, n67, n17, n5919, n5914, n5912}), .B({n6271, n6269, 
        n6267, n3, n6263, n6261, n6259, n6257, n6255, n6253, n6251, n6249, 
        n6247, n6245, n6243, n70, n6241, n6239, n6237, n5280, n6234, n6232, 
        n18, oprB[23], n6228, n6226, n6224, oprB[27], n5882, n5907, n6217, 
        n5267, n6215, n6213, n6211, n6209, oprB[36], n6205, n6203, n6201, 
        n6199, n6197, n6195, n6193, n6191, oprB[45], n6187, n6185, n6183, 
        n6181, n6179, n6177, n6175, n6173, n6171, n6169, n6167, n6165, n6163, 
        n5905, n5903, n5899, n5896, n8}), .CI(1'b0), .DIFF({n936, n935, n934, 
        n933, n932, n931, n930, n929, n928, n927, n926, n925, n924, n923, n922, 
        n921, n920, n919, n918, n917, n916, n915, n914, n913, n912, n911, n910, 
        n909, n908, n907, n906, n905, n904, n903, n902, n901, n900, n899, n898, 
        n897, n896, n895, n894, n893, n892, n891, n890, n889, n888, n887, n886, 
        n885, n884, n883, n882, n881, n880, n879, n878, n877, n876, n875, n874, 
        n873}), .CO() );
  alu_DW01_add_15 add_140 ( .A({n6061, n6058, n6057, n6054, n6051, n21, n5734, 
        n6042, n6039, n5277, n6034, n5885, n6032, n6342, n6026, n59, n5272, 
        n6022, n6018, n6016, n5269, n6009, n5270, n6328, n6003, n6001, n6000, 
        n44, n5276, n5995, n5993, n5879, n5988, n5987, n5983, oprA[35], n5980, 
        n5978, oprA[38], n5974, n5970, n5969, n5966, n5965, n5961, n5956, 
        n5954, n5952, n5948, n5946, n5944, n5942, n5941, n5938, n5935, n5932, 
        n5928, n5926, n5925, n67, n5922, n5919, n5914, n5911}), .B({n6271, 
        n6269, n6267, n3, n6263, n6261, n6259, n6257, n6255, n6253, n6251, 
        n6249, n6247, n6245, n6243, n70, n6241, n6239, n6237, n5280, n6234, 
        n22, oprB[22:23], n6228, n6226, n6224, oprB[27], n5882, n5908, n6217, 
        n5267, n6215, n6213, n6211, n6209, oprB[36], n6205, n6203, n6201, 
        n6199, n6197, n6195, n6193, n6191, oprB[45], n6187, n6185, n6183, 
        n6181, n6179, n6177, n6175, n6173, n6171, n6169, n6167, n6165, n6163, 
        n5905, n5902, n5900, n5896, n9}), .CI(1'b0), .SUM({n615, n614, n613, 
        n612, n611, n610, n609, n608, n607, n606, n605, n604, n603, n602, n601, 
        n600, n599, n598, n597, n596, n595, n594, n593, n592, n591, n590, n589, 
        n588, n587, n586, n585, n584, n583, n582, n581, n580, n579, n578, n577, 
        n576, n575, n574, n573, n572, n571, n570, n569, n568, n567, n566, n565, 
        n564, n563, n562, n561, n560, n559, n558, n557, n556, n555, n554, n553, 
        n552}), .CO() );
  alu_DW_mult_uns_37 mult_193 ( .a({n5989, n5987, n5985, oprA[35], n5980, 
        n5978, oprA[38], n5972, n5970, n5968, n5966, n5963, n5960, n5956, 
        n5954, n5951}), .b({n6215, n6213, n6211, n6209, oprB[36], n6205, n6203, 
        n6201, n6199, n6197, n6195, n6193, n6191, oprB[45], n6187, n6185}), 
        .product({n1129, n1128, n1127, n1126, n1125, n1124, n1123, n1122, 
        n1121, n1120, n1119, n1118, n1117, n1116, n1115, n1114, n1113, n1112, 
        n1111, n1110, n1109, n1108, n1107, n1106, n1105, n1104, n1103, n1102, 
        n1101, n1100, n1099, n1098}) );
  alu_DW_mult_uns_36 mult_192 ( .a({oprA[0], n6059, n6056, n6053, n6351, n29, 
        n6045, n6041, oprA[8], n6037, n6035, n37, n6031, n6342, n6025, 
        oprA[15]}), .b({n6271, n6269, n6267, n2, n6263, n6261, n6259, n6257, 
        n6255, n6253, n6251, n6249, n6247, oprB[13], n6243, oprB[15]}), 
        .product({n1097, n1096, n1095, n1094, n1093, n1092, n1091, n1090, 
        n1089, n1088, n1087, n1086, n1085, n1084, n1083, n1082, n1081, n1080, 
        n1079, n1078, n1077, n1076, n1075, n1074, n1073, n1072, n1071, n1070, 
        n1069, n1068, n1067, n1066}) );
  alu_DW_mult_uns_38 mult_219 ( .a({n5949, n5946, n5944, n5942, n5940, n5937, 
        n5935, n5931, n5928, n5927, n5925, n67, n17, n5919, n5914, n5910}), 
        .b({n6183, n6181, n6179, n6177, n6175, n6173, n6171, n6169, n6167, 
        n6165, n6163, n5905, n5903, n5899, n5896, n9}), .product({n1386, n1385, 
        n1384, n1383, n1382, n1381, n1380, n1379, n1378, n1377, n1376, n1375, 
        n1374, n1373, n1372, n1371, n1370, n1369, n1368, n1367, n1366, n1365, 
        n1364, n1363, n1362, n1361, n1360, n1359, n1358, n1357, n1356, n1355})
         );
  alu_DW01_sub_17 sub_170 ( .A({n5989, n5987, n5984, n5981, n5980, n6301, 
        n5975, n5973, n6297, n5968, n5966, n5964, n5960, n5958, n5955, n5952, 
        n5948, n6290, n5944, n5942, n5941, n5938, n5933, n5932, n6282, n5926, 
        n5924, n66, n6275, n5919, n5914, n5912}), .B({n6215, n6213, n6211, 
        n6209, n6207, n6205, n6203, n6201, n6199, n6197, n6195, n6193, n6191, 
        n6189, n6187, n6185, n6183, n6181, n6179, n6177, n6175, n6173, n6171, 
        n6169, n6167, n6165, n6163, n5905, n5902, n5900, n5897, n7}), .CI(1'b0), .DIFF({n872, n871, n870, n869, n868, n867, n866, n865, n864, n863, n862, 
        n861, n860, n859, n858, n857, n856, n855, n854, n853, n852, n851, n850, 
        n849, n848, n847, n846, n845, n844, n843, n842, n841}), .CO() );
  alu_DW01_add_16 add_135 ( .A({n6061, n6059, n6057, n6055, n6052, n6049, 
        n6046, n6042, n6039, n6037, n6034, n5885, n6032, n6029, n6026, n59, 
        n5271, n6022, n6018, n5286, n5269, n6332, n5270, n6328, n5274, n6001, 
        n6000, n6317, n5275, n6314, n5992, n5990}), .B({n6271, n6269, n6267, 
        n3, n6263, n6261, n6259, n6257, n6255, n6253, n6251, n6249, n6247, 
        n6245, n6243, n70, n6241, n6239, n6237, n5279, n6234, n6232, n20, n46, 
        n6228, n6226, n6224, oprB[27], n5882, n5907, n6217, oprB[31]}), .CI(
        1'b0), .SUM({n519, n518, n517, n516, n515, n514, n513, n512, n511, 
        n510, n509, n508, n507, n506, n505, n504, n503, n502, n501, n500, n499, 
        n498, n497, n496, n495, n494, n493, n492, n491, n490, n489, n488}), 
        .CO() );
  alu_DW01_add_17 add_136 ( .A({n5988, n5986, n5983, n5982, n5980, n5977, 
        n5975, n5974, n5970, n5969, n45, n5964, n5960, n5957, n5955, n5952, 
        n5949, n6290, n5945, n6288, n5940, n5938, n5933, n5932, n6282, n5927, 
        n5925, oprA[59], n16, n5919, n5914, n5912}), .B({n6215, n6213, n6211, 
        n6209, n6207, n6205, n6203, n6201, n6199, n6197, n6195, n6193, n6191, 
        n6189, n6187, n6185, n6183, n6181, n6179, n6177, n6175, n6173, n6171, 
        n6169, n6167, n6165, n6163, n5906, n5903, oprB[61], n5897, oprB[63]}), 
        .CI(1'b0), .SUM({n551, n550, n549, n548, n547, n546, n545, n544, n543, 
        n542, n541, n540, n539, n538, n537, n536, n535, n534, n533, n532, n531, 
        n530, n529, n528, n527, n526, n525, n524, n523, n522, n521, n520}), 
        .CO() );
  alu_DW01_sub_16 sub_169 ( .A({n6060, n6058, n6057, n6054, n6052, n6049, 
        n6046, n6043, n6039, n6037, n6034, n5885, n6032, n6029, n6026, n59, 
        n6024, n5282, n6018, n6016, n5285, n6332, n6330, n6004, n6003, n5283, 
        n5268, n27, n5275, n6314, n5993, n5991}), .B({n6271, n6269, n6267, n3, 
        n6263, n6261, n6259, n6257, n6255, n6253, n6251, n6249, n6247, n6245, 
        n6243, n70, n6241, n6239, n6237, n5280, n6234, n6232, n19, n46, n6228, 
        n6226, n6224, oprB[27], n5883, n5908, n6217, n5266}), .CI(1'b0), 
        .DIFF({n840, n839, n838, n837, n836, n835, n834, n833, n832, n831, 
        n830, n829, n828, n827, n826, n825, n824, n823, n822, n821, n820, n819, 
        n818, n817, n816, n815, n814, n813, n812, n811, n810, n809}), .CO() );
  alu_DW_mult_uns_25 mult_245 ( .a({n5989, n5987, n5983, n5982, n6303, n5978, 
        n5975, n5973, n6297, n5968, n5966, n5964, n5960, n5956, n5955, n5952}), 
        .b({n5988, n5986, n5984, oprA[35:36], n5978, oprA[38], n5972, n5970, 
        n5968, oprA[42], n5963, n5960, n5956, n5954, n5951}), .product({n1643, 
        n1642, n1641, n1640, n1639, n1638, n1637, n1636, n1635, n1634, n1633, 
        n1632, n1631, n1630, n1629, n1628, n1627, n1626, n1625, n1624, n1623, 
        n1622, n1621, n1620, n1619, n1618, n1617, n1616, n1615, n1614, 
        SYNOPSYS_UNCONNECTED_5, n1612}) );
  alu_DW_mult_uns_24 mult_244 ( .a({n6061, n6058, n6057, n6054, n6052, n21, 
        n6046, n6041, n6345, n6038, n6035, n37, n6031, n6342, n6025, n59}), 
        .b({n6060, n6059, n6057, n6053, n6350, n29, n6045, n6041, oprA[8:11], 
        n6031, n6028, n6025, oprA[15]}), .product({n1611, n1610, n1609, n1608, 
        n1607, n1606, n1605, n1604, n1603, n1602, n1601, n1600, n1599, n1598, 
        n1597, n1596, n1595, n1594, n1593, n1592, n1591, n1590, n1589, n1588, 
        n1587, n1586, n1585, n1584, n1583, n1582, SYNOPSYS_UNCONNECTED_6, 
        n1580}) );
  alu_DW_mult_uns_27 mult_270 ( .a({n5271, n5282, n6018, n5278, n5285, n6008, 
        n6007, n6328, n6003, n5283, n6319, n27, n5275, n6314, n5993, n5879}), 
        .b({n6024, n6021, n6019, oprA[19], n6012, n6009, n6006, n6327, 
        oprA[24], n52, n5268, n5998, n5275, n6314, n5992, n5990}), .product({
        n1836, n1835, n1834, n1833, n1832, n1831, n1830, n1829, n1828, n1827, 
        n1826, n1825, n1824, n1823, n1822, n1821, n1820, n1819, n1818, n1817, 
        n1816, n1815, n1814, n1813, n1812, n1811, n1810, n1809, n1808, n1807, 
        SYNOPSYS_UNCONNECTED_7, n1805}) );
  alu_DW_mult_uns_26 mult_271 ( .a({n5948, n5947, n5945, n5942, n6286, n5937, 
        n5934, n5931, n6282, n5927, n5925, n67, n6275, n5919, n5914, n5911}), 
        .b({n5948, n5947, n5945, n5942, n5941, n5938, n5935, n5931, n5928, 
        n6279, oprA[58], n66, n6275, n5919, n5914, n5910}), .product({n1868, 
        n1867, n1866, n1865, n1864, n1863, n1862, n1861, n1860, n1859, n1858, 
        n1857, n1856, n1855, n1854, n1853, n1852, n1851, n1850, n1849, n1848, 
        n1847, n1846, n1845, n1844, n1843, n1842, n1841, n1840, n1839, 
        SYNOPSYS_UNCONNECTED_8, n1837}) );
  alu_DW01_add_20 add_129 ( .A({n6024, n5282, n6018, n6016, n5285, n6008, 
        n6007, n6004, n6003, n6322, n5268, n5997, n5276, n5995, n5993, n5991}), 
        .B({n6241, n6239, n6237, n5279, n6234, n6232, n19, n46, n6228, n56, 
        n6224, n6222, n5883, n5908, n6217, n5266}), .CI(1'b0), .SUM({n455, 
        n454, n453, n452, n451, n450, n449, n448, n447, n446, n445, n444, n443, 
        n442, n441, n440}), .CO() );
  alu_DW01_add_18 add_131 ( .A({n5949, n5947, n5945, n5942, n5941, n5937, 
        n5933, n5932, n5929, n5927, n5924, n67, n6275, n5918, n5916, n5911}), 
        .B({n6183, n6181, n6179, n6177, n6175, n6173, n6171, n6169, n6167, 
        n6165, n6163, n5904, n5902, n5900, n5896, n9}), .CI(1'b0), .SUM({n487, 
        n486, n485, n484, n483, n482, n481, n480, n479, n478, n477, n476, n475, 
        n474, n473, n472}), .CO() );
  alu_DW01_sub_19 sub_164 ( .A({n5988, n6308, n5984, n5981, n5980, n5977, 
        n5975, n5972, n6297, n5969, n5966, n5965, n5960, n5958, n5953, n5952}), 
        .B({n6215, n6213, n6211, n6209, n6207, n6205, n6203, n6201, n6199, 
        n6197, n6195, n6193, n6191, oprB[45], n6187, n6185}), .CI(1'b0), 
        .DIFF({n792, n791, n790, n789, n788, n787, n786, n785, n784, n783, 
        n782, n781, n780, n779, n778, n777}), .CO() );
  alu_DW01_sub_18 sub_165 ( .A({n5948, n6290, n5944, n5942, n5940, n5938, 
        n5934, n5931, n5929, n5926, n6277, n67, n17, n5918, n5916, n5911}), 
        .B({n6183, n6181, n6179, n6177, n6175, n6173, n6171, n6169, n6167, 
        n6165, n6163, n5905, n5902, n5900, n5897, n9}), .CI(1'b0), .DIFF({n808, 
        n807, n806, n805, n804, n803, n802, n801, n800, n799, n798, n797, n796, 
        n795, n794, n793}), .CO() );
  alu_DW01_sub_21 sub_162 ( .A({n6061, n6059, n6057, n6054, n6052, n21, n6046, 
        n6042, n6039, n6038, n6034, n5885, n6032, n6029, n6026, n59}), .B({
        n6271, n6269, n6267, n3, n6263, n6261, n6259, n6257, n6255, n6253, 
        n6251, n6249, n6247, n15, n6243, oprB[15]}), .CI(1'b0), .DIFF({n760, 
        n759, n758, n757, n756, n755, n754, n753, n752, n751, n750, n749, n748, 
        n747, n746, n745}), .CO() );
  alu_DW01_sub_20 sub_163 ( .A({n5272, n6022, n6018, n5286, n5269, n6008, 
        n5270, n6004, n5274, n5283, n6319, n43, n5276, n6315, n5993, n5880}), 
        .B({n6241, n6239, n6237, n5280, n6234, n6232, n20, n46, n6228, n56, 
        n6224, n6222, n6220, n5907, n6217, n5266}), .CI(1'b0), .DIFF({n776, 
        n775, n774, n773, n772, n771, n770, n769, n768, n767, n766, n765, n764, 
        n763, n762, n761}), .CO() );
  alu_DW_mult_uns_29 mult_265 ( .a({n5970, n5969, n5966, n5965, n5961, n5957, 
        n5955, n5952}), .b({n5970, n6296, n45, n5964, n5961, n5957, n5955, 
        n5951}), .product({n1788, n1787, n1786, n1785, n1784, n1783, n1782, 
        n1781, n1780, n1779, n1778, n1777, n1776, n1775, 
        SYNOPSYS_UNCONNECTED_9, n1773}) );
  alu_DW_mult_uns_31 mult_263 ( .a({n6039, n5277, n6034, n5885, n6032, n6028, 
        n6026, n59}), .b({n6345, n6037, n6034, n5885, n6032, n6028, n6026, n59}), .product({n1756, n1755, n1754, n1753, n1752, n1751, n1750, n1749, n1748, 
        n1747, n1746, n1745, n1744, n1743, SYNOPSYS_UNCONNECTED_10, n1741}) );
  alu_DW_mult_uns_30 mult_264 ( .a({n6325, n58, n5268, n43, n5276, n5995, 
        n5992, n5879}), .b({n6003, n5283, n6000, n27, n5276, n6314, n5992, 
        n5990}), .product({n1772, n1771, n1770, n1769, n1768, n1767, n1766, 
        n1765, n1764, n1763, n1762, n1761, n1760, n1759, 
        SYNOPSYS_UNCONNECTED_11, n1757}) );
  alu_DW_mult_uns_28 mult_266 ( .a({n5929, n5926, n5925, n66, n5922, n5919, 
        n5916, n5911}), .b({n6282, n5926, n5924, n66, n6275, n5919, n5915, 
        n5910}), .product({n1804, n1803, n1802, n1801, n1800, n1799, n1798, 
        n1797, n1796, n1795, n1794, n1793, n1792, n1791, 
        SYNOPSYS_UNCONNECTED_12, n1789}) );
  alu_DW01_add_25 add_128 ( .A({n6060, n6059, n6057, n6055, n6051, n6049, 
        n5734, n6043, n6039, n5277, n6034, n5885, n6032, n6029, n6026, 
        oprA[15]}), .B({n6271, n6269, n6267, n3, n6263, n6261, n6259, n6257, 
        n6255, n6253, n6251, n6249, n6247, n6245, n6243, n23}), .CI(1'b0), 
        .SUM({n439, n438, n437, n436, n435, n434, n433, n432, n431, n430, n429, 
        n428, n427, n426, n425, n424}), .CO() );
  alu_DW01_add_26 add_130 ( .A({n5989, n5986, n5983, n5982, n6303, n5978, 
        n5976, n5974, n5970, n6296, n45, n5963, n5960, n5957, n5953, n5952}), 
        .B({n6215, n6213, n6211, n6209, n6207, n6205, n6203, n6201, n6199, 
        n6197, n6195, n6193, n6191, oprB[45], n6187, n6185}), .CI(1'b0), .SUM(
        {n471, n470, n469, n468, n467, n466, n465, n464, n463, n462, n461, 
        n460, n459, n458, n457, n456}), .CO() );
  alu_DW_mult_uns_105 mult_218 ( .a({oprA[16], n5281, n6019, n6015, n6013, 
        n6009, n6007, n6328, n6003, n5283, n6000, n27, n5275, n6314, n5993, 
        n5990}), .b({n6241, n6239, n6237, oprB[19], n6234, n6232, n19, n46, 
        n6228, n6226, n6224, oprB[27], n5883, n5907, n6217, n5266}), .product(
        {n1354, n1353, n1352, n1351, n1350, n1349, n1348, n1347, n1346, n1345, 
        n1344, n1343, n1342, n1341, n1340, n1339, n1338, n1337, n1336, n1335, 
        n1334, n1333, n1332, n1331, n1330, n1329, n1328, n1327, n1326, n1325, 
        n1324, n1323}) );
  INVX2 U6 ( .A(oprB[20]), .Y(n6235) );
  INVX2 U7 ( .A(n6040), .Y(n6043) );
  INVX2 U8 ( .A(oprB[19]), .Y(n6236) );
  INVX2 U9 ( .A(oprA[33]), .Y(n6309) );
  INVX2 U10 ( .A(n5909), .Y(n5910) );
  INVX2 U11 ( .A(oprA[15]), .Y(n5881) );
  INVX1 U12 ( .A(oprA[23]), .Y(n1) );
  INVX2 U13 ( .A(oprB[32]), .Y(n6216) );
  INVX4 U14 ( .A(n6359), .Y(n6061) );
  INVX2 U15 ( .A(n6329), .Y(n6327) );
  AND2X2 U16 ( .A(n19), .B(n1), .Y(n9176) );
  INVX2 U17 ( .A(n6289), .Y(n6288) );
  INVX2 U18 ( .A(oprA[47]), .Y(n5950) );
  INVX2 U19 ( .A(n6155), .Y(n5889) );
  INVX2 U20 ( .A(n6033), .Y(n6035) );
  INVX2 U21 ( .A(oprA[10]), .Y(n6033) );
  INVX8 U22 ( .A(n6020), .Y(n6021) );
  INVX8 U23 ( .A(n6186), .Y(n6185) );
  INVX2 U24 ( .A(oprA[41]), .Y(n5967) );
  INVX4 U25 ( .A(n6280), .Y(n5927) );
  INVX2 U26 ( .A(oprA[57]), .Y(n6280) );
  INVX4 U27 ( .A(n6353), .Y(n6053) );
  INVX2 U28 ( .A(oprA[3]), .Y(n6353) );
  INVX2 U29 ( .A(oprB[22]), .Y(n6231) );
  BUFX4 U30 ( .A(n6006), .Y(n5270) );
  INVX8 U31 ( .A(n6196), .Y(n6195) );
  INVX2 U32 ( .A(mult32_B[14]), .Y(n5593) );
  OR2X2 U33 ( .A(n6259), .B(n10210), .Y(n10507) );
  AND2X2 U34 ( .A(n6259), .B(n6257), .Y(n10216) );
  INVX8 U35 ( .A(n6194), .Y(n6193) );
  BUFX4 U36 ( .A(n6265), .Y(n2) );
  BUFX2 U37 ( .A(n6265), .Y(n3) );
  INVX1 U38 ( .A(n6266), .Y(n6265) );
  INVX1 U39 ( .A(n6349), .Y(n4) );
  INVX1 U40 ( .A(n4), .Y(n5) );
  INVX1 U41 ( .A(n4), .Y(n6) );
  INVX2 U42 ( .A(mult32_B[9]), .Y(n5657) );
  INVX2 U43 ( .A(mult32_B[11]), .Y(n5590) );
  INVX8 U44 ( .A(n6188), .Y(n6187) );
  INVX8 U45 ( .A(n6184), .Y(n6183) );
  AND2X2 U46 ( .A(n6185), .B(n5967), .Y(n7585) );
  AND2X2 U47 ( .A(n6185), .B(n6188), .Y(n7611) );
  AND2X2 U48 ( .A(n6187), .B(n6185), .Y(n7586) );
  INVX2 U49 ( .A(n6333), .Y(n6332) );
  BUFX2 U50 ( .A(n5893), .Y(n7) );
  BUFX2 U51 ( .A(n5893), .Y(n8) );
  BUFX2 U52 ( .A(n5893), .Y(n9) );
  INVX1 U53 ( .A(n5891), .Y(n5893) );
  INVX2 U54 ( .A(mult32_B[30]), .Y(n5460) );
  BUFX4 U55 ( .A(n6024), .Y(n5271) );
  INVX4 U56 ( .A(n6023), .Y(n6024) );
  INVX2 U57 ( .A(oprB[37]), .Y(n6206) );
  AND2X1 U58 ( .A(n268), .B(n7418), .Y(n7420) );
  AND2X1 U59 ( .A(n4647), .B(n4693), .Y(n10283) );
  AND2X1 U60 ( .A(n5888), .B(n6344), .Y(n9634) );
  AND2X1 U61 ( .A(n4641), .B(n4686), .Y(n9243) );
  INVX2 U62 ( .A(n5), .Y(n29) );
  AND2X1 U63 ( .A(n5821), .B(n6248), .Y(n9845) );
  AND2X1 U64 ( .A(n963), .B(n1461), .Y(n10569) );
  AND2X1 U65 ( .A(n4707), .B(n4689), .Y(n9564) );
  AND2X1 U66 ( .A(n4643), .B(n4687), .Y(n9335) );
  AND2X1 U67 ( .A(n4638), .B(n4680), .Y(n8526) );
  AND2X1 U68 ( .A(n4635), .B(n4678), .Y(n8231) );
  AND2X1 U69 ( .A(n4705), .B(n4673), .Y(n7537) );
  AND2X1 U70 ( .A(n6171), .B(n6170), .Y(n5792) );
  AND2X1 U71 ( .A(n4627), .B(n4663), .Y(n6478) );
  AND2X1 U72 ( .A(n5400), .B(n5731), .Y(n6505) );
  AND2X1 U73 ( .A(n4704), .B(n4664), .Y(n6496) );
  AND2X1 U74 ( .A(n5647), .B(n5646), .Y(mult32_A[15]) );
  AND2X1 U75 ( .A(n6076), .B(n6351), .Y(n6465) );
  AND2X1 U76 ( .A(n10373), .B(n5399), .Y(n5738) );
  AND2X1 U77 ( .A(n1138), .B(n1485), .Y(n10391) );
  AND2X1 U78 ( .A(n1000), .B(n1481), .Y(n10245) );
  AND2X1 U79 ( .A(n945), .B(n1450), .Y(n10396) );
  AND2X1 U80 ( .A(n948), .B(n1452), .Y(n10388) );
  AND2X1 U81 ( .A(n6247), .B(n10218), .Y(n9727) );
  AND2X1 U82 ( .A(n1157), .B(n5212), .Y(n9698) );
  AND2X1 U83 ( .A(n1158), .B(n1460), .Y(n9708) );
  INVX2 U84 ( .A(n6246), .Y(n6245) );
  AND2X1 U85 ( .A(n957), .B(n1458), .Y(n9653) );
  AND2X1 U86 ( .A(n628), .B(n1420), .Y(n9502) );
  AND2X1 U87 ( .A(n666), .B(n1441), .Y(n9205) );
  AND2X1 U88 ( .A(n357), .B(n1412), .Y(n9336) );
  AND2X1 U89 ( .A(n354), .B(n1410), .Y(n9344) );
  AND2X1 U90 ( .A(n620), .B(n1418), .Y(n8623) );
  AND2X1 U91 ( .A(n621), .B(n1419), .Y(n8639) );
  AND2X1 U92 ( .A(n619), .B(n1417), .Y(n8598) );
  AND2X1 U93 ( .A(n4706), .B(n4681), .Y(n8541) );
  AND2X1 U94 ( .A(n5656), .B(n5588), .Y(n10093) );
  AND2X1 U95 ( .A(n344), .B(n1405), .Y(n8424) );
  AND2X1 U96 ( .A(n4637), .B(n4679), .Y(n8325) );
  AND2X1 U97 ( .A(n329), .B(n1397), .Y(n8194) );
  AND2X1 U98 ( .A(n280), .B(n1237), .Y(n8326) );
  AND2X1 U99 ( .A(n277), .B(n1235), .Y(n8334) );
  INVX1 U100 ( .A(oprA[60]), .Y(n5920) );
  AND2X1 U101 ( .A(n1149), .B(n5210), .Y(n7666) );
  AND2X1 U102 ( .A(n1150), .B(n1245), .Y(n7675) );
  AND2X1 U103 ( .A(n287), .B(n1243), .Y(n7621) );
  AND2X1 U104 ( .A(n272), .B(n1233), .Y(n7481) );
  AND2X1 U105 ( .A(n232), .B(n1210), .Y(n6832) );
  AND2X1 U106 ( .A(n205), .B(n1193), .Y(n7318) );
  BUFX2 U107 ( .A(n5921), .Y(n16) );
  AND2X1 U111 ( .A(n2553), .B(n6102), .Y(n6674) );
  AND2X1 U112 ( .A(n215), .B(n1201), .Y(n6589) );
  AND2X1 U113 ( .A(n216), .B(n1202), .Y(n6606) );
  AND2X1 U114 ( .A(n214), .B(n1200), .Y(n6563) );
  AND2X1 U115 ( .A(n6731), .B(n5451), .Y(n5742) );
  AND2X1 U116 ( .A(n208), .B(n1195), .Y(n7310) );
  INVX2 U117 ( .A(n5920), .Y(n5922) );
  AND2X1 U118 ( .A(n199), .B(n1186), .Y(mult32_B[7]) );
  AND2X1 U119 ( .A(n6076), .B(n6011), .Y(n6446) );
  AND2X1 U120 ( .A(n197), .B(n1185), .Y(mult32_B[8]) );
  INVX2 U121 ( .A(n5894), .Y(n5897) );
  INVX1 U122 ( .A(n10453), .Y(n41) );
  AND2X1 U126 ( .A(n5469), .B(n5470), .Y(n10353) );
  AND2X1 U127 ( .A(n986), .B(n1474), .Y(n10052) );
  AND2X1 U128 ( .A(n984), .B(n1472), .Y(n10039) );
  INVX1 U129 ( .A(op[2]), .Y(n6472) );
  AND2X1 U130 ( .A(n339), .B(n1402), .Y(n8298) );
  AND2X1 U131 ( .A(n314), .B(n1258), .Y(n7993) );
  AND2X1 U132 ( .A(n5617), .B(n1388), .Y(n8006) );
  INVX2 U133 ( .A(oprA[58]), .Y(n5923) );
  INVX1 U134 ( .A(n5920), .Y(n5921) );
  AND2X1 U135 ( .A(n941), .B(n1449), .Y(n9464) );
  INVX1 U136 ( .A(n1386), .Y(n35) );
  AND2X1 U137 ( .A(n348), .B(n1408), .Y(n8463) );
  OR2X1 U141 ( .A(n105), .B(n2337), .Y(n8467) );
  AND2X1 U142 ( .A(n347), .B(n1676), .Y(n8459) );
  INVX1 U143 ( .A(n839), .Y(n54) );
  AND2X1 U144 ( .A(n1137), .B(n1736), .Y(n10344) );
  AND2X1 U145 ( .A(n1140), .B(n1737), .Y(n10407) );
  AND2X1 U146 ( .A(n1136), .B(n1735), .Y(n10337) );
  AND2X1 U147 ( .A(n1131), .B(n1734), .Y(n10277) );
  AND2X1 U148 ( .A(n1130), .B(n1733), .Y(n10270) );
  AND2X1 U149 ( .A(n998), .B(n1732), .Y(n10203) );
  AND2X1 U150 ( .A(n997), .B(n1731), .Y(n10196) );
  AND2X1 U151 ( .A(n995), .B(n1730), .Y(n10128) );
  AND2X1 U152 ( .A(n994), .B(n1729), .Y(n10121) );
  AND2X1 U183 ( .A(n988), .B(n1728), .Y(n10065) );
  AND2X1 U184 ( .A(n987), .B(n1727), .Y(n10058) );
  AND2X1 U185 ( .A(n982), .B(n1726), .Y(n10014) );
  AND2X1 U186 ( .A(n981), .B(n1725), .Y(n10007) );
  AND2X1 U187 ( .A(n980), .B(n1723), .Y(n9950) );
  AND2X1 U188 ( .A(n979), .B(n1722), .Y(n9943) );
  AND2X1 U189 ( .A(n974), .B(n1721), .Y(n9884) );
  AND2X1 U190 ( .A(n973), .B(n1720), .Y(n9877) );
  AND2X1 U191 ( .A(n968), .B(n1719), .Y(n9830) );
  AND2X1 U192 ( .A(n967), .B(n1718), .Y(n9823) );
  AND2X1 U193 ( .A(n962), .B(n1717), .Y(n9762) );
  AND2X1 U194 ( .A(n961), .B(n1716), .Y(n9755) );
  AND2X1 U195 ( .A(n960), .B(n1715), .Y(n9684) );
  AND2X1 U196 ( .A(n959), .B(n1714), .Y(n9677) );
  AND2X1 U197 ( .A(n955), .B(n1713), .Y(n9606) );
  AND2X1 U198 ( .A(n954), .B(n1712), .Y(n9599) );
  AND2X1 U199 ( .A(n944), .B(n1711), .Y(n9546) );
  AND2X1 U200 ( .A(n679), .B(n1702), .Y(n9355) );
  AND2X1 U201 ( .A(n675), .B(n1701), .Y(n9299) );
  AND2X1 U202 ( .A(n674), .B(n1700), .Y(n9292) );
  AND2X1 U203 ( .A(n669), .B(n1699), .Y(n9237) );
  AND2X1 U204 ( .A(n668), .B(n1698), .Y(n9230) );
  AND2X1 U205 ( .A(n664), .B(n1697), .Y(n9163) );
  AND2X1 U206 ( .A(n663), .B(n1696), .Y(n9156) );
  AND2X1 U207 ( .A(n661), .B(n1695), .Y(n9088) );
  AND2X1 U208 ( .A(n660), .B(n1694), .Y(n9081) );
  AND2X1 U209 ( .A(n654), .B(n1693), .Y(n9030) );
  AND2X1 U210 ( .A(n653), .B(n1692), .Y(n9023) );
  AND2X1 U211 ( .A(n648), .B(n1691), .Y(n8981) );
  AND2X1 U212 ( .A(n644), .B(n1687), .Y(n8904) );
  AND2X1 U213 ( .A(n639), .B(n1686), .Y(n8848) );
  AND2X1 U214 ( .A(n638), .B(n1685), .Y(n8841) );
  AND2X1 U215 ( .A(n633), .B(n1684), .Y(n8796) );
  AND2X1 U216 ( .A(n632), .B(n1683), .Y(n8789) );
  AND2X1 U217 ( .A(n627), .B(n1682), .Y(n8733) );
  AND2X1 U218 ( .A(n618), .B(n1679), .Y(n8575) );
  AND2X1 U219 ( .A(n353), .B(n1678), .Y(n8523) );
  AND2X1 U220 ( .A(n342), .B(n1674), .Y(n8345) );
  AND2X1 U221 ( .A(n337), .B(n1672), .Y(n8282) );
  AND2X1 U222 ( .A(n331), .B(n1670), .Y(n8218) );
  AND2X1 U223 ( .A(n327), .B(n1669), .Y(n8151) );
  AND2X1 U224 ( .A(n326), .B(n1668), .Y(n8144) );
  AND2X1 U225 ( .A(n324), .B(n1667), .Y(n8076) );
  AND2X1 U226 ( .A(n323), .B(n1666), .Y(n8069) );
  AND2X1 U227 ( .A(n317), .B(n1665), .Y(n8019) );
  AND2X1 U228 ( .A(n316), .B(n1664), .Y(n8012) );
  AND2X1 U229 ( .A(n312), .B(n1663), .Y(n7968) );
  AND2X1 U230 ( .A(n311), .B(n1662), .Y(n7961) );
  AND2X1 U231 ( .A(n310), .B(n1660), .Y(n7905) );
  AND2X1 U232 ( .A(n309), .B(n1659), .Y(n7898) );
  AND2X1 U233 ( .A(n304), .B(n1658), .Y(n7840) );
  AND2X1 U234 ( .A(n303), .B(n1657), .Y(n7833) );
  AND2X1 U235 ( .A(n298), .B(n1656), .Y(n7789) );
  AND2X1 U236 ( .A(n297), .B(n1655), .Y(n7782) );
  AND2X1 U237 ( .A(n292), .B(n1654), .Y(n7727) );
  AND2X1 U238 ( .A(n291), .B(n1653), .Y(n7720) );
  AND2X1 U239 ( .A(n290), .B(n1652), .Y(n7652) );
  AND2X1 U240 ( .A(n289), .B(n1651), .Y(n7645) );
  AND2X1 U241 ( .A(n285), .B(n1650), .Y(n7578) );
  AND2X1 U242 ( .A(n284), .B(n1649), .Y(n7571) );
  AND2X1 U243 ( .A(n276), .B(n1648), .Y(n7519) );
  AND2X1 U244 ( .A(n275), .B(n1647), .Y(n7512) );
  AND2X1 U245 ( .A(n270), .B(n1646), .Y(n7467) );
  AND2X1 U246 ( .A(n269), .B(n1645), .Y(n7460) );
  AND2X1 U247 ( .A(n267), .B(n1644), .Y(n7401) );
  AND2X1 U248 ( .A(n264), .B(n1565), .Y(n7329) );
  AND2X1 U249 ( .A(n260), .B(n1549), .Y(n7274) );
  AND2X1 U250 ( .A(n259), .B(n1533), .Y(n7267) );
  AND2X1 U251 ( .A(n5345), .B(n5344), .Y(n7208) );
  AND2X1 U252 ( .A(n254), .B(n1517), .Y(n7201) );
  AND2X1 U253 ( .A(n5322), .B(n5321), .Y(n7133) );
  AND2X1 U254 ( .A(n252), .B(n1515), .Y(n7126) );
  AND2X1 U255 ( .A(n251), .B(n1514), .Y(n7063) );
  AND2X1 U256 ( .A(n250), .B(n1513), .Y(n7056) );
  AND2X1 U257 ( .A(n244), .B(n1512), .Y(n7006) );
  AND2X1 U258 ( .A(n243), .B(n1511), .Y(n6999) );
  AND2X1 U259 ( .A(n5330), .B(n5329), .Y(n6953) );
  AND2X1 U260 ( .A(n236), .B(n1507), .Y(n6879) );
  AND2X1 U261 ( .A(n231), .B(n1506), .Y(n6823) );
  AND2X1 U262 ( .A(n230), .B(n1505), .Y(n6816) );
  AND2X1 U263 ( .A(n225), .B(n1504), .Y(n6767) );
  AND2X1 U264 ( .A(n224), .B(n1503), .Y(n6760) );
  AND2X1 U265 ( .A(n219), .B(n1502), .Y(n6699) );
  AND2X1 U266 ( .A(n218), .B(n1501), .Y(n6692) );
  AND2X1 U267 ( .A(n217), .B(n1500), .Y(n6621) );
  AND2X1 U268 ( .A(n213), .B(n1499), .Y(n6538) );
  AND2X1 U269 ( .A(n204), .B(n1498), .Y(n6475) );
  AND2X1 U270 ( .A(n5671), .B(n5670), .Y(n10567) );
  INVX1 U271 ( .A(n6334), .Y(n5273) );
  AND2X1 U272 ( .A(n1148), .B(n1489), .Y(n7433) );
  AND2X1 U273 ( .A(n2935), .B(n6086), .Y(n10583) );
  AND2X1 U274 ( .A(n2934), .B(n6086), .Y(n10528) );
  OR2X1 U275 ( .A(n10527), .B(n2334), .Y(n10529) );
  OR2X1 U276 ( .A(n2086), .B(n2339), .Y(n10591) );
  AND2X1 U277 ( .A(n1142), .B(n1739), .Y(n10590) );
  AND2X1 U278 ( .A(n70), .B(n6036), .Y(n9613) );
  AND2X1 U279 ( .A(n5267), .B(n6324), .Y(n8587) );
  OR2X1 U280 ( .A(n6282), .B(n6159), .Y(n6549) );
  AND2X1 U281 ( .A(n4712), .B(n4692), .Y(n10305) );
  AND2X1 U282 ( .A(n10355), .B(n6351), .Y(n10308) );
  AND2X1 U283 ( .A(n4645), .B(n4691), .Y(n10233) );
  AND2X1 U284 ( .A(n4644), .B(n4688), .Y(n9549) );
  AND2X1 U285 ( .A(n9688), .B(n6351), .Y(n10302) );
  AND2X1 U286 ( .A(n4711), .B(n4685), .Y(n9263) );
  OR2X1 U287 ( .A(n6064), .B(n6336), .Y(n8599) );
  OR2X1 U288 ( .A(n6217), .B(n8583), .Y(n8876) );
  OR2X1 U289 ( .A(n5988), .B(n6204), .Y(n8101) );
  AND2X1 U290 ( .A(n4634), .B(n4676), .Y(n8183) );
  AND2X1 U291 ( .A(n4633), .B(n4672), .Y(n7522) );
  AND2X1 U292 ( .A(n6171), .B(n6284), .Y(n7168) );
  AND2X1 U293 ( .A(n4704), .B(n4650), .Y(n7421) );
  AND2X1 U294 ( .A(n4628), .B(n4668), .Y(n7162) );
  AND2X1 U295 ( .A(n5577), .B(n5576), .Y(mult32_A[12]) );
  AND2X1 U296 ( .A(n6076), .B(n6342), .Y(n6454) );
  OR2X1 U297 ( .A(n6243), .B(n9609), .Y(n9913) );
  AND2X1 U298 ( .A(n6257), .B(n6358), .Y(n10156) );
  AND2X1 U299 ( .A(n6351), .B(n9639), .Y(n9701) );
  AND2X1 U300 ( .A(n4648), .B(n5629), .Y(n10430) );
  INVX1 U301 ( .A(oprB[7]), .Y(n6258) );
  AND2X1 U302 ( .A(n6351), .B(n9577), .Y(n10280) );
  AND2X1 U303 ( .A(n6246), .B(n6248), .Y(n5794) );
  AND2X1 U304 ( .A(n5448), .B(n6155), .Y(n5865) );
  AND2X1 U305 ( .A(n6243), .B(n24), .Y(n5769) );
  AND2X1 U306 ( .A(n4626), .B(n4712), .Y(n9932) );
  AND2X1 U307 ( .A(n4625), .B(n4690), .Y(n9931) );
  AND2X1 U308 ( .A(n4646), .B(n9846), .Y(n9915) );
  AND2X1 U309 ( .A(n46), .B(n6331), .Y(n9177) );
  AND2X1 U310 ( .A(n20), .B(n50), .Y(n5788) );
  AND2X1 U311 ( .A(n46), .B(n6231), .Y(n9114) );
  AND2X1 U312 ( .A(n46), .B(n6339), .Y(n9116) );
  AND2X1 U313 ( .A(n4642), .B(n4682), .Y(n9378) );
  AND2X1 U314 ( .A(n4624), .B(n4711), .Y(n8893) );
  AND2X1 U315 ( .A(n4623), .B(n4683), .Y(n8892) );
  AND2X1 U316 ( .A(n4640), .B(n9846), .Y(n8878) );
  AND2X1 U317 ( .A(n349), .B(n5666), .Y(n8479) );
  OR2X1 U318 ( .A(n6187), .B(n7581), .Y(n7869) );
  AND2X1 U319 ( .A(n4710), .B(n4677), .Y(n8252) );
  AND2X1 U320 ( .A(n8239), .B(n5519), .Y(n5756) );
  AND2X1 U321 ( .A(n4705), .B(n4653), .Y(n8447) );
  INVX1 U322 ( .A(oprB[39]), .Y(n6202) );
  AND2X1 U323 ( .A(n4622), .B(n4710), .Y(n7887) );
  INVX1 U324 ( .A(oprB[45]), .Y(n6190) );
  AND2X1 U325 ( .A(n4621), .B(n4675), .Y(n7886) );
  AND2X1 U326 ( .A(n271), .B(n5594), .Y(n7472) );
  AND2X1 U327 ( .A(n1959), .B(n3901), .Y(n7503) );
  AND2X1 U328 ( .A(n273), .B(n7497), .Y(n7502) );
  AND2X1 U329 ( .A(n274), .B(n1234), .Y(n7501) );
  AND2X1 U330 ( .A(n6173), .B(n5819), .Y(n5747) );
  AND2X1 U331 ( .A(n6551), .B(n67), .Y(n6966) );
  AND2X1 U332 ( .A(n4630), .B(n4670), .Y(n7214) );
  AND2X1 U333 ( .A(n4709), .B(n4669), .Y(n7238) );
  OR2X1 U334 ( .A(n6171), .B(n7141), .Y(n7405) );
  AND2X1 U335 ( .A(n4631), .B(n4666), .Y(n7352) );
  AND2X1 U336 ( .A(n2239), .B(n5838), .Y(n7109) );
  INVX1 U337 ( .A(oprB[55]), .Y(n6170) );
  AND2X1 U338 ( .A(n4620), .B(n4709), .Y(n6868) );
  AND2X1 U339 ( .A(n4619), .B(n4667), .Y(n6867) );
  AND2X1 U340 ( .A(n7224), .B(n5519), .Y(n5741) );
  AND2X1 U341 ( .A(n5720), .B(op[1]), .Y(n5878) );
  AND2X1 U342 ( .A(n1144), .B(n5208), .Y(n6638) );
  AND2X1 U343 ( .A(n4629), .B(n9846), .Y(n6853) );
  AND2X1 U344 ( .A(n5504), .B(n5732), .Y(n5736) );
  AND2X1 U345 ( .A(n186), .B(n1176), .Y(mult32_B[19]) );
  AND2X1 U346 ( .A(n79), .B(n91), .Y(mult32_B[13]) );
  AND2X1 U347 ( .A(n192), .B(n1179), .Y(mult32_B[15]) );
  AND2X1 U348 ( .A(n193), .B(n1181), .Y(mult32_B[12]) );
  AND2X1 U349 ( .A(n187), .B(n1177), .Y(mult32_B[18]) );
  AND2X1 U350 ( .A(n189), .B(n90), .Y(mult32_B[17]) );
  AND2X1 U351 ( .A(n1162), .B(n1497), .Y(mult32_A[27]) );
  AND2X1 U352 ( .A(n1161), .B(n1496), .Y(mult32_A[28]) );
  AND2X1 U353 ( .A(n181), .B(n1168), .Y(mult32_B[26]) );
  AND2X1 U354 ( .A(n182), .B(n1169), .Y(mult32_B[25]) );
  AND2X1 U355 ( .A(n183), .B(n1170), .Y(mult32_B[24]) );
  AND2X1 U356 ( .A(n184), .B(n1171), .Y(mult32_B[23]) );
  AND2X1 U357 ( .A(n76), .B(n1172), .Y(mult32_B[22]) );
  AND2X1 U358 ( .A(n77), .B(n1173), .Y(mult32_B[21]) );
  AND2X1 U359 ( .A(n185), .B(n1174), .Y(mult32_B[20]) );
  INVX1 U360 ( .A(n1531), .Y(n69) );
  AND2X1 U361 ( .A(n2838), .B(n6110), .Y(n10479) );
  AND2X1 U362 ( .A(n1134), .B(n94), .Y(n10321) );
  AND2X1 U363 ( .A(n1132), .B(n1482), .Y(n10287) );
  AND2X1 U364 ( .A(n5585), .B(n5586), .Y(n10226) );
  AND2X1 U365 ( .A(n999), .B(n1480), .Y(n10214) );
  AND2X1 U366 ( .A(n4649), .B(n4694), .Y(n10387) );
  AND2X1 U367 ( .A(n1160), .B(n1478), .Y(n10172) );
  AND2X1 U368 ( .A(n989), .B(n5424), .Y(n10079) );
  AND2X1 U369 ( .A(n983), .B(n1471), .Y(n10020) );
  AND2X1 U370 ( .A(n985), .B(n1473), .Y(n10042) );
  AND2X1 U371 ( .A(n977), .B(n1470), .Y(n9925) );
  OR2X1 U372 ( .A(n1965), .B(n6359), .Y(n9642) );
  INVX1 U373 ( .A(oprB[10]), .Y(n6252) );
  AND2X1 U374 ( .A(n969), .B(n1464), .Y(n9835) );
  INVX1 U375 ( .A(oprB[11]), .Y(n6250) );
  AND2X1 U376 ( .A(n6247), .B(n6245), .Y(n9792) );
  AND2X1 U377 ( .A(n965), .B(n1495), .Y(n9808) );
  AND2X1 U378 ( .A(n5800), .B(n6351), .Y(n9557) );
  AND2X1 U379 ( .A(n946), .B(n1451), .Y(n9561) );
  INVX1 U380 ( .A(oprB[16]), .Y(n6242) );
  AND2X1 U381 ( .A(n6232), .B(n5819), .Y(n9498) );
  AND2X1 U382 ( .A(n4639), .B(n4684), .Y(n9194) );
  AND2X1 U383 ( .A(n677), .B(n1446), .Y(n9339) );
  AND2X1 U384 ( .A(n670), .B(n1442), .Y(n9247) );
  AND2X1 U385 ( .A(n672), .B(n1493), .Y(n9278) );
  AND2X1 U386 ( .A(n665), .B(n1440), .Y(n9174) );
  AND2X1 U387 ( .A(n655), .B(n1434), .Y(n9043) );
  AND2X1 U388 ( .A(n651), .B(n1433), .Y(n9007) );
  AND2X1 U389 ( .A(n649), .B(n1431), .Y(n8986) );
  AND2X1 U390 ( .A(n642), .B(n1427), .Y(n8886) );
  OR2X1 U391 ( .A(n1964), .B(n6340), .Y(n8613) );
  INVX1 U392 ( .A(oprB[26]), .Y(n6225) );
  AND2X1 U393 ( .A(n634), .B(n1422), .Y(n8801) );
  INVX1 U394 ( .A(oprB[30]), .Y(n6218) );
  AND2X1 U395 ( .A(n355), .B(n1411), .Y(n8538) );
  AND2X1 U396 ( .A(n351), .B(n8502), .Y(n8507) );
  AND2X1 U397 ( .A(n352), .B(n1677), .Y(n8506) );
  AND2X1 U398 ( .A(n350), .B(n1409), .Y(n8489) );
  AND2X1 U399 ( .A(n340), .B(n1403), .Y(n8329) );
  AND2X1 U400 ( .A(n333), .B(n1399), .Y(n8235) );
  AND2X1 U401 ( .A(n328), .B(n1396), .Y(n8162) );
  AND2X1 U402 ( .A(n5653), .B(n5652), .Y(n8176) );
  AND2X1 U403 ( .A(n1152), .B(n1394), .Y(n8120) );
  AND2X1 U404 ( .A(n4636), .B(n4674), .Y(n8368) );
  AND2X1 U405 ( .A(n318), .B(n1389), .Y(n8032) );
  AND2X1 U406 ( .A(n315), .B(n1387), .Y(n7996) );
  AND2X1 U407 ( .A(n313), .B(n1257), .Y(n7974) );
  AND2X1 U408 ( .A(n307), .B(n1255), .Y(n7880) );
  OR2X1 U409 ( .A(n1963), .B(n6311), .Y(n7608) );
  AND2X1 U410 ( .A(n301), .B(n1251), .Y(n7817) );
  AND2X1 U411 ( .A(n299), .B(n1249), .Y(n7794) );
  AND2X1 U412 ( .A(n295), .B(n1491), .Y(n7767) );
  AND2X1 U413 ( .A(n82), .B(n7555), .Y(n7557) );
  AND2X1 U414 ( .A(n278), .B(n1236), .Y(n7534) );
  AND2X1 U415 ( .A(n262), .B(n1231), .Y(n7313) );
  AND2X1 U416 ( .A(n255), .B(n1225), .Y(n7218) );
  AND2X1 U417 ( .A(n6332), .B(n10502), .Y(n7189) );
  AND2X1 U418 ( .A(n253), .B(n1223), .Y(n7139) );
  AND2X1 U419 ( .A(n4632), .B(n4671), .Y(n7309) );
  AND2X1 U420 ( .A(n5640), .B(n6160), .Y(n5863) );
  AND2X1 U421 ( .A(n245), .B(n1219), .Y(n7019) );
  AND2X1 U422 ( .A(n242), .B(n1218), .Y(n6982) );
  AND2X1 U423 ( .A(n240), .B(n1216), .Y(n6958) );
  INVX1 U424 ( .A(op[3]), .Y(n6360) );
  AND2X1 U425 ( .A(n5820), .B(n67), .Y(n6925) );
  AND2X1 U426 ( .A(n234), .B(n1212), .Y(n6861) );
  AND2X1 U427 ( .A(n226), .B(n1206), .Y(n6772) );
  AND2X1 U428 ( .A(n206), .B(n1194), .Y(n6493) );
  INVX1 U429 ( .A(oprB[63]), .Y(n5891) );
  AND2X1 U430 ( .A(n195), .B(n1183), .Y(mult32_B[10]) );
  AND2X1 U431 ( .A(n200), .B(n1188), .Y(mult32_B[5]) );
  AND2X1 U432 ( .A(n81), .B(n1190), .Y(mult32_B[3]) );
  AND2X1 U433 ( .A(n78), .B(n1180), .Y(mult32_B[14]) );
  AND2X1 U434 ( .A(n201), .B(n1189), .Y(mult32_B[4]) );
  AND2X1 U435 ( .A(n5512), .B(n5511), .Y(mult32_A[31]) );
  AND2X1 U436 ( .A(n180), .B(n1167), .Y(mult32_B[27]) );
  AND2X1 U437 ( .A(n178), .B(n1165), .Y(mult32_B[29]) );
  INVX1 U438 ( .A(n439), .Y(n48) );
  INVX1 U439 ( .A(n5824), .Y(n13) );
  INVX1 U440 ( .A(n935), .Y(n12) );
  INVX1 U441 ( .A(oprB[2]), .Y(n6268) );
  INVX1 U442 ( .A(oprA[18]), .Y(n6017) );
  INVX1 U443 ( .A(oprB[3]), .Y(n6266) );
  AND2X1 U444 ( .A(n1139), .B(n1486), .Y(n10400) );
  AND2X1 U445 ( .A(n1955), .B(n4572), .Y(n10329) );
  AND2X1 U446 ( .A(n1135), .B(n1484), .Y(n10330) );
  AND2X1 U447 ( .A(n1133), .B(n1483), .Y(n10314) );
  OR2X1 U448 ( .A(n2061), .B(n2324), .Y(n10263) );
  AND2X1 U449 ( .A(n1001), .B(n5626), .Y(n10262) );
  OR2X1 U450 ( .A(n2085), .B(n2323), .Y(n10265) );
  AND2X1 U451 ( .A(n996), .B(n1479), .Y(n10188) );
  OR2X1 U452 ( .A(n2058), .B(n2320), .Y(n10192) );
  OR2X1 U453 ( .A(n2059), .B(n2321), .Y(n10191) );
  INVX1 U454 ( .A(n6007), .Y(n6331) );
  AND2X1 U455 ( .A(n992), .B(n1477), .Y(n10101) );
  AND2X1 U456 ( .A(n990), .B(n1475), .Y(n10098) );
  AND2X1 U457 ( .A(n993), .B(n5382), .Y(n10114) );
  AND2X1 U458 ( .A(n9967), .B(n1724), .Y(n9971) );
  OR2X1 U459 ( .A(n2054), .B(n2317), .Y(n10000) );
  OR2X1 U460 ( .A(n2053), .B(n2316), .Y(n10003) );
  AND2X1 U461 ( .A(n978), .B(n5619), .Y(n9936) );
  OR2X1 U462 ( .A(n2051), .B(n2314), .Y(n9938) );
  OR2X1 U463 ( .A(n2084), .B(n2313), .Y(n9939) );
  AND2X1 U464 ( .A(n975), .B(n1468), .Y(n9893) );
  AND2X1 U465 ( .A(n971), .B(n1466), .Y(n9860) );
  AND2X1 U466 ( .A(n970), .B(n1465), .Y(n9857) );
  AND2X1 U467 ( .A(n972), .B(n1467), .Y(n9870) );
  AND2X1 U468 ( .A(n966), .B(n1463), .Y(n9816) );
  AND2X1 U469 ( .A(n964), .B(n1462), .Y(n9801) );
  OR2X1 U470 ( .A(n2047), .B(n2308), .Y(n9748) );
  OR2X1 U471 ( .A(n2046), .B(n2307), .Y(n9750) );
  OR2X1 U472 ( .A(n2045), .B(n2338), .Y(n9751) );
  OR2X1 U473 ( .A(n2083), .B(n2304), .Y(n9672) );
  OR2X1 U474 ( .A(n2043), .B(n2305), .Y(n9670) );
  AND2X1 U475 ( .A(n958), .B(n1459), .Y(n9669) );
  OR2X1 U476 ( .A(n2082), .B(n2303), .Y(n9673) );
  AND2X1 U477 ( .A(n956), .B(n1457), .Y(n9624) );
  AND2X1 U478 ( .A(n949), .B(n1454), .Y(n9574) );
  AND2X1 U479 ( .A(n951), .B(n9582), .Y(n9584) );
  AND2X1 U480 ( .A(n952), .B(n1455), .Y(n9592) );
  AND2X1 U481 ( .A(n953), .B(n1456), .Y(n9591) );
  AND2X1 U482 ( .A(n947), .B(n1453), .Y(n9575) );
  AND2X1 U483 ( .A(n5363), .B(n5729), .Y(n10371) );
  AND2X1 U484 ( .A(n50), .B(n6231), .Y(n9310) );
  OR2X1 U485 ( .A(n2039), .B(n2301), .Y(n9412) );
  OR2X1 U486 ( .A(n2038), .B(n2299), .Y(n9414) );
  OR2X1 U487 ( .A(n2037), .B(n2298), .Y(n9415) );
  OR2X1 U488 ( .A(n2081), .B(n113), .Y(n9351) );
  AND2X1 U489 ( .A(n676), .B(n1445), .Y(n9308) );
  AND2X1 U490 ( .A(n678), .B(n1447), .Y(n9348) );
  OR2X1 U491 ( .A(n2035), .B(n114), .Y(n9350) );
  AND2X1 U492 ( .A(n673), .B(n1444), .Y(n9286) );
  AND2X1 U493 ( .A(n671), .B(n1443), .Y(n9272) );
  OR2X1 U494 ( .A(n2032), .B(n2165), .Y(n9223) );
  AND2X1 U495 ( .A(n667), .B(n5692), .Y(n9222) );
  OR2X1 U496 ( .A(n2080), .B(n2164), .Y(n9225) );
  INVX1 U497 ( .A(oprA[5]), .Y(n6349) );
  AND2X1 U498 ( .A(n662), .B(n1439), .Y(n9148) );
  AND2X1 U499 ( .A(n1156), .B(n1438), .Y(n9132) );
  OR2X1 U500 ( .A(n2030), .B(n2162), .Y(n9151) );
  OR2X1 U501 ( .A(n2029), .B(n2161), .Y(n9152) );
  AND2X1 U502 ( .A(n656), .B(n1435), .Y(n9059) );
  AND2X1 U503 ( .A(n659), .B(n5618), .Y(n9074) );
  AND2X1 U504 ( .A(n658), .B(n1437), .Y(n9062) );
  AND2X1 U505 ( .A(n650), .B(n1432), .Y(n9004) );
  AND2X1 U506 ( .A(n652), .B(n5551), .Y(n9017) );
  AND2X1 U507 ( .A(n5509), .B(n6155), .Y(n5860) );
  AND2X1 U508 ( .A(n5267), .B(n6218), .Y(n8610) );
  AND2X1 U509 ( .A(n6219), .B(n6221), .Y(n5798) );
  AND2X1 U510 ( .A(n643), .B(n1428), .Y(n8897) );
  OR2X1 U511 ( .A(n2025), .B(n2157), .Y(n8899) );
  OR2X1 U512 ( .A(n2079), .B(n2156), .Y(n8900) );
  AND2X1 U513 ( .A(n640), .B(n1425), .Y(n8857) );
  AND2X1 U514 ( .A(n636), .B(n1424), .Y(n8824) );
  AND2X1 U515 ( .A(n635), .B(n1423), .Y(n8821) );
  AND2X1 U516 ( .A(n637), .B(n5377), .Y(n8834) );
  AND2X1 U517 ( .A(n630), .B(n1492), .Y(n8774) );
  AND2X1 U518 ( .A(n631), .B(n5438), .Y(n8782) );
  AND2X1 U519 ( .A(n629), .B(n1421), .Y(n8768) );
  AND2X1 U520 ( .A(n5908), .B(n6221), .Y(n9127) );
  AND2X1 U521 ( .A(n5267), .B(n6217), .Y(n8588) );
  INVX1 U522 ( .A(oprB[28]), .Y(n6221) );
  OR2X1 U523 ( .A(n2078), .B(n2151), .Y(n8642) );
  OR2X1 U524 ( .A(n2021), .B(n2152), .Y(n8640) );
  OR2X1 U525 ( .A(n2077), .B(n2150), .Y(n8643) );
  AND2X1 U526 ( .A(n359), .B(n8559), .Y(n8561) );
  AND2X1 U527 ( .A(n356), .B(n1413), .Y(n8552) );
  AND2X1 U528 ( .A(n358), .B(n1414), .Y(n8551) );
  BUFX2 U529 ( .A(n5284), .Y(n5266) );
  AND2X1 U530 ( .A(n346), .B(n1407), .Y(n8452) );
  OR2X1 U531 ( .A(n2018), .B(n2148), .Y(n8453) );
  OR2X1 U532 ( .A(n2076), .B(n2147), .Y(n8432) );
  AND2X1 U533 ( .A(n345), .B(n1406), .Y(n8431) );
  OR2X1 U534 ( .A(n4452), .B(n8399), .Y(n4454) );
  AND2X1 U535 ( .A(n341), .B(n1404), .Y(n8338) );
  AND2X1 U536 ( .A(n335), .B(n92), .Y(n8267) );
  AND2X1 U537 ( .A(n336), .B(n1401), .Y(n8275) );
  AND2X1 U538 ( .A(n334), .B(n1400), .Y(n8261) );
  OR2X1 U539 ( .A(n101), .B(n2138), .Y(n8211) );
  AND2X1 U540 ( .A(n330), .B(n1398), .Y(n8210) );
  OR2X1 U541 ( .A(n2074), .B(n2137), .Y(n8213) );
  AND2X1 U542 ( .A(n325), .B(n1395), .Y(n8136) );
  OR2X1 U543 ( .A(n2012), .B(n2135), .Y(n8139) );
  OR2X1 U544 ( .A(n2011), .B(n2134), .Y(n8140) );
  AND2X1 U545 ( .A(n321), .B(n1392), .Y(n8051) );
  AND2X1 U546 ( .A(n319), .B(n1390), .Y(n8048) );
  AND2X1 U547 ( .A(n322), .B(n1393), .Y(n8063) );
  AND2X1 U548 ( .A(n7922), .B(n1661), .Y(n7925) );
  OR2X1 U549 ( .A(n2007), .B(n2131), .Y(n7954) );
  OR2X1 U550 ( .A(n2006), .B(n2130), .Y(n7957) );
  AND2X1 U551 ( .A(n308), .B(n1256), .Y(n7891) );
  OR2X1 U552 ( .A(n2004), .B(n2128), .Y(n7893) );
  OR2X1 U553 ( .A(n2073), .B(n2127), .Y(n7894) );
  AND2X1 U554 ( .A(n305), .B(n1253), .Y(n7849) );
  AND2X1 U555 ( .A(n300), .B(n1250), .Y(n7814) );
  AND2X1 U556 ( .A(n302), .B(n1252), .Y(n7827) );
  AND2X1 U557 ( .A(n296), .B(n1248), .Y(n7775) );
  AND2X1 U558 ( .A(n294), .B(n1247), .Y(n7761) );
  OR2X1 U559 ( .A(n2000), .B(n2122), .Y(n7713) );
  OR2X1 U560 ( .A(n1999), .B(n2121), .Y(n7715) );
  OR2X1 U561 ( .A(n1998), .B(n2336), .Y(n7716) );
  OR2X1 U562 ( .A(n2072), .B(n2118), .Y(n7640) );
  OR2X1 U563 ( .A(n1996), .B(n2119), .Y(n7638) );
  AND2X1 U564 ( .A(n288), .B(n1244), .Y(n7637) );
  OR2X1 U565 ( .A(n2071), .B(n2117), .Y(n7641) );
  AND2X1 U566 ( .A(n286), .B(n1242), .Y(n7596) );
  AND2X1 U567 ( .A(n282), .B(n1240), .Y(n7565) );
  AND2X1 U568 ( .A(n283), .B(n1241), .Y(n7564) );
  AND2X1 U569 ( .A(n279), .B(n1238), .Y(n7548) );
  AND2X1 U570 ( .A(n281), .B(n1239), .Y(n7547) );
  INVX1 U571 ( .A(n1065), .Y(n31) );
  OR2X1 U572 ( .A(n1990), .B(n2113), .Y(n7389) );
  OR2X1 U573 ( .A(n1989), .B(n2112), .Y(n7390) );
  OR2X1 U574 ( .A(n2070), .B(n2109), .Y(n7325) );
  AND2X1 U575 ( .A(n261), .B(n1230), .Y(n7283) );
  OR2X1 U576 ( .A(n1987), .B(n2110), .Y(n7324) );
  AND2X1 U577 ( .A(n263), .B(n1232), .Y(n7322) );
  AND2X1 U578 ( .A(n258), .B(n1229), .Y(n7260) );
  AND2X1 U579 ( .A(n256), .B(n1227), .Y(n7247) );
  AND2X1 U580 ( .A(n257), .B(n1228), .Y(n7250) );
  OR2X1 U581 ( .A(n1984), .B(n2106), .Y(n7194) );
  OR2X1 U582 ( .A(n1983), .B(n2105), .Y(n7196) );
  OR2X1 U583 ( .A(n1980), .B(n2102), .Y(n7121) );
  OR2X1 U584 ( .A(n1981), .B(n2103), .Y(n7119) );
  AND2X1 U585 ( .A(n248), .B(n1222), .Y(n7038) );
  AND2X1 U586 ( .A(n246), .B(n1220), .Y(n7035) );
  AND2X1 U587 ( .A(n249), .B(n5540), .Y(n7050) );
  AND2X1 U588 ( .A(n241), .B(n1217), .Y(n6979) );
  INVX1 U589 ( .A(oprA[40]), .Y(n6298) );
  AND2X1 U590 ( .A(n5721), .B(n5012), .Y(n5739) );
  AND2X1 U591 ( .A(n6160), .B(n6161), .Y(n5841) );
  AND2X1 U592 ( .A(n5897), .B(n5892), .Y(n6551) );
  AND2X1 U593 ( .A(n235), .B(n1213), .Y(n6872) );
  OR2X1 U594 ( .A(n1976), .B(n2098), .Y(n6874) );
  OR2X1 U595 ( .A(n2069), .B(n2097), .Y(n6875) );
  AND2X1 U596 ( .A(n228), .B(n1208), .Y(n6798) );
  AND2X1 U597 ( .A(n227), .B(n1207), .Y(n6795) );
  AND2X1 U598 ( .A(n229), .B(n1209), .Y(n6808) );
  INVX1 U599 ( .A(oprA[43]), .Y(n5962) );
  AND2X1 U600 ( .A(n222), .B(n1488), .Y(n6745) );
  AND2X1 U601 ( .A(n223), .B(n5389), .Y(n6754) );
  AND2X1 U602 ( .A(n221), .B(n1205), .Y(n6739) );
  OR2X1 U603 ( .A(n1972), .B(n2093), .Y(n6685) );
  OR2X1 U604 ( .A(n1971), .B(n2092), .Y(n6687) );
  OR2X1 U605 ( .A(n1970), .B(n2335), .Y(n6688) );
  AND2X1 U606 ( .A(n1145), .B(n1203), .Y(n6647) );
  OR2X1 U607 ( .A(n2068), .B(n2089), .Y(n6609) );
  OR2X1 U608 ( .A(n1968), .B(n2090), .Y(n6607) );
  OR2X1 U609 ( .A(n2067), .B(n2088), .Y(n6610) );
  AND2X1 U610 ( .A(n210), .B(n6522), .Y(n6524) );
  AND2X1 U611 ( .A(n209), .B(n1197), .Y(n6513) );
  AND2X1 U612 ( .A(n207), .B(n1196), .Y(n6514) );
  AND2X1 U613 ( .A(n203), .B(n1192), .Y(mult32_B[1]) );
  AND2X1 U614 ( .A(n202), .B(n1191), .Y(mult32_B[2]) );
  AND2X1 U615 ( .A(n179), .B(n1166), .Y(mult32_B[28]) );
  INVX1 U616 ( .A(oprB[0]), .Y(n6272) );
  INVX1 U617 ( .A(oprB[1]), .Y(n6270) );
  OR2X1 U618 ( .A(n2065), .B(n2331), .Y(n10470) );
  OR2X1 U619 ( .A(n10458), .B(n2333), .Y(n10467) );
  OR2X1 U620 ( .A(n2066), .B(n2332), .Y(n10469) );
  OR2X1 U621 ( .A(n5468), .B(n2329), .Y(n10403) );
  OR2X1 U622 ( .A(n2064), .B(n2330), .Y(n10402) );
  AND2X1 U623 ( .A(n10054), .B(n10053), .Y(n10055) );
  OR2X1 U624 ( .A(n20), .B(n9170), .Y(n9474) );
  AND2X1 U625 ( .A(n10290), .B(n6233), .Y(n9168) );
  AND2X1 U626 ( .A(n939), .B(n1705), .Y(n9438) );
  AND2X1 U627 ( .A(n616), .B(n1415), .Y(n8569) );
  AND2X1 U628 ( .A(n617), .B(n1416), .Y(n8568) );
  INVX1 U629 ( .A(oprB[33]), .Y(n6214) );
  OR2X1 U630 ( .A(n2016), .B(n2144), .Y(n8404) );
  OR2X1 U631 ( .A(n2017), .B(n2145), .Y(n8403) );
  OR2X1 U632 ( .A(n102), .B(n2141), .Y(n8340) );
  OR2X1 U633 ( .A(n2075), .B(n2140), .Y(n8341) );
  AND2X1 U634 ( .A(n8008), .B(n8007), .Y(n8009) );
  BUFX2 U635 ( .A(n5921), .Y(n17) );
  AND2X1 U636 ( .A(n211), .B(n1198), .Y(n6532) );
  AND2X1 U637 ( .A(n212), .B(n1199), .Y(n6531) );
  AND2X1 U638 ( .A(n177), .B(n1164), .Y(mult32_B[30]) );
  AND2X1 U639 ( .A(n6142), .B(n150), .Y(n10549) );
  AND2X1 U640 ( .A(n83), .B(n1708), .Y(n9470) );
  AND2X1 U641 ( .A(n9467), .B(n1707), .Y(n9482) );
  AND2X1 U642 ( .A(n1961), .B(n4054), .Y(n9435) );
  AND2X1 U643 ( .A(n938), .B(n1448), .Y(n9433) );
  AND2X1 U644 ( .A(n940), .B(n1706), .Y(n9450) );
  AND2X1 U645 ( .A(n5478), .B(n8923), .Y(n8925) );
  AND2X1 U646 ( .A(n647), .B(n1430), .Y(n8932) );
  AND2X1 U647 ( .A(n5687), .B(n1689), .Y(n8933) );
  AND2X1 U648 ( .A(n8958), .B(n1690), .Y(n8974) );
  AND2X1 U649 ( .A(n5525), .B(n5524), .Y(n8961) );
  AND2X1 U650 ( .A(n645), .B(n1688), .Y(n8920) );
  AND2X1 U651 ( .A(n646), .B(n1429), .Y(n8919) );
  AND2X1 U652 ( .A(n624), .B(n8665), .Y(n8667) );
  AND2X1 U653 ( .A(n625), .B(n5668), .Y(n8674) );
  AND2X1 U654 ( .A(n5490), .B(n1680), .Y(n8675) );
  AND2X1 U655 ( .A(n622), .B(n5667), .Y(n8662) );
  AND2X1 U656 ( .A(n623), .B(n5554), .Y(n8661) );
  AND2X1 U657 ( .A(n626), .B(n5495), .Y(n8712) );
  AND2X1 U658 ( .A(n1163), .B(n1681), .Y(n8726) );
  AND2X1 U659 ( .A(n5421), .B(n6897), .Y(n6899) );
  AND2X1 U660 ( .A(n239), .B(n1215), .Y(n6906) );
  AND2X1 U661 ( .A(n5620), .B(n1509), .Y(n6907) );
  AND2X1 U662 ( .A(n6931), .B(n1510), .Y(n6946) );
  AND2X1 U663 ( .A(n5366), .B(n5365), .Y(n6934) );
  AND2X1 U664 ( .A(n237), .B(n1508), .Y(n6894) );
  AND2X1 U665 ( .A(n238), .B(n1214), .Y(n6893) );
  AND2X1 U666 ( .A(n1141), .B(n1738), .Y(n10474) );
  AND2X1 U667 ( .A(n943), .B(n1710), .Y(n9539) );
  AND2X1 U668 ( .A(n942), .B(n1709), .Y(n9489) );
  AND2X1 U669 ( .A(n937), .B(n1704), .Y(n9419) );
  AND2X1 U670 ( .A(n680), .B(n1703), .Y(n9362) );
  AND2X1 U671 ( .A(n8517), .B(n95), .Y(n8519) );
  INVX1 U672 ( .A(n8467), .Y(n63) );
  AND2X1 U673 ( .A(n343), .B(n1675), .Y(n8408) );
  AND2X1 U674 ( .A(n5463), .B(n5464), .Y(n8352) );
  AND2X1 U675 ( .A(n266), .B(n1613), .Y(n7394) );
  AND2X1 U676 ( .A(n265), .B(n1581), .Y(n7336) );
  OR2X1 U677 ( .A(n2063), .B(n118), .Y(result[3]) );
  OR2X1 U678 ( .A(n2062), .B(n2328), .Y(result[4]) );
  OR2X1 U679 ( .A(n2060), .B(n2326), .Y(result[5]) );
  OR2X1 U680 ( .A(n2057), .B(n2322), .Y(result[6]) );
  OR2X1 U681 ( .A(n2056), .B(n2319), .Y(result[7]) );
  OR2X1 U682 ( .A(n2055), .B(n117), .Y(result[8]) );
  OR2X1 U683 ( .A(n2052), .B(n2318), .Y(result[9]) );
  OR2X1 U684 ( .A(n2050), .B(n2315), .Y(result[10]) );
  OR2X1 U685 ( .A(n2049), .B(n2312), .Y(result[11]) );
  OR2X1 U686 ( .A(n2048), .B(n2310), .Y(result[12]) );
  OR2X1 U687 ( .A(n2044), .B(n2309), .Y(result[13]) );
  OR2X1 U688 ( .A(n2042), .B(n2306), .Y(result[14]) );
  OR2X1 U689 ( .A(n2041), .B(n2302), .Y(result[15]) );
  AND2X1 U690 ( .A(n87), .B(n6141), .Y(result[17]) );
  OR2X1 U691 ( .A(n2034), .B(n2297), .Y(result[19]) );
  OR2X1 U692 ( .A(n2033), .B(n2296), .Y(result[20]) );
  OR2X1 U693 ( .A(n2031), .B(n2294), .Y(result[21]) );
  OR2X1 U694 ( .A(n2028), .B(n2163), .Y(result[22]) );
  OR2X1 U695 ( .A(n2027), .B(n2160), .Y(result[23]) );
  OR2X1 U696 ( .A(n2026), .B(n2159), .Y(result[24]) );
  AND2X1 U697 ( .A(n1154), .B(n6141), .Y(result[25]) );
  OR2X1 U698 ( .A(n2024), .B(n2158), .Y(result[26]) );
  OR2X1 U699 ( .A(n2023), .B(n2155), .Y(result[27]) );
  OR2X1 U700 ( .A(n2022), .B(n2154), .Y(result[28]) );
  AND2X1 U701 ( .A(n1153), .B(n6141), .Y(result[29]) );
  OR2X1 U702 ( .A(n2020), .B(n2153), .Y(result[30]) );
  OR2X1 U703 ( .A(n2019), .B(n2149), .Y(result[31]) );
  OR2X1 U704 ( .A(n2015), .B(n2143), .Y(result[35]) );
  OR2X1 U705 ( .A(n2014), .B(n111), .Y(result[36]) );
  OR2X1 U706 ( .A(n2013), .B(n2139), .Y(result[37]) );
  OR2X1 U707 ( .A(n2010), .B(n2136), .Y(result[38]) );
  OR2X1 U708 ( .A(n2009), .B(n2133), .Y(result[39]) );
  OR2X1 U709 ( .A(n2008), .B(n110), .Y(result[40]) );
  OR2X1 U710 ( .A(n2005), .B(n2132), .Y(result[41]) );
  OR2X1 U711 ( .A(n2003), .B(n2129), .Y(result[42]) );
  OR2X1 U712 ( .A(n2002), .B(n2126), .Y(result[43]) );
  OR2X1 U713 ( .A(n2001), .B(n2124), .Y(result[44]) );
  OR2X1 U714 ( .A(n1997), .B(n2123), .Y(result[45]) );
  OR2X1 U715 ( .A(n1995), .B(n2120), .Y(result[46]) );
  OR2X1 U716 ( .A(n1994), .B(n2116), .Y(result[47]) );
  OR2X1 U717 ( .A(n1993), .B(n109), .Y(result[48]) );
  OR2X1 U718 ( .A(n1992), .B(n108), .Y(result[49]) );
  OR2X1 U719 ( .A(n1986), .B(n2111), .Y(result[51]) );
  OR2X1 U720 ( .A(n1985), .B(n2108), .Y(result[52]) );
  OR2X1 U721 ( .A(n1982), .B(n2107), .Y(result[53]) );
  OR2X1 U722 ( .A(n1979), .B(n2104), .Y(result[54]) );
  OR2X1 U723 ( .A(n1978), .B(n2101), .Y(result[55]) );
  OR2X1 U724 ( .A(n1977), .B(n2100), .Y(result[56]) );
  AND2X1 U725 ( .A(n1146), .B(n6141), .Y(result[57]) );
  OR2X1 U726 ( .A(n1975), .B(n2099), .Y(result[58]) );
  OR2X1 U727 ( .A(n1974), .B(n2096), .Y(result[59]) );
  OR2X1 U728 ( .A(n1973), .B(n2095), .Y(result[60]) );
  OR2X1 U729 ( .A(n1969), .B(n2094), .Y(result[61]) );
  OR2X1 U730 ( .A(n1967), .B(n2091), .Y(result[62]) );
  OR2X1 U731 ( .A(n1966), .B(n2087), .Y(result[63]) );
  AND2X2 U732 ( .A(n8554), .B(n5991), .Y(n5740) );
  AND2X2 U733 ( .A(n5991), .B(n9632), .Y(n8592) );
  INVX2 U734 ( .A(n6283), .Y(n5929) );
  INVX2 U735 ( .A(n5278), .Y(n6014) );
  INVX1 U736 ( .A(n6331), .Y(n10) );
  BUFX4 U737 ( .A(oprB[31]), .Y(n5284) );
  OAI21X1 U738 ( .A(n12), .B(n13), .C(n14), .Y(n11) );
  INVX1 U739 ( .A(n11), .Y(n10544) );
  INVX1 U740 ( .A(n10543), .Y(n14) );
  INVX4 U741 ( .A(oprA[2]), .Y(n6355) );
  INVX1 U742 ( .A(shift_amount[4]), .Y(n6152) );
  BUFX2 U743 ( .A(oprB[13]), .Y(n15) );
  BUFX2 U744 ( .A(oprB[15]), .Y(n23) );
  INVX4 U745 ( .A(oprA[4]), .Y(n6352) );
  INVX4 U746 ( .A(n6333), .Y(n6008) );
  INVX1 U747 ( .A(oprA[20]), .Y(n6010) );
  AND2X1 U748 ( .A(n936), .B(n6133), .Y(n10604) );
  INVX1 U749 ( .A(n5913), .Y(n5916) );
  INVX8 U750 ( .A(n65), .Y(n67) );
  BUFX2 U751 ( .A(n6230), .Y(n18) );
  BUFX2 U752 ( .A(n6230), .Y(n19) );
  BUFX2 U753 ( .A(n6230), .Y(n20) );
  INVX1 U754 ( .A(n6231), .Y(n6230) );
  BUFX2 U755 ( .A(n6047), .Y(n21) );
  INVX4 U756 ( .A(n6227), .Y(n6226) );
  INVX1 U757 ( .A(oprB[25]), .Y(n6227) );
  INVX8 U758 ( .A(n5923), .Y(n5925) );
  AND2X1 U759 ( .A(n6158), .B(n6159), .Y(n6517) );
  AND2X1 U760 ( .A(n6243), .B(n70), .Y(n9614) );
  INVX2 U761 ( .A(n72), .Y(n6319) );
  AND2X1 U762 ( .A(n70), .B(n6244), .Y(n9639) );
  INVX1 U763 ( .A(oprB[61]), .Y(n6160) );
  INVX1 U764 ( .A(oprA[50]), .Y(n5943) );
  AND2X1 U765 ( .A(n9), .B(n6159), .Y(n6579) );
  AND2X1 U766 ( .A(n7222), .B(n5451), .Y(n6791) );
  AND2X1 U767 ( .A(n8811), .B(n5908), .Y(n9046) );
  INVX1 U768 ( .A(n5998), .Y(n5996) );
  INVX1 U769 ( .A(oprA[12]), .Y(n6030) );
  AND2X1 U770 ( .A(n5819), .B(n51), .Y(n10356) );
  AND2X1 U771 ( .A(n10290), .B(n51), .Y(n10208) );
  AND2X1 U772 ( .A(n5562), .B(n5393), .Y(n6071) );
  INVX1 U773 ( .A(oprA[42]), .Y(n6295) );
  AND2X1 U774 ( .A(n6257), .B(n6260), .Y(n10154) );
  INVX1 U775 ( .A(oprA[36]), .Y(n5979) );
  INVX1 U776 ( .A(oprA[44]), .Y(n5959) );
  AND2X1 U777 ( .A(n5819), .B(n6174), .Y(n7285) );
  INVX2 U778 ( .A(oprA[32]), .Y(n6311) );
  AND2X1 U779 ( .A(n306), .B(n1254), .Y(n8127) );
  AND2X1 U780 ( .A(n233), .B(n1211), .Y(n7089) );
  INVX2 U781 ( .A(oprA[14]), .Y(n6341) );
  INVX1 U782 ( .A(n6), .Y(n6048) );
  INVX1 U783 ( .A(oprA[52]), .Y(n5939) );
  INVX2 U784 ( .A(n6017), .Y(n6019) );
  AND2X1 U785 ( .A(n6247), .B(n6246), .Y(n10034) );
  INVX2 U786 ( .A(n6285), .Y(n5934) );
  INVX1 U787 ( .A(oprA[24]), .Y(n6002) );
  INVX1 U788 ( .A(oprA[55]), .Y(n5930) );
  AND2X1 U789 ( .A(n6261), .B(n5819), .Y(n10498) );
  AND2X1 U790 ( .A(n976), .B(n1469), .Y(n10179) );
  AND2X1 U791 ( .A(n641), .B(n1426), .Y(n9139) );
  INVX2 U792 ( .A(n5959), .Y(n5961) );
  INVX2 U793 ( .A(n5962), .Y(n5964) );
  AND2X1 U794 ( .A(n7224), .B(n1226), .Y(n8239) );
  AND2X1 U795 ( .A(n247), .B(n1221), .Y(n7308) );
  AND2X1 U796 ( .A(n320), .B(n1391), .Y(n8324) );
  AND2X1 U797 ( .A(n657), .B(n1436), .Y(n9334) );
  AND2X1 U798 ( .A(n991), .B(n1476), .Y(n10386) );
  AND2X1 U799 ( .A(n1151), .B(n5732), .Y(n8497) );
  AND2X1 U800 ( .A(n9310), .B(n6011), .Y(n9266) );
  AND2X1 U801 ( .A(n8554), .B(n6315), .Y(n8701) );
  AND2X1 U802 ( .A(n8610), .B(n6334), .Y(n8685) );
  AND2X1 U803 ( .A(n8554), .B(n6011), .Y(n9240) );
  AND2X1 U804 ( .A(n6011), .B(n9688), .Y(n9260) );
  AND2X1 U805 ( .A(n6043), .B(n9577), .Y(n10073) );
  AND2X1 U806 ( .A(n5821), .B(n6221), .Y(n8811) );
  AND2X1 U807 ( .A(n5720), .B(n5870), .Y(n5818) );
  AND2X1 U808 ( .A(n6247), .B(n5821), .Y(n10424) );
  AND2X1 U809 ( .A(n6655), .B(n6159), .Y(n6662) );
  AND2X1 U810 ( .A(n8703), .B(n6218), .Y(n8717) );
  AND2X1 U811 ( .A(n44), .B(n9688), .Y(n8805) );
  AND2X1 U812 ( .A(n6085), .B(n5504), .Y(n9803) );
  AND2X1 U813 ( .A(n6171), .B(n6169), .Y(n7167) );
  INVX1 U814 ( .A(oprA[38]), .Y(n6300) );
  INVX2 U815 ( .A(oprA[48]), .Y(n6292) );
  AND2X1 U816 ( .A(n10291), .B(n51), .Y(n10436) );
  INVX1 U817 ( .A(oprA[56]), .Y(n6283) );
  INVX1 U818 ( .A(oprA[60]), .Y(n6276) );
  INVX1 U819 ( .A(oprA[16]), .Y(n6340) );
  AND2X1 U820 ( .A(n5392), .B(n5440), .Y(n6457) );
  OR2X1 U821 ( .A(n4387), .B(n4388), .Y(n4385) );
  INVX1 U822 ( .A(n6338), .Y(n6337) );
  AND2X1 U823 ( .A(n9996), .B(n6246), .Y(n10486) );
  AND2X1 U824 ( .A(n1147), .B(n5732), .Y(n7492) );
  AND2X1 U825 ( .A(n1155), .B(n5732), .Y(n9509) );
  AND2X1 U826 ( .A(n1159), .B(n5732), .Y(n10556) );
  AND2X1 U827 ( .A(n6011), .B(n5800), .Y(n8534) );
  AND2X1 U828 ( .A(n5581), .B(n5580), .Y(n9187) );
  AND2X1 U829 ( .A(n8610), .B(n5992), .Y(n8677) );
  AND2X1 U830 ( .A(n6579), .B(n5916), .Y(n6628) );
  AND2X1 U831 ( .A(n8610), .B(n6315), .Y(n8754) );
  AND2X1 U832 ( .A(n1956), .B(n1948), .Y(n4577) );
  OR2X1 U833 ( .A(n4160), .B(n7823), .Y(n4162) );
  OR2X1 U834 ( .A(n4168), .B(n8002), .Y(n4170) );
  OR2X1 U835 ( .A(n4217), .B(n10048), .Y(n4219) );
  AND2X1 U836 ( .A(n5430), .B(n1946), .Y(n4054) );
  AND2X1 U837 ( .A(n4707), .B(n4659), .Y(n10499) );
  INVX1 U838 ( .A(oprA[9]), .Y(n6344) );
  INVX2 U839 ( .A(n6317), .Y(n26) );
  INVX1 U840 ( .A(oprA[8]), .Y(n6346) );
  OR2X1 U841 ( .A(n4161), .B(n4162), .Y(n4159) );
  OR2X1 U842 ( .A(n4169), .B(n4170), .Y(n4167) );
  OR2X1 U843 ( .A(n4218), .B(n4219), .Y(n4216) );
  AND2X1 U844 ( .A(n5834), .B(n5451), .Y(n8968) );
  AND2X1 U845 ( .A(n5833), .B(n5451), .Y(n9774) );
  AND2X1 U846 ( .A(n220), .B(n1204), .Y(n7475) );
  INVX1 U847 ( .A(oprA[45]), .Y(n6294) );
  INVX1 U848 ( .A(oprA[46]), .Y(n6293) );
  INVX2 U849 ( .A(oprA[34]), .Y(n6307) );
  AND2X1 U850 ( .A(n6245), .B(n6248), .Y(n10167) );
  INVX2 U851 ( .A(oprA[53]), .Y(n5936) );
  AND2X1 U852 ( .A(n10355), .B(n6), .Y(n10217) );
  AND2X1 U853 ( .A(n6029), .B(n9614), .Y(n9912) );
  AND2X1 U854 ( .A(n5800), .B(n6026), .Y(n9840) );
  AND2X1 U855 ( .A(n6334), .B(n6081), .Y(n8617) );
  AND2X1 U856 ( .A(n9626), .B(n6351), .Y(n9646) );
  AND2X1 U857 ( .A(n5915), .B(n6080), .Y(n6777) );
  AND2X1 U858 ( .A(n5992), .B(n6080), .Y(n8806) );
  BUFX2 U859 ( .A(oprA[28]), .Y(n5275) );
  INVX2 U860 ( .A(oprA[61]), .Y(n6274) );
  INVX1 U861 ( .A(oprA[54]), .Y(n6285) );
  AND2X1 U862 ( .A(n6658), .B(n6159), .Y(n6913) );
  AND2X1 U863 ( .A(n9721), .B(n6244), .Y(n9996) );
  INVX1 U864 ( .A(oprA[37]), .Y(n6302) );
  AND2X1 U865 ( .A(n9688), .B(n5936), .Y(n7157) );
  AND2X1 U866 ( .A(n9688), .B(n6333), .Y(n9199) );
  AND2X1 U867 ( .A(n9688), .B(n6), .Y(n10238) );
  INVX1 U868 ( .A(oprA[9]), .Y(n6036) );
  OR2X1 U869 ( .A(n3910), .B(n3911), .Y(n3907) );
  OR2X1 U870 ( .A(n4047), .B(n4048), .Y(n4044) );
  OR2X1 U871 ( .A(n4210), .B(n4211), .Y(n4208) );
  AND2X1 U872 ( .A(n5574), .B(n5364), .Y(n5766) );
  AND2X1 U873 ( .A(n5907), .B(n7491), .Y(n9324) );
  AND2X1 U874 ( .A(n4706), .B(n4656), .Y(n9475) );
  AND2X1 U875 ( .A(n5516), .B(n5517), .Y(n7148) );
  AND2X1 U876 ( .A(n45), .B(n6065), .Y(n7759) );
  AND2X1 U877 ( .A(n293), .B(n1246), .Y(n8482) );
  AND2X1 U878 ( .A(n8692), .B(n6218), .Y(n8939) );
  AND2X1 U879 ( .A(n5587), .B(n4665), .Y(n5801) );
  INVX1 U880 ( .A(n6233), .Y(n22) );
  INVX2 U881 ( .A(oprB[21]), .Y(n6233) );
  INVX8 U882 ( .A(n6314), .Y(n5994) );
  INVX8 U883 ( .A(n6311), .Y(n5988) );
  AND2X2 U884 ( .A(n6205), .B(n5988), .Y(n5761) );
  INVX4 U885 ( .A(n6307), .Y(n5983) );
  INVX2 U886 ( .A(oprB[34]), .Y(n6212) );
  INVX4 U887 ( .A(n6005), .Y(n6006) );
  INVX8 U888 ( .A(n5881), .Y(n59) );
  INVX1 U889 ( .A(n70), .Y(n24) );
  INVX2 U890 ( .A(n6208), .Y(n6207) );
  INVX1 U891 ( .A(oprB[23]), .Y(n25) );
  INVX8 U892 ( .A(n6172), .Y(n6171) );
  INVX1 U893 ( .A(n6010), .Y(n6334) );
  INVX8 U894 ( .A(n26), .Y(n27) );
  INVX1 U895 ( .A(oprB[53]), .Y(n6174) );
  INVX8 U896 ( .A(n6174), .Y(n6173) );
  INVX1 U897 ( .A(n28), .Y(n33) );
  INVX1 U898 ( .A(n6010), .Y(n6013) );
  BUFX2 U899 ( .A(n10603), .Y(n28) );
  INVX8 U900 ( .A(n65), .Y(n66) );
  INVX4 U901 ( .A(n6030), .Y(n6032) );
  INVX1 U902 ( .A(oprA[1]), .Y(n6357) );
  INVX4 U903 ( .A(oprB[60]), .Y(n6161) );
  INVX2 U904 ( .A(n6352), .Y(n6350) );
  INVX8 U905 ( .A(n6180), .Y(n6179) );
  INVX2 U906 ( .A(n6027), .Y(n6029) );
  INVX8 U907 ( .A(n6005), .Y(n6007) );
  INVX8 U908 ( .A(n6329), .Y(n6328) );
  OAI21X1 U909 ( .A(n31), .B(n6130), .C(n7506), .Y(n30) );
  AND2X1 U910 ( .A(n7505), .B(n7504), .Y(n7506) );
  INVX1 U911 ( .A(n32), .Y(n10605) );
  INVX4 U912 ( .A(n5930), .Y(n5932) );
  INVX4 U913 ( .A(n5930), .Y(n5931) );
  INVX8 U914 ( .A(n6313), .Y(n5993) );
  NOR3X1 U915 ( .A(n10604), .B(n47), .C(n33), .Y(n32) );
  INVX2 U916 ( .A(n5898), .Y(n5900) );
  OAI21X1 U917 ( .A(n6140), .B(n35), .C(n2347), .Y(n34) );
  INVX1 U918 ( .A(n34), .Y(n8517) );
  INVX1 U919 ( .A(oprA[11]), .Y(n36) );
  INVX8 U920 ( .A(n36), .Y(n37) );
  INVX8 U921 ( .A(n26), .Y(n44) );
  INVX2 U922 ( .A(n6300), .Y(n5976) );
  OR2X1 U923 ( .A(n4453), .B(n4454), .Y(n4451) );
  INVX1 U924 ( .A(n10465), .Y(n38) );
  AND2X1 U925 ( .A(n1957), .B(n4577), .Y(n10465) );
  INVX1 U926 ( .A(oprB[62]), .Y(n6159) );
  AND2X2 U927 ( .A(n6187), .B(n6186), .Y(n5767) );
  INVX2 U928 ( .A(n6320), .Y(n6000) );
  INVX1 U929 ( .A(n9411), .Y(n39) );
  AND2X1 U930 ( .A(n99), .B(n4516), .Y(n9411) );
  INVX2 U931 ( .A(n6306), .Y(n5982) );
  INVX1 U932 ( .A(n6273), .Y(n5917) );
  INVX4 U933 ( .A(n6307), .Y(n5984) );
  INVX1 U934 ( .A(n6320), .Y(n5999) );
  INVX8 U935 ( .A(n6027), .Y(n6028) );
  INVX2 U936 ( .A(oprA[13]), .Y(n6027) );
  INVX8 U937 ( .A(n5936), .Y(n5938) );
  INVX8 U938 ( .A(n5936), .Y(n5937) );
  INVX8 U939 ( .A(n6312), .Y(n5990) );
  INVX4 U940 ( .A(n6276), .Y(n6275) );
  NOR3X1 U941 ( .A(n41), .B(n10452), .C(n42), .Y(n40) );
  INVX2 U942 ( .A(n40), .Y(n10458) );
  INVX1 U943 ( .A(n10451), .Y(n42) );
  OR2X2 U944 ( .A(n104), .B(n2146), .Y(n8401) );
  INVX1 U945 ( .A(n26), .Y(n43) );
  INVX8 U946 ( .A(n6311), .Y(n5989) );
  AND2X2 U947 ( .A(n6042), .B(n6080), .Y(n10303) );
  INVX1 U948 ( .A(n6295), .Y(n45) );
  INVX4 U949 ( .A(n5917), .Y(n5918) );
  INVX4 U950 ( .A(n25), .Y(n46) );
  OAI21X1 U951 ( .A(n48), .B(n6132), .C(n49), .Y(n47) );
  INVX1 U952 ( .A(n10602), .Y(n49) );
  INVX8 U953 ( .A(n5909), .Y(n5912) );
  INVX2 U954 ( .A(n6166), .Y(n6165) );
  INVX1 U955 ( .A(n6316), .Y(n6315) );
  INVX2 U956 ( .A(oprA[29]), .Y(n6316) );
  INVX1 U957 ( .A(n6019), .Y(n6336) );
  INVX1 U958 ( .A(n46), .Y(n50) );
  BUFX2 U959 ( .A(n6262), .Y(n51) );
  INVX2 U960 ( .A(oprB[5]), .Y(n6262) );
  INVX4 U961 ( .A(n6348), .Y(n6347) );
  OR2X2 U962 ( .A(n6061), .B(n6260), .Y(n10153) );
  AND2X2 U963 ( .A(n6258), .B(n6260), .Y(n10355) );
  INVX8 U964 ( .A(n6341), .Y(n6025) );
  INVX4 U965 ( .A(n6302), .Y(n5978) );
  BUFX2 U966 ( .A(n6037), .Y(n5277) );
  INVX2 U967 ( .A(oprB[6]), .Y(n6260) );
  INVX4 U968 ( .A(n6312), .Y(n5991) );
  INVX8 U969 ( .A(n6236), .Y(n5280) );
  INVX8 U970 ( .A(n5943), .Y(n5944) );
  INVX8 U971 ( .A(n6192), .Y(n6191) );
  INVX1 U972 ( .A(n6323), .Y(n52) );
  INVX1 U973 ( .A(n57), .Y(n58) );
  OAI21X1 U974 ( .A(n54), .B(n6146), .C(n55), .Y(n53) );
  INVX1 U975 ( .A(n53), .Y(n10552) );
  INVX1 U976 ( .A(n10551), .Y(n55) );
  BUFX2 U977 ( .A(n6226), .Y(n56) );
  INVX1 U978 ( .A(n840), .Y(n61) );
  INVX1 U979 ( .A(oprA[17]), .Y(n6338) );
  INVX1 U980 ( .A(n6221), .Y(n6220) );
  AND2X1 U981 ( .A(n98), .B(n1944), .Y(n3901) );
  AND2X2 U982 ( .A(n5915), .B(n9969), .Y(n7106) );
  INVX2 U983 ( .A(oprA[26]), .Y(n6320) );
  INVX8 U984 ( .A(n6161), .Y(n5902) );
  INVX8 U985 ( .A(n5979), .Y(n5980) );
  INVX4 U986 ( .A(oprA[63]), .Y(n5909) );
  INVX2 U987 ( .A(n6293), .Y(n5953) );
  INVX8 U988 ( .A(n6298), .Y(n5970) );
  INVX1 U989 ( .A(n6321), .Y(n57) );
  INVX1 U990 ( .A(n57), .Y(n6001) );
  BUFX4 U991 ( .A(oprA[24]), .Y(n5274) );
  INVX4 U992 ( .A(n6161), .Y(n5903) );
  AND2X2 U993 ( .A(n6076), .B(n6314), .Y(n6435) );
  INVX8 U994 ( .A(n6310), .Y(n5986) );
  INVX4 U995 ( .A(n6359), .Y(n6060) );
  INVX4 U996 ( .A(oprA[59]), .Y(n65) );
  INVX2 U997 ( .A(n6223), .Y(n6222) );
  INVX2 U998 ( .A(n6293), .Y(n5954) );
  OAI21X1 U999 ( .A(n61), .B(n6146), .C(n10608), .Y(n60) );
  INVX1 U1000 ( .A(n60), .Y(n10610) );
  INVX8 U1001 ( .A(n6242), .Y(n6241) );
  INVX1 U1002 ( .A(oprA[58]), .Y(n6278) );
  INVX8 U1003 ( .A(n6219), .Y(n5908) );
  INVX8 U1004 ( .A(n6002), .Y(n6003) );
  INVX2 U1005 ( .A(n6285), .Y(n5933) );
  INVX8 U1006 ( .A(n6200), .Y(n6199) );
  OAI21X1 U1007 ( .A(n63), .B(op[0]), .C(n64), .Y(n62) );
  INVX1 U1008 ( .A(n62), .Y(n8469) );
  INVX1 U1009 ( .A(n8466), .Y(n64) );
  OAI21X1 U1010 ( .A(n69), .B(n6124), .C(n2362), .Y(n68) );
  INVX1 U1011 ( .A(n68), .Y(n10601) );
  INVX8 U1012 ( .A(n6033), .Y(n6034) );
  INVX2 U1013 ( .A(n6198), .Y(n6197) );
  BUFX2 U1014 ( .A(n23), .Y(n70) );
  INVX8 U1015 ( .A(n6292), .Y(n5949) );
  INVX2 U1016 ( .A(n5909), .Y(n5911) );
  INVX2 U1017 ( .A(oprA[30]), .Y(n6313) );
  INVX2 U1018 ( .A(oprB[27]), .Y(n6223) );
  INVX2 U1019 ( .A(n6294), .Y(n5957) );
  BUFX2 U1020 ( .A(n6227), .Y(n71) );
  INVX1 U1021 ( .A(oprA[6]), .Y(n6348) );
  INVX8 U1022 ( .A(n6030), .Y(n6031) );
  INVX4 U1023 ( .A(n6353), .Y(n6054) );
  AND2X2 U1024 ( .A(n5819), .B(n6233), .Y(n9309) );
  INVX8 U1025 ( .A(n6210), .Y(n6209) );
  INVX8 U1026 ( .A(n6355), .Y(n6057) );
  INVX1 U1027 ( .A(oprA[1]), .Y(n6358) );
  INVX8 U1028 ( .A(n6309), .Y(n5987) );
  INVX8 U1029 ( .A(n6295), .Y(n5966) );
  INVX8 U1030 ( .A(n6014), .Y(n6016) );
  INVX4 U1031 ( .A(n6294), .Y(n5956) );
  INVX2 U1032 ( .A(n6044), .Y(n5734) );
  INVX2 U1033 ( .A(n5971), .Y(n5973) );
  INVX8 U1034 ( .A(n6178), .Y(n6177) );
  INVX2 U1035 ( .A(n6), .Y(n6049) );
  BUFX4 U1036 ( .A(n6012), .Y(n5269) );
  INVX4 U1037 ( .A(oprA[23]), .Y(n6329) );
  INVX8 U1038 ( .A(n6214), .Y(n6213) );
  INVX8 U1039 ( .A(n6170), .Y(n6169) );
  INVX8 U1040 ( .A(n6235), .Y(n6234) );
  INVX4 U1041 ( .A(n6355), .Y(n6056) );
  INVX8 U1042 ( .A(n6212), .Y(n6211) );
  BUFX4 U1043 ( .A(n6013), .Y(n5285) );
  INVX1 U1044 ( .A(oprA[25]), .Y(n6323) );
  INVX2 U1045 ( .A(oprA[31]), .Y(n6312) );
  INVX8 U1046 ( .A(n5967), .Y(n5968) );
  INVX8 U1047 ( .A(n5967), .Y(n5969) );
  INVX2 U1048 ( .A(oprA[13]), .Y(n6343) );
  INVX4 U1049 ( .A(n6343), .Y(n6342) );
  INVX2 U1050 ( .A(n6050), .Y(n6052) );
  INVX8 U1051 ( .A(n6182), .Y(n6181) );
  INVX2 U1052 ( .A(oprB[38]), .Y(n6204) );
  INVX8 U1053 ( .A(n6204), .Y(n6203) );
  INVX2 U1054 ( .A(oprB[17]), .Y(n6240) );
  INVX8 U1055 ( .A(n6240), .Y(n6239) );
  INVX1 U1056 ( .A(n5268), .Y(n72) );
  BUFX4 U1057 ( .A(n5999), .Y(n5268) );
  INVX8 U1058 ( .A(n5962), .Y(n5963) );
  INVX8 U1059 ( .A(n6206), .Y(n6205) );
  INVX8 U1060 ( .A(n6352), .Y(n6351) );
  INVX2 U1061 ( .A(n6044), .Y(n6045) );
  INVX2 U1062 ( .A(oprB[36]), .Y(n6208) );
  INVX8 U1063 ( .A(n6252), .Y(n6251) );
  INVX8 U1064 ( .A(n6256), .Y(n6255) );
  INVX4 U1065 ( .A(oprA[62]), .Y(n5913) );
  INVX8 U1066 ( .A(n5913), .Y(n5914) );
  AND2X2 U1067 ( .A(n24), .B(n6244), .Y(n9577) );
  AND2X2 U1068 ( .A(n6319), .B(n9632), .Y(n8936) );
  INVX8 U1069 ( .A(n6292), .Y(n5948) );
  INVX8 U1070 ( .A(n6202), .Y(n6201) );
  INVX2 U1071 ( .A(oprB[24]), .Y(n6229) );
  INVX8 U1072 ( .A(n6229), .Y(n6228) );
  INVX8 U1073 ( .A(n5950), .Y(n5951) );
  INVX8 U1074 ( .A(n6036), .Y(n6037) );
  INVX8 U1075 ( .A(n5943), .Y(n5945) );
  INVX2 U1076 ( .A(oprB[4]), .Y(n6264) );
  INVX4 U1077 ( .A(n6281), .Y(n5926) );
  INVX2 U1078 ( .A(n5913), .Y(n5915) );
  INVX8 U1079 ( .A(n6274), .Y(n5919) );
  INVX4 U1080 ( .A(n5950), .Y(n5952) );
  INVX4 U1081 ( .A(n6285), .Y(n5935) );
  INVX8 U1082 ( .A(n6289), .Y(n5942) );
  INVX4 U1083 ( .A(oprA[7]), .Y(n6040) );
  INVX8 U1084 ( .A(n6357), .Y(n6059) );
  INVX8 U1085 ( .A(n6341), .Y(n6026) );
  INVX4 U1086 ( .A(n6050), .Y(n6051) );
  INVX8 U1087 ( .A(n6254), .Y(n6253) );
  INVX4 U1088 ( .A(oprA[22]), .Y(n6005) );
  INVX8 U1089 ( .A(n6216), .Y(n6215) );
  INVX8 U1090 ( .A(n5939), .Y(n5940) );
  INVX4 U1091 ( .A(n5962), .Y(n5965) );
  INVX8 U1092 ( .A(n1), .Y(n6004) );
  INVX8 U1093 ( .A(n5939), .Y(n5941) );
  INVX8 U1094 ( .A(n6272), .Y(n6271) );
  INVX8 U1095 ( .A(n5959), .Y(n5960) );
  INVX8 U1096 ( .A(n5923), .Y(n5924) );
  INVX8 U1097 ( .A(n6316), .Y(n6314) );
  INVX8 U1098 ( .A(n6268), .Y(n6267) );
  INVX8 U1099 ( .A(n6017), .Y(n6018) );
  INVX4 U1100 ( .A(oprA[21]), .Y(n6333) );
  INVX8 U1101 ( .A(n6250), .Y(n6249) );
  INVX8 U1102 ( .A(n6260), .Y(n6259) );
  AND2X2 U1103 ( .A(n6259), .B(n6258), .Y(n5793) );
  INVX8 U1104 ( .A(n6262), .Y(n6261) );
  INVX8 U1105 ( .A(n6333), .Y(n6009) );
  INVX4 U1106 ( .A(oprB[14]), .Y(n6244) );
  INVX8 U1107 ( .A(n6244), .Y(n6243) );
  BUFX4 U1108 ( .A(n5284), .Y(n5267) );
  INVX8 U1109 ( .A(n6233), .Y(n6232) );
  INVX2 U1110 ( .A(n6294), .Y(n5958) );
  INVX2 U1111 ( .A(n6291), .Y(n6290) );
  INVX1 U1112 ( .A(n7503), .Y(n73) );
  INVX1 U1113 ( .A(n9435), .Y(n74) );
  INVX1 U1114 ( .A(n10329), .Y(n75) );
  BUFX2 U1115 ( .A(n6384), .Y(n76) );
  BUFX2 U1116 ( .A(n6386), .Y(n77) );
  BUFX2 U1117 ( .A(n6400), .Y(n78) );
  BUFX2 U1118 ( .A(n6402), .Y(n79) );
  BUFX2 U1119 ( .A(n6416), .Y(n80) );
  BUFX2 U1120 ( .A(n6422), .Y(n81) );
  BUFX2 U1121 ( .A(n7556), .Y(n82) );
  BUFX2 U1122 ( .A(n9469), .Y(n83) );
  BUFX2 U1123 ( .A(n10607), .Y(n84) );
  BUFX2 U1124 ( .A(n10615), .Y(result[33]) );
  BUFX2 U1125 ( .A(n10614), .Y(result[32]) );
  BUFX2 U1126 ( .A(n9486), .Y(n87) );
  AND2X2 U1127 ( .A(n10552), .B(n100), .Y(n10613) );
  INVX1 U1128 ( .A(n10613), .Y(result[1]) );
  AND2X2 U1129 ( .A(n10610), .B(n97), .Y(n10612) );
  INVX1 U1130 ( .A(n10612), .Y(result[0]) );
  BUFX2 U1131 ( .A(n6393), .Y(n90) );
  BUFX2 U1132 ( .A(n6401), .Y(n91) );
  BUFX2 U1133 ( .A(n8265), .Y(n92) );
  BUFX2 U1134 ( .A(n9535), .Y(n93) );
  BUFX2 U1135 ( .A(n10319), .Y(n94) );
  AND2X2 U1136 ( .A(n6142), .B(n148), .Y(n8516) );
  INVX1 U1137 ( .A(n8516), .Y(n95) );
  AND2X1 U1138 ( .A(n519), .B(n5773), .Y(n10606) );
  INVX1 U1139 ( .A(n10606), .Y(n96) );
  BUFX2 U1140 ( .A(n10609), .Y(n97) );
  BUFX2 U1141 ( .A(n7487), .Y(n98) );
  BUFX2 U1142 ( .A(n9408), .Y(n99) );
  BUFX2 U1143 ( .A(n10553), .Y(n100) );
  BUFX2 U1144 ( .A(n8204), .Y(n101) );
  BUFX2 U1145 ( .A(n8311), .Y(n102) );
  BUFX2 U1146 ( .A(n8412), .Y(n103) );
  BUFX2 U1147 ( .A(n8394), .Y(n104) );
  BUFX2 U1148 ( .A(n8460), .Y(n105) );
  BUFX2 U1149 ( .A(n10478), .Y(n106) );
  BUFX2 U1150 ( .A(n7397), .Y(n107) );
  BUFX2 U1151 ( .A(n7463), .Y(n108) );
  BUFX2 U1152 ( .A(n7515), .Y(n109) );
  BUFX2 U1153 ( .A(n8015), .Y(n110) );
  BUFX2 U1154 ( .A(n8285), .Y(n111) );
  BUFX2 U1155 ( .A(n8411), .Y(n112) );
  BUFX2 U1156 ( .A(n9307), .Y(n113) );
  BUFX2 U1157 ( .A(n9320), .Y(n114) );
  BUFX2 U1158 ( .A(n9422), .Y(n115) );
  BUFX2 U1159 ( .A(n9542), .Y(n116) );
  BUFX2 U1160 ( .A(n10061), .Y(n117) );
  BUFX2 U1161 ( .A(n10410), .Y(n118) );
  BUFX2 U1162 ( .A(n10477), .Y(n119) );
  BUFX2 U1163 ( .A(n7453), .Y(n120) );
  BUFX2 U1164 ( .A(n8511), .Y(n121) );
  BUFX2 U1165 ( .A(n9533), .Y(n122) );
  BUFX2 U1166 ( .A(n10539), .Y(n123) );
  AND2X2 U1167 ( .A(n96), .B(n84), .Y(n10608) );
  BUFX2 U1168 ( .A(n7514), .Y(n124) );
  BUFX2 U1169 ( .A(n8014), .Y(n125) );
  BUFX2 U1170 ( .A(n8410), .Y(n126) );
  BUFX2 U1171 ( .A(n8470), .Y(n127) );
  BUFX2 U1172 ( .A(n8465), .Y(n128) );
  BUFX2 U1173 ( .A(n9421), .Y(n129) );
  BUFX2 U1174 ( .A(n9541), .Y(n130) );
  BUFX2 U1175 ( .A(n10060), .Y(n131) );
  BUFX2 U1176 ( .A(n10409), .Y(n132) );
  BUFX2 U1177 ( .A(n10461), .Y(n133) );
  BUFX2 U1178 ( .A(n10476), .Y(n134) );
  BUFX2 U1179 ( .A(n10542), .Y(n135) );
  INVX1 U1180 ( .A(n10549), .Y(n136) );
  BUFX2 U1181 ( .A(n8405), .Y(n137) );
  BUFX2 U1182 ( .A(n9416), .Y(n138) );
  BUFX2 U1183 ( .A(n10471), .Y(n139) );
  AND2X2 U1184 ( .A(n5411), .B(n93), .Y(n9536) );
  INVX1 U1185 ( .A(n9536), .Y(n140) );
  AND2X1 U1186 ( .A(n1274), .B(n5785), .Y(n10600) );
  INVX1 U1187 ( .A(n10600), .Y(n141) );
  BUFX2 U1188 ( .A(n8468), .Y(n142) );
  BUFX2 U1189 ( .A(n8518), .Y(n143) );
  BUFX2 U1190 ( .A(n10599), .Y(n144) );
  BUFX2 U1191 ( .A(n9481), .Y(n145) );
  BUFX2 U1192 ( .A(n10466), .Y(n146) );
  INVX8 U1193 ( .A(n5994), .Y(n5995) );
  AND2X2 U1194 ( .A(n6232), .B(n5272), .Y(n5762) );
  INVX8 U1195 ( .A(n6264), .Y(n6263) );
  AND2X1 U1196 ( .A(n9626), .B(n5885), .Y(n9987) );
  AND2X1 U1197 ( .A(n5800), .B(n5885), .Y(n10025) );
  INVX1 U1198 ( .A(n8515), .Y(n147) );
  INVX1 U1199 ( .A(n147), .Y(n148) );
  INVX1 U1200 ( .A(n10547), .Y(n149) );
  INVX1 U1201 ( .A(n149), .Y(n150) );
  AND2X2 U1202 ( .A(n6151), .B(n6218), .Y(n8554) );
  INVX1 U1203 ( .A(n8554), .Y(n151) );
  OR2X1 U1204 ( .A(n3692), .B(n3693), .Y(n3689) );
  OR2X1 U1205 ( .A(n3690), .B(n3691), .Y(n3693) );
  OR2X1 U1206 ( .A(n3697), .B(n3698), .Y(n3694) );
  OR2X1 U1207 ( .A(n3695), .B(n3696), .Y(n3698) );
  OR2X1 U1208 ( .A(n3701), .B(n3702), .Y(n3699) );
  OR2X1 U1209 ( .A(n6714), .B(n3700), .Y(n3702) );
  OR2X1 U1210 ( .A(n3706), .B(n3707), .Y(n3703) );
  OR2X1 U1211 ( .A(n3704), .B(n3705), .Y(n3707) );
  OR2X1 U1212 ( .A(n3711), .B(n3712), .Y(n3708) );
  OR2X1 U1213 ( .A(n3709), .B(n3710), .Y(n3712) );
  OR2X1 U1214 ( .A(n3717), .B(n3718), .Y(n3714) );
  OR2X1 U1215 ( .A(n3715), .B(n3716), .Y(n3718) );
  OR2X1 U1216 ( .A(n3721), .B(n3722), .Y(n3719) );
  OR2X1 U1217 ( .A(n3720), .B(n6887), .Y(n3722) );
  OR2X1 U1218 ( .A(n3727), .B(n3728), .Y(n3724) );
  OR2X1 U1219 ( .A(n3725), .B(n3726), .Y(n3728) );
  OR2X1 U1220 ( .A(n3732), .B(n3733), .Y(n3729) );
  OR2X1 U1221 ( .A(n3730), .B(n3731), .Y(n3733) );
  OR2X1 U1222 ( .A(n3737), .B(n3738), .Y(n3734) );
  OR2X1 U1223 ( .A(n3735), .B(n3736), .Y(n3738) );
  OR2X1 U1224 ( .A(n3742), .B(n3743), .Y(n3739) );
  OR2X1 U1225 ( .A(n3740), .B(n3741), .Y(n3743) );
  OR2X1 U1226 ( .A(n3746), .B(n3747), .Y(n3744) );
  OR2X1 U1227 ( .A(n3745), .B(n7078), .Y(n3747) );
  OR2X1 U1228 ( .A(n3750), .B(n3751), .Y(n3748) );
  OR2X1 U1229 ( .A(n3749), .B(n7144), .Y(n3751) );
  OR2X1 U1230 ( .A(n3755), .B(n3756), .Y(n3752) );
  OR2X1 U1231 ( .A(n3753), .B(n3754), .Y(n3756) );
  OR2X1 U1232 ( .A(n3761), .B(n3762), .Y(n3758) );
  OR2X1 U1233 ( .A(n3759), .B(n3760), .Y(n3762) );
  OR2X1 U1234 ( .A(n3766), .B(n3767), .Y(n3763) );
  OR2X1 U1235 ( .A(n3764), .B(n3765), .Y(n3767) );
  OR2X1 U1236 ( .A(n3899), .B(n3900), .Y(n3768) );
  OR2X1 U1237 ( .A(n3769), .B(n3770), .Y(n3900) );
  OR2X1 U1238 ( .A(n3905), .B(n3906), .Y(n3902) );
  OR2X1 U1239 ( .A(n3903), .B(n3904), .Y(n3906) );
  OR2X1 U1240 ( .A(n3908), .B(n3909), .Y(n3911) );
  OR2X1 U1241 ( .A(n3914), .B(n3915), .Y(n3912) );
  OR2X1 U1242 ( .A(n7741), .B(n3913), .Y(n3915) );
  OR2X1 U1243 ( .A(n3920), .B(n3921), .Y(n3917) );
  OR2X1 U1244 ( .A(n3918), .B(n3919), .Y(n3921) );
  OR2X1 U1245 ( .A(n3925), .B(n3926), .Y(n3922) );
  OR2X1 U1246 ( .A(n3923), .B(n3924), .Y(n3926) );
  OR2X1 U1247 ( .A(n3930), .B(n3931), .Y(n3927) );
  OR2X1 U1248 ( .A(n3928), .B(n3929), .Y(n3931) );
  OR2X1 U1249 ( .A(n3934), .B(n3935), .Y(n3932) );
  OR2X1 U1250 ( .A(n3933), .B(n7917), .Y(n3935) );
  OR2X1 U1251 ( .A(n3939), .B(n3940), .Y(n3936) );
  OR2X1 U1252 ( .A(n3937), .B(n3938), .Y(n3940) );
  OR2X1 U1253 ( .A(n3944), .B(n3945), .Y(n3941) );
  OR2X1 U1254 ( .A(n3942), .B(n3943), .Y(n3945) );
  OR2X1 U1255 ( .A(n3949), .B(n3950), .Y(n3946) );
  OR2X1 U1256 ( .A(n3947), .B(n3948), .Y(n3950) );
  OR2X1 U1257 ( .A(n3954), .B(n3955), .Y(n3951) );
  OR2X1 U1258 ( .A(n3952), .B(n3953), .Y(n3955) );
  OR2X1 U1259 ( .A(n3959), .B(n3960), .Y(n3957) );
  OR2X1 U1260 ( .A(n3958), .B(n8169), .Y(n3960) );
  OR2X1 U1261 ( .A(n3964), .B(n3965), .Y(n3961) );
  OR2X1 U1262 ( .A(n3962), .B(n3963), .Y(n3965) );
  OR2X1 U1263 ( .A(n3970), .B(n3971), .Y(n3967) );
  OR2X1 U1264 ( .A(n3968), .B(n3969), .Y(n3971) );
  OR2X1 U1265 ( .A(n3975), .B(n3976), .Y(n3972) );
  OR2X1 U1266 ( .A(n3973), .B(n3974), .Y(n3976) );
  OR2X1 U1267 ( .A(n3980), .B(n3981), .Y(n3977) );
  OR2X1 U1268 ( .A(n3978), .B(n3979), .Y(n3981) );
  OR2X1 U1269 ( .A(n3985), .B(n3986), .Y(n3982) );
  OR2X1 U1270 ( .A(n3983), .B(n3984), .Y(n3986) );
  OR2X1 U1271 ( .A(n3990), .B(n3991), .Y(n3987) );
  OR2X1 U1272 ( .A(n3988), .B(n3989), .Y(n3991) );
  OR2X1 U1273 ( .A(n3994), .B(n3995), .Y(n3992) );
  OR2X1 U1274 ( .A(n3993), .B(n8655), .Y(n3995) );
  OR2X1 U1275 ( .A(n3999), .B(n4000), .Y(n3997) );
  OR2X1 U1276 ( .A(n8748), .B(n3998), .Y(n4000) );
  OR2X1 U1277 ( .A(n4005), .B(n4006), .Y(n4002) );
  OR2X1 U1278 ( .A(n4003), .B(n4004), .Y(n4006) );
  OR2X1 U1279 ( .A(n4011), .B(n4012), .Y(n4008) );
  OR2X1 U1280 ( .A(n4009), .B(n4010), .Y(n4012) );
  OR2X1 U1281 ( .A(n4015), .B(n4016), .Y(n4013) );
  OR2X1 U1282 ( .A(n4014), .B(n8913), .Y(n4016) );
  OR2X1 U1283 ( .A(n4021), .B(n4022), .Y(n4018) );
  OR2X1 U1284 ( .A(n4019), .B(n4020), .Y(n4022) );
  OR2X1 U1285 ( .A(n4026), .B(n4027), .Y(n4023) );
  OR2X1 U1286 ( .A(n4024), .B(n4025), .Y(n4027) );
  OR2X1 U1287 ( .A(n4031), .B(n4032), .Y(n4028) );
  OR2X1 U1288 ( .A(n4029), .B(n4030), .Y(n4032) );
  OR2X1 U1289 ( .A(n4037), .B(n4038), .Y(n4035) );
  OR2X1 U1290 ( .A(n4036), .B(n9181), .Y(n4038) );
  OR2X1 U1291 ( .A(n4042), .B(n4043), .Y(n4039) );
  OR2X1 U1292 ( .A(n4040), .B(n4041), .Y(n4043) );
  OR2X1 U1293 ( .A(n4045), .B(n4046), .Y(n4048) );
  OR2X1 U1294 ( .A(n4052), .B(n4053), .Y(n4049) );
  OR2X1 U1295 ( .A(n4050), .B(n4051), .Y(n4053) );
  OR2X1 U1296 ( .A(n4057), .B(n4058), .Y(n4055) );
  OR2X1 U1297 ( .A(n4056), .B(n9439), .Y(n4058) );
  OR2X1 U1298 ( .A(n4061), .B(n4062), .Y(n4059) );
  OR2X1 U1299 ( .A(n4060), .B(n9494), .Y(n4062) );
  OR2X1 U1300 ( .A(n4066), .B(n4067), .Y(n4063) );
  OR2X1 U1301 ( .A(n4064), .B(n4065), .Y(n4067) );
  OR2X1 U1302 ( .A(n4071), .B(n4072), .Y(n4069) );
  OR2X1 U1303 ( .A(n9777), .B(n4070), .Y(n4072) );
  OR2X1 U1304 ( .A(n4077), .B(n4078), .Y(n4074) );
  OR2X1 U1305 ( .A(n4075), .B(n4076), .Y(n4078) );
  OR2X1 U1306 ( .A(n4083), .B(n4084), .Y(n4080) );
  OR2X1 U1307 ( .A(n4081), .B(n4082), .Y(n4084) );
  OR2X1 U1308 ( .A(n4087), .B(n4088), .Y(n4085) );
  OR2X1 U1309 ( .A(n4086), .B(n9962), .Y(n4088) );
  OR2X1 U1310 ( .A(n4092), .B(n4093), .Y(n4089) );
  OR2X1 U1311 ( .A(n4090), .B(n4091), .Y(n4093) );
  OR2X1 U1312 ( .A(n4097), .B(n4098), .Y(n4094) );
  OR2X1 U1313 ( .A(n4095), .B(n4096), .Y(n4098) );
  OR2X1 U1314 ( .A(n4102), .B(n4103), .Y(n4099) );
  OR2X1 U1315 ( .A(n4100), .B(n4101), .Y(n4103) );
  OR2X1 U1316 ( .A(n4108), .B(n4109), .Y(n4106) );
  OR2X1 U1317 ( .A(n4107), .B(n10220), .Y(n4109) );
  OR2X1 U1318 ( .A(n4113), .B(n4114), .Y(n4110) );
  OR2X1 U1319 ( .A(n4111), .B(n4112), .Y(n4114) );
  OR2X1 U1320 ( .A(n4119), .B(n4120), .Y(n4116) );
  OR2X1 U1321 ( .A(n4117), .B(n4118), .Y(n4120) );
  OR2X1 U1322 ( .A(n4133), .B(n4134), .Y(n4131) );
  OR2X1 U1323 ( .A(n4132), .B(n6989), .Y(n4134) );
  OR2X1 U1324 ( .A(n4137), .B(n4138), .Y(n4135) );
  OR2X1 U1325 ( .A(n4136), .B(n7046), .Y(n4138) );
  OR2X1 U1326 ( .A(n4141), .B(n4142), .Y(n4139) );
  OR2X1 U1327 ( .A(n4140), .B(n7114), .Y(n4142) );
  OR2X1 U1328 ( .A(n4145), .B(n4146), .Y(n4143) );
  OR2X1 U1329 ( .A(n4144), .B(n7189), .Y(n4146) );
  OR2X1 U1330 ( .A(n4149), .B(n4150), .Y(n4147) );
  OR2X1 U1331 ( .A(n4148), .B(n7256), .Y(n4150) );
  OR2X1 U1332 ( .A(n4153), .B(n4154), .Y(n4151) );
  OR2X1 U1333 ( .A(n4152), .B(n7382), .Y(n4154) );
  OR2X1 U1334 ( .A(n4157), .B(n4158), .Y(n4155) );
  OR2X1 U1335 ( .A(n4156), .B(n7708), .Y(n4158) );
  OR2X1 U1336 ( .A(n4165), .B(n4166), .Y(n4163) );
  OR2X1 U1337 ( .A(n4164), .B(n7948), .Y(n4166) );
  OR2X1 U1338 ( .A(n4173), .B(n4174), .Y(n4171) );
  OR2X1 U1339 ( .A(n4172), .B(n8059), .Y(n4174) );
  OR2X1 U1340 ( .A(n4177), .B(n4178), .Y(n4175) );
  OR2X1 U1341 ( .A(n4176), .B(n8396), .Y(n4178) );
  OR2X1 U1342 ( .A(n4181), .B(n4182), .Y(n4179) );
  OR2X1 U1343 ( .A(n4180), .B(n8713), .Y(n4182) );
  OR2X1 U1344 ( .A(n4185), .B(n4186), .Y(n4183) );
  OR2X1 U1345 ( .A(n4184), .B(n8830), .Y(n4186) );
  OR2X1 U1346 ( .A(n4190), .B(n4191), .Y(n4188) );
  OR2X1 U1347 ( .A(n4189), .B(n9013), .Y(n4191) );
  OR2X1 U1348 ( .A(n4194), .B(n4195), .Y(n4192) );
  OR2X1 U1349 ( .A(n4193), .B(n9070), .Y(n4195) );
  OR2X1 U1350 ( .A(n4198), .B(n4199), .Y(n4196) );
  OR2X1 U1351 ( .A(n4197), .B(n9406), .Y(n4199) );
  OR2X1 U1352 ( .A(n4202), .B(n4203), .Y(n4200) );
  OR2X1 U1353 ( .A(n4201), .B(n9446), .Y(n4203) );
  OR2X1 U1354 ( .A(n4206), .B(n4207), .Y(n4204) );
  OR2X1 U1355 ( .A(n4205), .B(n9743), .Y(n4207) );
  OR2X1 U1356 ( .A(n4209), .B(n9866), .Y(n4211) );
  OR2X1 U1357 ( .A(n4214), .B(n4215), .Y(n4212) );
  OR2X1 U1358 ( .A(n4213), .B(n9994), .Y(n4215) );
  OR2X1 U1359 ( .A(n4222), .B(n4223), .Y(n4220) );
  OR2X1 U1360 ( .A(n4221), .B(n10110), .Y(n4223) );
  OR2X1 U1361 ( .A(n4297), .B(n4298), .Y(n4295) );
  OR2X1 U1362 ( .A(n4296), .B(n6604), .Y(n4298) );
  OR2X1 U1363 ( .A(n4304), .B(n4305), .Y(n4299) );
  OR2X1 U1364 ( .A(n4300), .B(n6682), .Y(n4305) );
  OR2X1 U1365 ( .A(n4308), .B(n4309), .Y(n4306) );
  OR2X1 U1366 ( .A(n4307), .B(n6737), .Y(n4309) );
  OR2X1 U1367 ( .A(n5036), .B(n4313), .Y(n4311) );
  OR2X1 U1368 ( .A(n4312), .B(n6794), .Y(n4313) );
  OR2X1 U1369 ( .A(n4319), .B(n4320), .Y(n4314) );
  OR2X1 U1370 ( .A(n4315), .B(n6870), .Y(n4320) );
  OR2X1 U1371 ( .A(n4324), .B(n4325), .Y(n4321) );
  OR2X1 U1372 ( .A(n4322), .B(n4323), .Y(n4325) );
  OR2X1 U1373 ( .A(n6978), .B(n4328), .Y(n4326) );
  OR2X1 U1374 ( .A(n4327), .B(n7233), .Y(n4328) );
  OR2X1 U1375 ( .A(n4334), .B(n4335), .Y(n4329) );
  OR2X1 U1376 ( .A(n4330), .B(n7033), .Y(n4335) );
  OR2X1 U1377 ( .A(n4338), .B(n4339), .Y(n4336) );
  OR2X1 U1378 ( .A(n4337), .B(n7117), .Y(n4339) );
  OR2X1 U1379 ( .A(n7151), .B(n4342), .Y(n4340) );
  OR2X1 U1380 ( .A(n7153), .B(n4341), .Y(n4342) );
  OR2X1 U1381 ( .A(n4345), .B(n4376), .Y(n4343) );
  OR2X1 U1382 ( .A(n4344), .B(n7192), .Y(n4376) );
  OR2X1 U1383 ( .A(n4379), .B(n4380), .Y(n4377) );
  OR2X1 U1384 ( .A(n4378), .B(n7245), .Y(n4380) );
  OR2X1 U1385 ( .A(n4383), .B(n4384), .Y(n4381) );
  OR2X1 U1386 ( .A(n4382), .B(n7320), .Y(n4384) );
  OR2X1 U1387 ( .A(n4386), .B(n7385), .Y(n4388) );
  OR2X1 U1388 ( .A(n4392), .B(n4393), .Y(n4389) );
  OR2X1 U1389 ( .A(n4390), .B(n4391), .Y(n4393) );
  OR2X1 U1390 ( .A(n4396), .B(n4397), .Y(n4394) );
  OR2X1 U1391 ( .A(n4395), .B(n7635), .Y(n4397) );
  OR2X1 U1392 ( .A(n4400), .B(n4401), .Y(n4398) );
  OR2X1 U1393 ( .A(n4399), .B(n7711), .Y(n4401) );
  OR2X1 U1394 ( .A(n4404), .B(n4405), .Y(n4402) );
  OR2X1 U1395 ( .A(n4403), .B(n7759), .Y(n4405) );
  OR2X1 U1396 ( .A(n4408), .B(n4409), .Y(n4406) );
  OR2X1 U1397 ( .A(n4407), .B(n7773), .Y(n4409) );
  OR2X1 U1398 ( .A(n4718), .B(n4412), .Y(n4410) );
  OR2X1 U1399 ( .A(n4411), .B(n7813), .Y(n4412) );
  OR2X1 U1400 ( .A(n4415), .B(n4416), .Y(n4413) );
  OR2X1 U1401 ( .A(n4414), .B(n7889), .Y(n4416) );
  OR2X1 U1402 ( .A(n4718), .B(n4420), .Y(n4417) );
  OR2X1 U1403 ( .A(n4418), .B(n4419), .Y(n4420) );
  OR2X1 U1404 ( .A(n7992), .B(n4423), .Y(n4421) );
  OR2X1 U1405 ( .A(n4422), .B(n8247), .Y(n4423) );
  OR2X1 U1406 ( .A(n4426), .B(n4427), .Y(n4424) );
  OR2X1 U1407 ( .A(n4425), .B(n8046), .Y(n4427) );
  OR2X1 U1408 ( .A(n4430), .B(n4431), .Y(n4428) );
  OR2X1 U1409 ( .A(n4429), .B(n8134), .Y(n4431) );
  OR2X1 U1410 ( .A(n8175), .B(n4434), .Y(n4432) );
  OR2X1 U1411 ( .A(n8177), .B(n4433), .Y(n4434) );
  OR2X1 U1412 ( .A(n4437), .B(n4438), .Y(n4435) );
  OR2X1 U1413 ( .A(n4436), .B(n8208), .Y(n4438) );
  OR2X1 U1414 ( .A(n4441), .B(n4442), .Y(n4439) );
  OR2X1 U1415 ( .A(n4440), .B(n8259), .Y(n4442) );
  OR2X1 U1416 ( .A(n4445), .B(n4446), .Y(n4443) );
  OR2X1 U1417 ( .A(n4444), .B(n8273), .Y(n4446) );
  OR2X1 U1418 ( .A(n4449), .B(n4450), .Y(n4447) );
  OR2X1 U1419 ( .A(n4448), .B(n8336), .Y(n4450) );
  OR2X1 U1420 ( .A(n4720), .B(n4458), .Y(n4455) );
  OR2X1 U1421 ( .A(n4456), .B(n4457), .Y(n4458) );
  OR2X1 U1422 ( .A(n4462), .B(n4463), .Y(n4460) );
  OR2X1 U1423 ( .A(n4461), .B(n8637), .Y(n4463) );
  OR2X1 U1424 ( .A(n4467), .B(n4468), .Y(n4464) );
  OR2X1 U1425 ( .A(n4465), .B(n4466), .Y(n4468) );
  OR2X1 U1426 ( .A(n4471), .B(n4472), .Y(n4469) );
  OR2X1 U1427 ( .A(n4470), .B(n8766), .Y(n4472) );
  OR2X1 U1428 ( .A(n4475), .B(n4476), .Y(n4473) );
  OR2X1 U1429 ( .A(n4474), .B(n8780), .Y(n4476) );
  OR2X1 U1430 ( .A(n5039), .B(n4479), .Y(n4477) );
  OR2X1 U1431 ( .A(n4478), .B(n8820), .Y(n4479) );
  OR2X1 U1432 ( .A(n4482), .B(n4483), .Y(n4480) );
  OR2X1 U1433 ( .A(n4481), .B(n8895), .Y(n4483) );
  OR2X1 U1434 ( .A(n4487), .B(n4488), .Y(n4484) );
  OR2X1 U1435 ( .A(n4485), .B(n4486), .Y(n4488) );
  OR2X1 U1436 ( .A(n9003), .B(n4491), .Y(n4489) );
  OR2X1 U1437 ( .A(n4490), .B(n9258), .Y(n4491) );
  OR2X1 U1438 ( .A(n4494), .B(n4495), .Y(n4492) );
  OR2X1 U1439 ( .A(n4493), .B(n9057), .Y(n4495) );
  OR2X1 U1440 ( .A(n4498), .B(n4499), .Y(n4496) );
  OR2X1 U1441 ( .A(n4497), .B(n9146), .Y(n4499) );
  OR2X1 U1442 ( .A(n9186), .B(n4502), .Y(n4500) );
  OR2X1 U1443 ( .A(n9188), .B(n4501), .Y(n4502) );
  OR2X1 U1444 ( .A(n4506), .B(n4507), .Y(n4504) );
  OR2X1 U1445 ( .A(n4505), .B(n9270), .Y(n4507) );
  OR2X1 U1446 ( .A(n4510), .B(n4511), .Y(n4508) );
  OR2X1 U1447 ( .A(n4509), .B(n9284), .Y(n4511) );
  OR2X1 U1448 ( .A(n4514), .B(n4515), .Y(n4512) );
  OR2X1 U1449 ( .A(n4513), .B(n9346), .Y(n4515) );
  AND2X1 U1450 ( .A(n1952), .B(n1945), .Y(n4516) );
  OR2X1 U1451 ( .A(n4520), .B(n4521), .Y(n4517) );
  OR2X1 U1452 ( .A(n4518), .B(n4519), .Y(n4521) );
  OR2X1 U1453 ( .A(n4524), .B(n4525), .Y(n4522) );
  OR2X1 U1454 ( .A(n9504), .B(n4523), .Y(n4525) );
  OR2X1 U1455 ( .A(n4528), .B(n4529), .Y(n4526) );
  OR2X1 U1456 ( .A(n4527), .B(n9667), .Y(n4529) );
  OR2X1 U1457 ( .A(n4532), .B(n4533), .Y(n4530) );
  OR2X1 U1458 ( .A(n4531), .B(n9746), .Y(n4533) );
  OR2X1 U1459 ( .A(n4536), .B(n4537), .Y(n4534) );
  OR2X1 U1460 ( .A(n4535), .B(n9799), .Y(n4537) );
  OR2X1 U1461 ( .A(n4540), .B(n4541), .Y(n4538) );
  OR2X1 U1462 ( .A(n4539), .B(n9814), .Y(n4541) );
  OR2X1 U1463 ( .A(n4721), .B(n4544), .Y(n4542) );
  OR2X1 U1464 ( .A(n4543), .B(n9856), .Y(n4544) );
  OR2X1 U1465 ( .A(n4547), .B(n4548), .Y(n4545) );
  OR2X1 U1466 ( .A(n4546), .B(n9934), .Y(n4548) );
  OR2X1 U1467 ( .A(n4721), .B(n4552), .Y(n4549) );
  OR2X1 U1468 ( .A(n4550), .B(n4551), .Y(n4552) );
  OR2X1 U1469 ( .A(n10038), .B(n4555), .Y(n4553) );
  OR2X1 U1470 ( .A(n4554), .B(n10300), .Y(n4555) );
  OR2X1 U1471 ( .A(n4558), .B(n4559), .Y(n4556) );
  OR2X1 U1472 ( .A(n4557), .B(n10096), .Y(n4559) );
  OR2X1 U1473 ( .A(n4562), .B(n4563), .Y(n4560) );
  OR2X1 U1474 ( .A(n4561), .B(n10186), .Y(n4563) );
  OR2X1 U1475 ( .A(n10225), .B(n4566), .Y(n4564) );
  OR2X1 U1476 ( .A(n10227), .B(n4565), .Y(n4566) );
  OR2X1 U1477 ( .A(n4570), .B(n4571), .Y(n4568) );
  OR2X1 U1478 ( .A(n4569), .B(n10312), .Y(n4571) );
  AND2X1 U1479 ( .A(n1953), .B(n1947), .Y(n4572) );
  OR2X1 U1480 ( .A(n4575), .B(n4576), .Y(n4573) );
  OR2X1 U1481 ( .A(n4574), .B(n10398), .Y(n4576) );
  OR2X1 U1482 ( .A(n4580), .B(n4581), .Y(n4578) );
  OR2X1 U1483 ( .A(n4579), .B(n10509), .Y(n4581) );
  OR2X1 U1484 ( .A(n4584), .B(n4585), .Y(n4582) );
  OR2X1 U1485 ( .A(n4583), .B(n10577), .Y(n4585) );
  OR2X1 U1486 ( .A(n7157), .B(n4652), .Y(n4650) );
  OR2X1 U1487 ( .A(n4651), .B(n6079), .Y(n4652) );
  OR2X1 U1488 ( .A(n8188), .B(n4655), .Y(n4653) );
  OR2X1 U1489 ( .A(n4654), .B(n6079), .Y(n4655) );
  OR2X1 U1490 ( .A(n9199), .B(n4658), .Y(n4656) );
  INVX1 U1491 ( .A(n4656), .Y(n152) );
  OR2X1 U1492 ( .A(n4657), .B(n6079), .Y(n4658) );
  OR2X1 U1493 ( .A(n10238), .B(n4662), .Y(n4660) );
  INVX1 U1494 ( .A(n4660), .Y(n153) );
  OR2X1 U1495 ( .A(n4661), .B(n6079), .Y(n4662) );
  OR2X1 U1496 ( .A(n10217), .B(n4794), .Y(n4792) );
  INVX1 U1497 ( .A(n4792), .Y(n154) );
  OR2X1 U1498 ( .A(n4793), .B(n10216), .Y(n4794) );
  OR2X1 U1499 ( .A(n7213), .B(n4810), .Y(n4808) );
  OR2X1 U1500 ( .A(n4809), .B(n6708), .Y(n4810) );
  OR2X1 U1501 ( .A(n8230), .B(n4814), .Y(n4812) );
  INVX1 U1502 ( .A(n4812), .Y(n155) );
  OR2X1 U1503 ( .A(n4813), .B(n7735), .Y(n4814) );
  OR2X1 U1504 ( .A(n9242), .B(n4817), .Y(n4815) );
  OR2X1 U1505 ( .A(n4816), .B(n8742), .Y(n4817) );
  OR2X1 U1506 ( .A(n9266), .B(n4821), .Y(n4819) );
  INVX1 U1507 ( .A(n4819), .Y(n156) );
  OR2X1 U1508 ( .A(n4820), .B(n9255), .Y(n4821) );
  OR2X1 U1509 ( .A(n10282), .B(n4825), .Y(n4823) );
  INVX1 U1510 ( .A(n4823), .Y(n157) );
  OR2X1 U1511 ( .A(n4824), .B(n9770), .Y(n4825) );
  OR2X1 U1512 ( .A(n6850), .B(n4851), .Y(n4849) );
  OR2X1 U1513 ( .A(n4850), .B(n6849), .Y(n4851) );
  OR2X1 U1514 ( .A(n9195), .B(n4854), .Y(n4852) );
  OR2X1 U1515 ( .A(n9193), .B(n4853), .Y(n4854) );
  OR2X1 U1516 ( .A(n7163), .B(n4862), .Y(n4860) );
  OR2X1 U1517 ( .A(n7161), .B(n4861), .Y(n4862) );
  OR2X1 U1518 ( .A(n10308), .B(n4865), .Y(n4863) );
  OR2X1 U1519 ( .A(n4864), .B(n10297), .Y(n4865) );
  OR2X1 U1520 ( .A(n8875), .B(n4879), .Y(n4877) );
  OR2X1 U1521 ( .A(n4878), .B(n8874), .Y(n4879) );
  OR2X1 U1522 ( .A(n7087), .B(n4882), .Y(n4880) );
  OR2X1 U1523 ( .A(n4881), .B(n7237), .Y(n4882) );
  OR2X1 U1524 ( .A(n7241), .B(n4885), .Y(n4883) );
  OR2X1 U1525 ( .A(n4884), .B(n7230), .Y(n4885) );
  OR2X1 U1526 ( .A(n8131), .B(n4888), .Y(n4886) );
  OR2X1 U1527 ( .A(n4887), .B(n8251), .Y(n4888) );
  OR2X1 U1528 ( .A(n8232), .B(n4891), .Y(n4889) );
  OR2X1 U1529 ( .A(n8230), .B(n4890), .Y(n4891) );
  OR2X1 U1530 ( .A(n9143), .B(n4894), .Y(n4892) );
  OR2X1 U1531 ( .A(n4893), .B(n9262), .Y(n4894) );
  OR2X1 U1532 ( .A(n10183), .B(n4897), .Y(n4895) );
  OR2X1 U1533 ( .A(n4896), .B(n10304), .Y(n4897) );
  OR2X1 U1534 ( .A(n7868), .B(n4905), .Y(n4903) );
  OR2X1 U1535 ( .A(n4904), .B(n7867), .Y(n4905) );
  OR2X1 U1536 ( .A(n9912), .B(n4908), .Y(n4906) );
  OR2X1 U1537 ( .A(n4907), .B(n9911), .Y(n4908) );
  OR2X1 U1538 ( .A(n7016), .B(n4911), .Y(n4909) );
  OR2X1 U1539 ( .A(n4910), .B(n7015), .Y(n4911) );
  OR2X1 U1540 ( .A(n7093), .B(n4914), .Y(n4912) );
  OR2X1 U1541 ( .A(n4913), .B(n7092), .Y(n4914) );
  OR2X1 U1542 ( .A(n8029), .B(n4917), .Y(n4915) );
  OR2X1 U1543 ( .A(n4916), .B(n8028), .Y(n4917) );
  OR2X1 U1544 ( .A(n8184), .B(n4920), .Y(n4918) );
  OR2X1 U1545 ( .A(n8182), .B(n4919), .Y(n4920) );
  OR2X1 U1546 ( .A(n8255), .B(n4923), .Y(n4921) );
  OR2X1 U1547 ( .A(n4922), .B(n8244), .Y(n4923) );
  OR2X1 U1548 ( .A(n9040), .B(n4926), .Y(n4924) );
  OR2X1 U1549 ( .A(n4925), .B(n9039), .Y(n4926) );
  OR2X1 U1550 ( .A(n9244), .B(n4929), .Y(n4927) );
  OR2X1 U1551 ( .A(n9242), .B(n4928), .Y(n4929) );
  OR2X1 U1552 ( .A(n10076), .B(n4932), .Y(n4930) );
  OR2X1 U1553 ( .A(n4931), .B(n10075), .Y(n4932) );
  OR2X1 U1554 ( .A(n10234), .B(n4935), .Y(n4933) );
  OR2X1 U1555 ( .A(n10232), .B(n4934), .Y(n4935) );
  OR2X1 U1556 ( .A(n10284), .B(n4938), .Y(n4936) );
  OR2X1 U1557 ( .A(n10282), .B(n4937), .Y(n4938) );
  OR2X1 U1558 ( .A(n6910), .B(n4951), .Y(n4949) );
  OR2X1 U1559 ( .A(n7011), .B(n4950), .Y(n4951) );
  OR2X1 U1560 ( .A(n7940), .B(n4954), .Y(n4952) );
  OR2X1 U1561 ( .A(n8024), .B(n4953), .Y(n4954) );
  OR2X1 U1562 ( .A(n8936), .B(n4957), .Y(n4955) );
  OR2X1 U1563 ( .A(n9035), .B(n4956), .Y(n4957) );
  OR2X1 U1564 ( .A(n9986), .B(n4961), .Y(n4959) );
  OR2X1 U1565 ( .A(n10070), .B(n4960), .Y(n4961) );
  OR2X1 U1566 ( .A(n6662), .B(n4975), .Y(n4974) );
  OR2X1 U1567 ( .A(n6661), .B(n7161), .Y(n4975) );
  OR2X1 U1568 ( .A(n7012), .B(n4978), .Y(n4976) );
  OR2X1 U1569 ( .A(n4977), .B(n7011), .Y(n4978) );
  OR2X1 U1570 ( .A(n7215), .B(n4981), .Y(n4979) );
  OR2X1 U1571 ( .A(n7213), .B(n4980), .Y(n4981) );
  OR2X1 U1572 ( .A(n7691), .B(n4983), .Y(n4982) );
  OR2X1 U1573 ( .A(n7690), .B(n8182), .Y(n4983) );
  OR2X1 U1574 ( .A(n8025), .B(n4986), .Y(n4984) );
  OR2X1 U1575 ( .A(n4985), .B(n8024), .Y(n4986) );
  OR2X1 U1576 ( .A(n8126), .B(n4989), .Y(n4987) );
  OR2X1 U1577 ( .A(n4988), .B(n8125), .Y(n4989) );
  OR2X1 U1578 ( .A(n8717), .B(n4991), .Y(n4990) );
  OR2X1 U1579 ( .A(n8716), .B(n9193), .Y(n4991) );
  OR2X1 U1580 ( .A(n9036), .B(n4994), .Y(n4992) );
  OR2X1 U1581 ( .A(n4993), .B(n9035), .Y(n4994) );
  OR2X1 U1582 ( .A(n9138), .B(n4997), .Y(n4995) );
  OR2X1 U1583 ( .A(n4996), .B(n9137), .Y(n4997) );
  OR2X1 U1584 ( .A(n9725), .B(n4999), .Y(n4998) );
  OR2X1 U1585 ( .A(n9724), .B(n10232), .Y(n4999) );
  OR2X1 U1586 ( .A(n10071), .B(n5002), .Y(n5000) );
  OR2X1 U1587 ( .A(n5001), .B(n10070), .Y(n5002) );
  OR2X1 U1588 ( .A(n10178), .B(n5005), .Y(n5003) );
  OR2X1 U1589 ( .A(n5004), .B(n10177), .Y(n5005) );
  OR2X1 U1590 ( .A(n6707), .B(n5015), .Y(n5013) );
  INVX1 U1591 ( .A(n5013), .Y(n158) );
  OR2X1 U1592 ( .A(n5014), .B(n7235), .Y(n5015) );
  OR2X1 U1593 ( .A(n7734), .B(n5018), .Y(n5016) );
  INVX1 U1594 ( .A(n5016), .Y(n159) );
  OR2X1 U1595 ( .A(n5017), .B(n8249), .Y(n5018) );
  OR2X1 U1596 ( .A(n8741), .B(n5021), .Y(n5019) );
  INVX1 U1597 ( .A(n5019), .Y(n160) );
  OR2X1 U1598 ( .A(n5020), .B(n9260), .Y(n5021) );
  OR2X1 U1599 ( .A(n9769), .B(n5024), .Y(n5022) );
  INVX1 U1600 ( .A(n5022), .Y(n161) );
  OR2X1 U1601 ( .A(n5023), .B(n10302), .Y(n5024) );
  OR2X1 U1602 ( .A(n6583), .B(n5027), .Y(n5025) );
  INVX1 U1603 ( .A(n5025), .Y(n162) );
  OR2X1 U1604 ( .A(n5026), .B(n7239), .Y(n5027) );
  OR2X1 U1605 ( .A(n8951), .B(n5035), .Y(n5033) );
  INVX1 U1606 ( .A(n5033), .Y(n163) );
  OR2X1 U1607 ( .A(n5034), .B(n8950), .Y(n5035) );
  OR2X1 U1608 ( .A(n6788), .B(n5038), .Y(n5036) );
  OR2X1 U1609 ( .A(n5037), .B(n6787), .Y(n5038) );
  OR2X1 U1610 ( .A(n8817), .B(n5041), .Y(n5039) );
  OR2X1 U1611 ( .A(n5040), .B(n8816), .Y(n5041) );
  OR2X1 U1612 ( .A(n6911), .B(n5045), .Y(n5043) );
  INVX1 U1613 ( .A(n5043), .Y(n164) );
  OR2X1 U1614 ( .A(n5044), .B(n6910), .Y(n5045) );
  OR2X1 U1615 ( .A(n8937), .B(n5048), .Y(n5046) );
  INVX1 U1616 ( .A(n5046), .Y(n165) );
  OR2X1 U1617 ( .A(n5047), .B(n8936), .Y(n5048) );
  OR2X1 U1618 ( .A(n9991), .B(n5052), .Y(n5050) );
  OR2X1 U1619 ( .A(n5051), .B(n9990), .Y(n5052) );
  OR2X1 U1620 ( .A(n8995), .B(n5055), .Y(n5053) );
  OR2X1 U1621 ( .A(n5054), .B(n8994), .Y(n5055) );
  OR2X1 U1622 ( .A(n7945), .B(n5058), .Y(n5056) );
  OR2X1 U1623 ( .A(n5057), .B(n7944), .Y(n5058) );
  OR2X1 U1624 ( .A(n6925), .B(n5061), .Y(n5059) );
  OR2X1 U1625 ( .A(n5060), .B(n6924), .Y(n5061) );
  OR2X1 U1626 ( .A(n9840), .B(n5064), .Y(n5062) );
  OR2X1 U1627 ( .A(n5063), .B(n9839), .Y(n5064) );
  OR2X1 U1628 ( .A(n7799), .B(n5067), .Y(n5065) );
  OR2X1 U1629 ( .A(n5066), .B(n7798), .Y(n5067) );
  OR2X1 U1630 ( .A(n6963), .B(n5070), .Y(n5068) );
  OR2X1 U1631 ( .A(n5069), .B(n6962), .Y(n5070) );
  OR2X1 U1632 ( .A(n7615), .B(n5073), .Y(n5071) );
  OR2X1 U1633 ( .A(n5072), .B(n8253), .Y(n5073) );
  OR2X1 U1634 ( .A(n8617), .B(n5076), .Y(n5074) );
  OR2X1 U1635 ( .A(n5075), .B(n9264), .Y(n5076) );
  OR2X1 U1636 ( .A(n9646), .B(n5079), .Y(n5077) );
  OR2X1 U1637 ( .A(n5078), .B(n10306), .Y(n5079) );
  OR2X1 U1638 ( .A(n7013), .B(n5082), .Y(n5080) );
  OR2X1 U1639 ( .A(n5081), .B(n7160), .Y(n5082) );
  OR2X1 U1640 ( .A(n7983), .B(n5085), .Y(n5083) );
  OR2X1 U1641 ( .A(n5084), .B(n7982), .Y(n5085) );
  OR2X1 U1642 ( .A(n9037), .B(n5088), .Y(n5086) );
  OR2X1 U1643 ( .A(n5087), .B(n9192), .Y(n5088) );
  OR2X1 U1644 ( .A(n8744), .B(n5091), .Y(n5089) );
  OR2X1 U1645 ( .A(n5090), .B(n9240), .Y(n5091) );
  OR2X1 U1646 ( .A(n10029), .B(n5094), .Y(n5092) );
  OR2X1 U1647 ( .A(n5093), .B(n10028), .Y(n5094) );
  OR2X1 U1648 ( .A(n6777), .B(n5097), .Y(n5095) );
  OR2X1 U1649 ( .A(n5096), .B(n6776), .Y(n5097) );
  OR2X1 U1650 ( .A(n8806), .B(n5100), .Y(n5098) );
  OR2X1 U1651 ( .A(n5099), .B(n8805), .Y(n5100) );
  OR2X1 U1652 ( .A(n7941), .B(n5103), .Y(n5101) );
  OR2X1 U1653 ( .A(n5102), .B(n7940), .Y(n5103) );
  OR2X1 U1654 ( .A(n6710), .B(n5109), .Y(n5107) );
  OR2X1 U1655 ( .A(n5108), .B(n7211), .Y(n5109) );
  OR2X1 U1656 ( .A(n6967), .B(n5112), .Y(n5110) );
  OR2X1 U1657 ( .A(n5111), .B(n6966), .Y(n5112) );
  OR2X1 U1658 ( .A(n8026), .B(n5115), .Y(n5113) );
  OR2X1 U1659 ( .A(n5114), .B(n8181), .Y(n5115) );
  OR2X1 U1660 ( .A(n8125), .B(n5118), .Y(n5116) );
  OR2X1 U1661 ( .A(n5117), .B(n8229), .Y(n5118) );
  OR2X1 U1662 ( .A(n7737), .B(n5121), .Y(n5119) );
  OR2X1 U1663 ( .A(n5120), .B(n8228), .Y(n5121) );
  OR2X1 U1664 ( .A(n7803), .B(n5124), .Y(n5122) );
  OR2X1 U1665 ( .A(n5123), .B(n7802), .Y(n5124) );
  OR2X1 U1666 ( .A(n10073), .B(n5127), .Y(n5125) );
  OR2X1 U1667 ( .A(n5126), .B(n10231), .Y(n5127) );
  OR2X1 U1668 ( .A(n10177), .B(n5130), .Y(n5128) );
  OR2X1 U1669 ( .A(n5129), .B(n10281), .Y(n5130) );
  OR2X1 U1670 ( .A(n9772), .B(n5133), .Y(n5131) );
  OR2X1 U1671 ( .A(n5132), .B(n10280), .Y(n5133) );
  OR2X1 U1672 ( .A(n9844), .B(n5136), .Y(n5134) );
  OR2X1 U1673 ( .A(n5135), .B(n9843), .Y(n5136) );
  OR2X1 U1674 ( .A(n9987), .B(n5139), .Y(n5137) );
  OR2X1 U1675 ( .A(n5138), .B(n9986), .Y(n5139) );
  OR2X1 U1676 ( .A(n6486), .B(n5142), .Y(n5140) );
  OR2X1 U1677 ( .A(n5141), .B(n7009), .Y(n5142) );
  OR2X1 U1678 ( .A(n7530), .B(n5145), .Y(n5143) );
  OR2X1 U1679 ( .A(n5144), .B(n8022), .Y(n5145) );
  OR2X1 U1680 ( .A(n8534), .B(n5148), .Y(n5146) );
  OR2X1 U1681 ( .A(n5147), .B(n9033), .Y(n5148) );
  OR2X1 U1682 ( .A(n9557), .B(n5151), .Y(n5149) );
  OR2X1 U1683 ( .A(n5150), .B(n10068), .Y(n5151) );
  OR2X1 U1684 ( .A(n7979), .B(n5154), .Y(n5152) );
  OR2X1 U1685 ( .A(n5153), .B(n7978), .Y(n5154) );
  OR2X1 U1686 ( .A(n8991), .B(n5157), .Y(n5155) );
  OR2X1 U1687 ( .A(n5156), .B(n8990), .Y(n5157) );
  OR2X1 U1688 ( .A(n7092), .B(n5161), .Y(n5159) );
  OR2X1 U1689 ( .A(n5160), .B(n7212), .Y(n5161) );
  OR2X1 U1690 ( .A(n6781), .B(n5164), .Y(n5162) );
  OR2X1 U1691 ( .A(n5163), .B(n6780), .Y(n5164) );
  OR2X1 U1692 ( .A(n9137), .B(n5167), .Y(n5165) );
  OR2X1 U1693 ( .A(n5166), .B(n9241), .Y(n5167) );
  OR2X1 U1694 ( .A(n8810), .B(n5170), .Y(n5168) );
  OR2X1 U1695 ( .A(n5169), .B(n8809), .Y(n5170) );
  OR2X1 U1696 ( .A(n10025), .B(n5173), .Y(n5171) );
  OR2X1 U1697 ( .A(n5172), .B(n10024), .Y(n5173) );
  OR2X1 U1698 ( .A(n10379), .B(n5177), .Y(n5175) );
  INVX1 U1699 ( .A(n5175), .Y(n166) );
  OR2X1 U1700 ( .A(n5176), .B(n10378), .Y(n5177) );
  OR2X1 U1701 ( .A(n8678), .B(n5179), .Y(n5178) );
  INVX1 U1702 ( .A(n5178), .Y(n167) );
  OR2X1 U1703 ( .A(n8701), .B(n8677), .Y(n5179) );
  OR2X1 U1704 ( .A(n10369), .B(n5182), .Y(n5180) );
  INVX1 U1705 ( .A(n5180), .Y(n168) );
  OR2X1 U1706 ( .A(n5181), .B(n10368), .Y(n5182) );
  OR2X1 U1707 ( .A(n9323), .B(n5187), .Y(n5185) );
  INVX1 U1708 ( .A(n5185), .Y(n169) );
  OR2X1 U1709 ( .A(n5186), .B(n10368), .Y(n5187) );
  OR2X1 U1710 ( .A(n6641), .B(n5190), .Y(n5188) );
  INVX1 U1711 ( .A(n5188), .Y(n170) );
  OR2X1 U1712 ( .A(n5189), .B(n7159), .Y(n5190) );
  OR2X1 U1713 ( .A(n7669), .B(n5193), .Y(n5191) );
  INVX1 U1714 ( .A(n5191), .Y(n171) );
  OR2X1 U1715 ( .A(n5192), .B(n8180), .Y(n5193) );
  OR2X1 U1716 ( .A(n8685), .B(n5196), .Y(n5194) );
  INVX1 U1717 ( .A(n5194), .Y(n172) );
  OR2X1 U1718 ( .A(n5195), .B(n9191), .Y(n5196) );
  OR2X1 U1719 ( .A(n9701), .B(n5199), .Y(n5197) );
  INVX1 U1720 ( .A(n5197), .Y(n173) );
  OR2X1 U1721 ( .A(n5198), .B(n10230), .Y(n5199) );
  OR2X1 U1722 ( .A(n8756), .B(n5202), .Y(n5200) );
  OR2X1 U1723 ( .A(n5201), .B(n8754), .Y(n5202) );
  OR2X1 U1724 ( .A(n9691), .B(n5204), .Y(n5203) );
  OR2X1 U1725 ( .A(n9692), .B(n9690), .Y(n5204) );
  OR2X1 U1726 ( .A(n7658), .B(n5206), .Y(n5205) );
  OR2X1 U1727 ( .A(n7659), .B(n7657), .Y(n5206) );
  OR2X1 U1728 ( .A(n6854), .B(n5209), .Y(n5208) );
  OR2X1 U1729 ( .A(n6920), .B(n6866), .Y(n5209) );
  OR2X1 U1730 ( .A(n7872), .B(n5211), .Y(n5210) );
  OR2X1 U1731 ( .A(n7873), .B(n7885), .Y(n5211) );
  OR2X1 U1732 ( .A(n9918), .B(n5213), .Y(n5212) );
  OR2X1 U1733 ( .A(n9917), .B(n9930), .Y(n5213) );
  OR2X1 U1734 ( .A(n9331), .B(n5219), .Y(n5217) );
  OR2X1 U1735 ( .A(n5218), .B(n10381), .Y(n5219) );
  OR2X1 U1736 ( .A(n10382), .B(n5222), .Y(n5220) );
  OR2X1 U1737 ( .A(n5221), .B(n10381), .Y(n5222) );
  OR2X1 U1738 ( .A(n9329), .B(n5225), .Y(n5223) );
  OR2X1 U1739 ( .A(n5224), .B(n10378), .Y(n5225) );
  OR2X1 U1740 ( .A(n7297), .B(n5228), .Y(n5226) );
  OR2X1 U1741 ( .A(n5227), .B(n10368), .Y(n5228) );
  OR2X1 U1742 ( .A(n8313), .B(n5231), .Y(n5229) );
  OR2X1 U1743 ( .A(n5230), .B(n10368), .Y(n5231) );
  OR2X1 U1744 ( .A(n9785), .B(n5234), .Y(n5232) );
  OR2X1 U1745 ( .A(n5233), .B(n9783), .Y(n5234) );
  OR2X1 U1746 ( .A(n7303), .B(n5241), .Y(n5239) );
  OR2X1 U1747 ( .A(n5240), .B(n10378), .Y(n5241) );
  OR2X1 U1748 ( .A(n7305), .B(n5244), .Y(n5242) );
  OR2X1 U1749 ( .A(n5243), .B(n10381), .Y(n5244) );
  OR2X1 U1750 ( .A(n7749), .B(n5247), .Y(n5245) );
  OR2X1 U1751 ( .A(n5246), .B(n7747), .Y(n5247) );
  OR2X1 U1752 ( .A(n8319), .B(n5250), .Y(n5248) );
  OR2X1 U1753 ( .A(n5249), .B(n10378), .Y(n5250) );
  OR2X1 U1754 ( .A(n8321), .B(n5253), .Y(n5251) );
  OR2X1 U1755 ( .A(n5252), .B(n10381), .Y(n5253) );
  OR2X1 U1756 ( .A(n8879), .B(n5257), .Y(n5256) );
  OR2X1 U1757 ( .A(n8946), .B(n8891), .Y(n5257) );
  OR2X1 U1758 ( .A(n6629), .B(n5259), .Y(n5258) );
  OR2X1 U1759 ( .A(n6630), .B(n6628), .Y(n5259) );
  OR2X1 U1760 ( .A(n6724), .B(n5262), .Y(n5260) );
  OR2X1 U1761 ( .A(n5261), .B(n6720), .Y(n5262) );
  AND2X1 U1762 ( .A(n1949), .B(n1942), .Y(mult32_B[31]) );
  INVX1 U1763 ( .A(mult32_B[31]), .Y(n174) );
  AND2X1 U1764 ( .A(n1951), .B(n1943), .Y(mult32_B[0]) );
  INVX1 U1765 ( .A(mult32_B[0]), .Y(n175) );
  AND2X1 U1766 ( .A(n6286), .B(n6079), .Y(n6486) );
  AND2X1 U1767 ( .A(n6286), .B(n6081), .Y(n6583) );
  AND2X1 U1768 ( .A(n1051), .B(n6129), .Y(n6604) );
  AND2X1 U1769 ( .A(n5820), .B(n5912), .Y(n6629) );
  AND2X1 U1770 ( .A(n6579), .B(n6286), .Y(n6641) );
  AND2X1 U1771 ( .A(n6551), .B(n5934), .Y(n6661) );
  AND2X1 U1772 ( .A(n1052), .B(n6129), .Y(n6682) );
  AND2X1 U1773 ( .A(n6290), .B(n6080), .Y(n6707) );
  AND2X1 U1774 ( .A(n6579), .B(n6288), .Y(n6710) );
  OR2X1 U1775 ( .A(n6713), .B(n6712), .Y(n6714) );
  AND2X1 U1776 ( .A(n6277), .B(n6065), .Y(n6737) );
  AND2X1 U1777 ( .A(n5948), .B(n6730), .Y(n6788) );
  AND2X1 U1778 ( .A(n5912), .B(n9853), .Y(n6794) );
  AND2X1 U1779 ( .A(n6551), .B(n6273), .Y(n6850) );
  AND2X1 U1780 ( .A(n6866), .B(n4866), .Y(n6870) );
  AND2X1 U1781 ( .A(n526), .B(n5849), .Y(n6887) );
  AND2X1 U1782 ( .A(n67), .B(n6081), .Y(n6911) );
  AND2X1 U1783 ( .A(n67), .B(n6080), .Y(n6963) );
  AND2X1 U1784 ( .A(n5949), .B(n6975), .Y(n6978) );
  AND2X1 U1785 ( .A(n1105), .B(n6127), .Y(n6989) );
  AND2X1 U1786 ( .A(n6282), .B(n9632), .Y(n7012) );
  AND2X1 U1787 ( .A(n5214), .B(n10087), .Y(n7033) );
  AND2X1 U1788 ( .A(n1106), .B(n6127), .Y(n7046) );
  AND2X1 U1789 ( .A(n5764), .B(n7360), .Y(n7078) );
  AND2X1 U1790 ( .A(n5944), .B(n9500), .Y(n7114) );
  AND2X1 U1791 ( .A(n1798), .B(n5777), .Y(n7117) );
  AND2X1 U1792 ( .A(n5764), .B(n5704), .Y(n7144) );
  AND2X1 U1793 ( .A(n6173), .B(n7152), .Y(n7153) );
  AND2X1 U1794 ( .A(n1060), .B(n6129), .Y(n7192) );
  AND2X1 U1795 ( .A(n5013), .B(n6073), .Y(n7245) );
  AND2X1 U1796 ( .A(n1109), .B(n6127), .Y(n7256) );
  AND2X1 U1797 ( .A(n6627), .B(n6579), .Y(n7297) );
  AND2X1 U1798 ( .A(n5820), .B(n6627), .Y(n7303) );
  AND2X1 U1799 ( .A(n6551), .B(n6627), .Y(n7305) );
  AND2X1 U1800 ( .A(n5911), .B(n5735), .Y(n7320) );
  AND2X1 U1801 ( .A(n6018), .B(n10502), .Y(n7382) );
  AND2X1 U1802 ( .A(n1802), .B(n5777), .Y(n7385) );
  AND2X1 U1803 ( .A(n6303), .B(n6080), .Y(n7530) );
  AND2X1 U1804 ( .A(n6303), .B(n6081), .Y(n7615) );
  AND2X1 U1805 ( .A(n1035), .B(n6129), .Y(n7635) );
  AND2X1 U1806 ( .A(n5767), .B(n5952), .Y(n7658) );
  AND2X1 U1807 ( .A(n7611), .B(n6303), .Y(n7669) );
  AND2X1 U1808 ( .A(n7586), .B(n5975), .Y(n7690) );
  AND2X1 U1809 ( .A(n10502), .B(n6029), .Y(n7708) );
  AND2X1 U1810 ( .A(n1036), .B(n6129), .Y(n7711) );
  AND2X1 U1811 ( .A(n6308), .B(n6080), .Y(n7734) );
  AND2X1 U1812 ( .A(n7611), .B(n6305), .Y(n7737) );
  OR2X1 U1813 ( .A(n7740), .B(n7739), .Y(n7741) );
  AND2X1 U1814 ( .A(n1294), .B(n6125), .Y(n7773) );
  AND2X1 U1815 ( .A(n5953), .B(n6080), .Y(n7799) );
  AND2X1 U1816 ( .A(n5951), .B(n9853), .Y(n7813) );
  AND2X1 U1817 ( .A(n1118), .B(n5826), .Y(n7823) );
  AND2X1 U1818 ( .A(n7586), .B(n5957), .Y(n7868) );
  AND2X1 U1819 ( .A(n7885), .B(n4867), .Y(n7889) );
  AND2X1 U1820 ( .A(n2252), .B(n5838), .Y(n7917) );
  AND2X1 U1821 ( .A(n5964), .B(n6081), .Y(n7941) );
  AND2X1 U1822 ( .A(n7985), .B(n5056), .Y(n7948) );
  AND2X1 U1823 ( .A(n5965), .B(n5800), .Y(n7979) );
  AND2X1 U1824 ( .A(n5989), .B(n7989), .Y(n7992) );
  AND2X1 U1825 ( .A(n1121), .B(n5826), .Y(n8002) );
  AND2X1 U1826 ( .A(n6297), .B(n9632), .Y(n8025) );
  AND2X1 U1827 ( .A(n5215), .B(n10087), .Y(n8046) );
  AND2X1 U1828 ( .A(n1122), .B(n5826), .Y(n8059) );
  AND2X1 U1829 ( .A(n6626), .B(n5712), .Y(n8134) );
  AND2X1 U1830 ( .A(n5796), .B(n5205), .Y(n8169) );
  AND2X1 U1831 ( .A(n5651), .B(n10505), .Y(n8177) );
  AND2X1 U1832 ( .A(n9688), .B(n6302), .Y(n8188) );
  AND2X1 U1833 ( .A(n1301), .B(n6125), .Y(n8208) );
  AND2X1 U1834 ( .A(n5016), .B(n6073), .Y(n8259) );
  AND2X1 U1835 ( .A(n1302), .B(n6125), .Y(n8273) );
  AND2X1 U1836 ( .A(n7656), .B(n7611), .Y(n8313) );
  AND2X1 U1837 ( .A(n5767), .B(n7656), .Y(n8319) );
  AND2X1 U1838 ( .A(n7586), .B(n7656), .Y(n8321) );
  AND2X1 U1839 ( .A(n5951), .B(n5735), .Y(n8336) );
  AND2X1 U1840 ( .A(n6354), .B(n10502), .Y(n8396) );
  AND2X1 U1841 ( .A(n1786), .B(n5777), .Y(n8399) );
  AND2X1 U1842 ( .A(n1019), .B(n6129), .Y(n8637) );
  AND2X1 U1843 ( .A(n5768), .B(n5880), .Y(n8678) );
  AND2X1 U1844 ( .A(n1020), .B(n5786), .Y(n8713) );
  AND2X1 U1845 ( .A(n8588), .B(n6330), .Y(n8716) );
  AND2X1 U1846 ( .A(n6337), .B(n6080), .Y(n8741) );
  AND2X1 U1847 ( .A(n8610), .B(n5286), .Y(n8744) );
  OR2X1 U1848 ( .A(n8747), .B(n8746), .Y(n8748) );
  AND2X1 U1849 ( .A(n6319), .B(n6065), .Y(n8766) );
  AND2X1 U1850 ( .A(n1278), .B(n6125), .Y(n8780) );
  AND2X1 U1851 ( .A(n6730), .B(n6024), .Y(n8817) );
  AND2X1 U1852 ( .A(n5880), .B(n9853), .Y(n8820) );
  AND2X1 U1853 ( .A(n1070), .B(n5826), .Y(n8830) );
  AND2X1 U1854 ( .A(n8588), .B(n5995), .Y(n8875) );
  AND2X1 U1855 ( .A(n8891), .B(n4868), .Y(n8895) );
  AND2X1 U1856 ( .A(n494), .B(n5849), .Y(n8913) );
  AND2X1 U1857 ( .A(n43), .B(n9626), .Y(n8937) );
  AND2X1 U1858 ( .A(n43), .B(n6080), .Y(n8991) );
  AND2X1 U1859 ( .A(n5271), .B(n9000), .Y(n9003) );
  AND2X1 U1860 ( .A(n1073), .B(n6127), .Y(n9013) );
  AND2X1 U1861 ( .A(n6325), .B(n9632), .Y(n9036) );
  AND2X1 U1862 ( .A(n5216), .B(n10087), .Y(n9057) );
  AND2X1 U1863 ( .A(n1074), .B(n6127), .Y(n9070) );
  AND2X1 U1864 ( .A(n6626), .B(n5714), .Y(n9146) );
  AND2X1 U1865 ( .A(n9460), .B(n5178), .Y(n9181) );
  AND2X1 U1866 ( .A(n5579), .B(n10505), .Y(n9188) );
  AND2X1 U1867 ( .A(n5019), .B(n6073), .Y(n9270) );
  AND2X1 U1868 ( .A(n1286), .B(n6125), .Y(n9284) );
  AND2X1 U1869 ( .A(n8679), .B(n8610), .Y(n9323) );
  AND2X1 U1870 ( .A(n8679), .B(n5768), .Y(n9329) );
  AND2X1 U1871 ( .A(n6217), .B(n6151), .Y(n5768) );
  AND2X1 U1872 ( .A(n8679), .B(n8588), .Y(n9331) );
  AND2X1 U1873 ( .A(n5991), .B(n5735), .Y(n9346) );
  AND2X1 U1874 ( .A(n5945), .B(n10502), .Y(n9406) );
  AND2X1 U1875 ( .A(n3143), .B(n5776), .Y(n9439) );
  AND2X1 U1876 ( .A(n1819), .B(n5783), .Y(n9446) );
  AND2X1 U1877 ( .A(n5286), .B(n5217), .Y(n9494) );
  AND2X1 U1878 ( .A(n5805), .B(n5200), .Y(n9504) );
  AND2X1 U1879 ( .A(n1003), .B(n6129), .Y(n9667) );
  AND2X1 U1880 ( .A(n59), .B(n5769), .Y(n9691) );
  AND2X1 U1881 ( .A(n6347), .B(n9614), .Y(n9724) );
  AND2X1 U1882 ( .A(n5958), .B(n10502), .Y(n9743) );
  AND2X1 U1883 ( .A(n1004), .B(n6129), .Y(n9746) );
  AND2X1 U1884 ( .A(n5800), .B(n6356), .Y(n9769) );
  AND2X1 U1885 ( .A(n6055), .B(n9639), .Y(n9772) );
  OR2X1 U1886 ( .A(n9776), .B(n9775), .Y(n9777) );
  AND2X1 U1887 ( .A(n6034), .B(n6065), .Y(n9799) );
  AND2X1 U1888 ( .A(n1262), .B(n6125), .Y(n9814) );
  AND2X1 U1889 ( .A(n59), .B(n9853), .Y(n9856) );
  AND2X1 U1890 ( .A(n1086), .B(n6127), .Y(n9866) );
  AND2X1 U1891 ( .A(n9930), .B(n4869), .Y(n9934) );
  AND2X1 U1892 ( .A(n10030), .B(n5050), .Y(n9994) );
  AND2X1 U1893 ( .A(n6060), .B(n10035), .Y(n10038) );
  AND2X1 U1894 ( .A(n1089), .B(n6127), .Y(n10048) );
  AND2X1 U1895 ( .A(n6345), .B(n6077), .Y(n10071) );
  AND2X1 U1896 ( .A(n10087), .B(n5207), .Y(n10096) );
  AND2X1 U1897 ( .A(n1090), .B(n6127), .Y(n10110) );
  AND2X1 U1898 ( .A(n6626), .B(n5713), .Y(n10186) );
  AND2X1 U1899 ( .A(n5797), .B(n5203), .Y(n10220) );
  AND2X1 U1900 ( .A(n5584), .B(n10505), .Y(n10227) );
  AND2X1 U1901 ( .A(n5022), .B(n6073), .Y(n10312) );
  AND2X1 U1902 ( .A(n9689), .B(n9639), .Y(n10369) );
  AND2X1 U1903 ( .A(n5769), .B(n9689), .Y(n10379) );
  AND2X1 U1904 ( .A(n9614), .B(n9689), .Y(n10382) );
  AND2X1 U1905 ( .A(n5735), .B(n59), .Y(n10398) );
  AND2X1 U1906 ( .A(n10506), .B(n10505), .Y(n10509) );
  AND2X1 U1907 ( .A(n10498), .B(n4863), .Y(n10577) );
  INVX1 U1908 ( .A(n6368), .Y(n176) );
  INVX1 U1909 ( .A(n176), .Y(n177) );
  BUFX2 U1910 ( .A(n6370), .Y(n178) );
  BUFX2 U1911 ( .A(n6372), .Y(n179) );
  BUFX2 U1912 ( .A(n6374), .Y(n180) );
  BUFX2 U1913 ( .A(n6376), .Y(n181) );
  BUFX2 U1914 ( .A(n6378), .Y(n182) );
  BUFX2 U1915 ( .A(n6380), .Y(n183) );
  BUFX2 U1916 ( .A(n6382), .Y(n184) );
  BUFX2 U1917 ( .A(n6388), .Y(n185) );
  BUFX2 U1918 ( .A(n6390), .Y(n186) );
  BUFX2 U1919 ( .A(n6392), .Y(n187) );
  INVX1 U1920 ( .A(n6394), .Y(n188) );
  INVX1 U1921 ( .A(n188), .Y(n189) );
  INVX1 U1922 ( .A(n6396), .Y(n190) );
  INVX1 U1923 ( .A(n190), .Y(n191) );
  BUFX2 U1924 ( .A(n6398), .Y(n192) );
  BUFX2 U1925 ( .A(n6404), .Y(n193) );
  BUFX2 U1926 ( .A(n6406), .Y(n194) );
  BUFX2 U1927 ( .A(n6408), .Y(n195) );
  BUFX2 U1928 ( .A(n6410), .Y(n196) );
  BUFX2 U1929 ( .A(n6412), .Y(n197) );
  INVX1 U1930 ( .A(n6414), .Y(n198) );
  INVX1 U1931 ( .A(n198), .Y(n199) );
  BUFX2 U1932 ( .A(n6418), .Y(n200) );
  BUFX2 U1933 ( .A(n6420), .Y(n201) );
  BUFX2 U1934 ( .A(n6424), .Y(n202) );
  BUFX2 U1935 ( .A(n6426), .Y(n203) );
  BUFX2 U1936 ( .A(n6474), .Y(n204) );
  BUFX2 U1937 ( .A(n6482), .Y(n205) );
  BUFX2 U1938 ( .A(n6492), .Y(n206) );
  BUFX2 U1939 ( .A(n6504), .Y(n207) );
  BUFX2 U1940 ( .A(n6501), .Y(n208) );
  BUFX2 U1941 ( .A(n6512), .Y(n209) );
  BUFX2 U1942 ( .A(n6523), .Y(n210) );
  BUFX2 U1943 ( .A(n6528), .Y(n211) );
  BUFX2 U1944 ( .A(n6530), .Y(n212) );
  BUFX2 U1945 ( .A(n6537), .Y(n213) );
  BUFX2 U1946 ( .A(n6554), .Y(n214) );
  BUFX2 U1947 ( .A(n6574), .Y(n215) );
  BUFX2 U1948 ( .A(n6602), .Y(n216) );
  BUFX2 U1949 ( .A(n6620), .Y(n217) );
  BUFX2 U1950 ( .A(n6691), .Y(n218) );
  BUFX2 U1951 ( .A(n6698), .Y(n219) );
  BUFX2 U1952 ( .A(n6718), .Y(n220) );
  BUFX2 U1953 ( .A(n6729), .Y(n221) );
  BUFX2 U1954 ( .A(n6744), .Y(n222) );
  BUFX2 U1955 ( .A(n6749), .Y(n223) );
  BUFX2 U1956 ( .A(n6759), .Y(n224) );
  BUFX2 U1957 ( .A(n6766), .Y(n225) );
  BUFX2 U1958 ( .A(n6771), .Y(n226) );
  BUFX2 U1959 ( .A(n6785), .Y(n227) );
  BUFX2 U1960 ( .A(n6797), .Y(n228) );
  BUFX2 U1961 ( .A(n6807), .Y(n229) );
  BUFX2 U1962 ( .A(n6815), .Y(n230) );
  BUFX2 U1963 ( .A(n6822), .Y(n231) );
  BUFX2 U1964 ( .A(n6827), .Y(n232) );
  BUFX2 U1965 ( .A(n6845), .Y(n233) );
  BUFX2 U1966 ( .A(n6860), .Y(n234) );
  BUFX2 U1967 ( .A(n6865), .Y(n235) );
  BUFX2 U1968 ( .A(n6878), .Y(n236) );
  BUFX2 U1969 ( .A(n6890), .Y(n237) );
  BUFX2 U1970 ( .A(n6892), .Y(n238) );
  BUFX2 U1971 ( .A(n6905), .Y(n239) );
  BUFX2 U1972 ( .A(n6957), .Y(n240) );
  BUFX2 U1973 ( .A(n6970), .Y(n241) );
  BUFX2 U1974 ( .A(n6981), .Y(n242) );
  BUFX2 U1975 ( .A(n6998), .Y(n243) );
  BUFX2 U1976 ( .A(n7005), .Y(n244) );
  BUFX2 U1977 ( .A(n7018), .Y(n245) );
  BUFX2 U1978 ( .A(n7024), .Y(n246) );
  BUFX2 U1979 ( .A(n7029), .Y(n247) );
  BUFX2 U1980 ( .A(n7037), .Y(n248) );
  BUFX2 U1981 ( .A(n7049), .Y(n249) );
  BUFX2 U1982 ( .A(n7055), .Y(n250) );
  BUFX2 U1983 ( .A(n7062), .Y(n251) );
  BUFX2 U1984 ( .A(n7125), .Y(n252) );
  BUFX2 U1985 ( .A(n7137), .Y(n253) );
  BUFX2 U1986 ( .A(n7200), .Y(n254) );
  BUFX2 U1987 ( .A(n7217), .Y(n255) );
  BUFX2 U1988 ( .A(n7232), .Y(n256) );
  BUFX2 U1989 ( .A(n7249), .Y(n257) );
  BUFX2 U1990 ( .A(n7259), .Y(n258) );
  BUFX2 U1991 ( .A(n7266), .Y(n259) );
  BUFX2 U1992 ( .A(n7273), .Y(n260) );
  BUFX2 U1993 ( .A(n7278), .Y(n261) );
  BUFX2 U1994 ( .A(n7312), .Y(n262) );
  BUFX2 U1995 ( .A(n7317), .Y(n263) );
  BUFX2 U1996 ( .A(n7328), .Y(n264) );
  BUFX2 U1997 ( .A(n7335), .Y(n265) );
  BUFX2 U1998 ( .A(n7393), .Y(n266) );
  BUFX2 U1999 ( .A(n7400), .Y(n267) );
  BUFX2 U2000 ( .A(n7419), .Y(n268) );
  BUFX2 U2001 ( .A(n7459), .Y(n269) );
  BUFX2 U2002 ( .A(n7466), .Y(n270) );
  BUFX2 U2003 ( .A(n7471), .Y(n271) );
  BUFX2 U2004 ( .A(n7480), .Y(n272) );
  BUFX2 U2005 ( .A(n7498), .Y(n273) );
  BUFX2 U2006 ( .A(n7500), .Y(n274) );
  BUFX2 U2007 ( .A(n7511), .Y(n275) );
  BUFX2 U2008 ( .A(n7518), .Y(n276) );
  BUFX2 U2009 ( .A(n7526), .Y(n277) );
  BUFX2 U2010 ( .A(n7533), .Y(n278) );
  BUFX2 U2011 ( .A(n7543), .Y(n279) );
  BUFX2 U2012 ( .A(n7540), .Y(n280) );
  BUFX2 U2013 ( .A(n7546), .Y(n281) );
  BUFX2 U2014 ( .A(n7561), .Y(n282) );
  BUFX2 U2015 ( .A(n7563), .Y(n283) );
  BUFX2 U2016 ( .A(n7570), .Y(n284) );
  BUFX2 U2017 ( .A(n7577), .Y(n285) );
  BUFX2 U2018 ( .A(n7589), .Y(n286) );
  BUFX2 U2019 ( .A(n7606), .Y(n287) );
  BUFX2 U2020 ( .A(n7633), .Y(n288) );
  BUFX2 U2021 ( .A(n7644), .Y(n289) );
  BUFX2 U2022 ( .A(n7651), .Y(n290) );
  BUFX2 U2023 ( .A(n7719), .Y(n291) );
  BUFX2 U2024 ( .A(n7726), .Y(n292) );
  BUFX2 U2025 ( .A(n7745), .Y(n293) );
  BUFX2 U2026 ( .A(n7754), .Y(n294) );
  BUFX2 U2027 ( .A(n7766), .Y(n295) );
  BUFX2 U2028 ( .A(n7771), .Y(n296) );
  BUFX2 U2029 ( .A(n7781), .Y(n297) );
  BUFX2 U2030 ( .A(n7788), .Y(n298) );
  BUFX2 U2031 ( .A(n7793), .Y(n299) );
  BUFX2 U2032 ( .A(n7807), .Y(n300) );
  BUFX2 U2033 ( .A(n7816), .Y(n301) );
  BUFX2 U2034 ( .A(n7826), .Y(n302) );
  BUFX2 U2035 ( .A(n7832), .Y(n303) );
  BUFX2 U2036 ( .A(n7839), .Y(n304) );
  BUFX2 U2037 ( .A(n7844), .Y(n305) );
  BUFX2 U2038 ( .A(n7863), .Y(n306) );
  BUFX2 U2039 ( .A(n7879), .Y(n307) );
  BUFX2 U2040 ( .A(n7884), .Y(n308) );
  BUFX2 U2041 ( .A(n7897), .Y(n309) );
  BUFX2 U2042 ( .A(n7904), .Y(n310) );
  BUFX2 U2043 ( .A(n7960), .Y(n311) );
  BUFX2 U2044 ( .A(n7967), .Y(n312) );
  BUFX2 U2045 ( .A(n7973), .Y(n313) );
  BUFX2 U2046 ( .A(n7987), .Y(n314) );
  BUFX2 U2047 ( .A(n7995), .Y(n315) );
  BUFX2 U2048 ( .A(n8011), .Y(n316) );
  BUFX2 U2049 ( .A(n8018), .Y(n317) );
  BUFX2 U2050 ( .A(n8031), .Y(n318) );
  BUFX2 U2051 ( .A(n8037), .Y(n319) );
  BUFX2 U2052 ( .A(n8042), .Y(n320) );
  BUFX2 U2053 ( .A(n8050), .Y(n321) );
  BUFX2 U2054 ( .A(n8062), .Y(n322) );
  BUFX2 U2055 ( .A(n8068), .Y(n323) );
  BUFX2 U2056 ( .A(n8075), .Y(n324) );
  BUFX2 U2057 ( .A(n8129), .Y(n325) );
  BUFX2 U2058 ( .A(n8143), .Y(n326) );
  BUFX2 U2059 ( .A(n8150), .Y(n327) );
  BUFX2 U2060 ( .A(n8155), .Y(n328) );
  BUFX2 U2061 ( .A(n8186), .Y(n329) );
  BUFX2 U2062 ( .A(n8206), .Y(n330) );
  BUFX2 U2063 ( .A(n8217), .Y(n331) );
  BUFX2 U2064 ( .A(n8224), .Y(n332) );
  BUFX2 U2065 ( .A(n8234), .Y(n333) );
  BUFX2 U2066 ( .A(n8246), .Y(n334) );
  BUFX2 U2067 ( .A(n8266), .Y(n335) );
  BUFX2 U2068 ( .A(n8271), .Y(n336) );
  BUFX2 U2069 ( .A(n8281), .Y(n337) );
  BUFX2 U2070 ( .A(n8288), .Y(n338) );
  BUFX2 U2071 ( .A(n8293), .Y(n339) );
  BUFX2 U2072 ( .A(n8328), .Y(n340) );
  BUFX2 U2073 ( .A(n8333), .Y(n341) );
  BUFX2 U2074 ( .A(n8344), .Y(n342) );
  BUFX2 U2075 ( .A(n8407), .Y(n343) );
  BUFX2 U2076 ( .A(n8417), .Y(n344) );
  BUFX2 U2077 ( .A(n8428), .Y(n345) );
  BUFX2 U2078 ( .A(n8446), .Y(n346) );
  BUFX2 U2079 ( .A(n8458), .Y(n347) );
  BUFX2 U2080 ( .A(n8462), .Y(n348) );
  BUFX2 U2081 ( .A(n8478), .Y(n349) );
  BUFX2 U2082 ( .A(n8488), .Y(n350) );
  BUFX2 U2083 ( .A(n8503), .Y(n351) );
  BUFX2 U2084 ( .A(n8505), .Y(n352) );
  BUFX2 U2085 ( .A(n8522), .Y(n353) );
  BUFX2 U2086 ( .A(n8530), .Y(n354) );
  BUFX2 U2087 ( .A(n8537), .Y(n355) );
  BUFX2 U2088 ( .A(n8547), .Y(n356) );
  BUFX2 U2089 ( .A(n8544), .Y(n357) );
  BUFX2 U2090 ( .A(n8550), .Y(n358) );
  BUFX2 U2091 ( .A(n8560), .Y(n359) );
  BUFX2 U2092 ( .A(n8565), .Y(n616) );
  BUFX2 U2093 ( .A(n8567), .Y(n617) );
  BUFX2 U2094 ( .A(n8574), .Y(n618) );
  BUFX2 U2095 ( .A(n8591), .Y(n619) );
  BUFX2 U2096 ( .A(n8608), .Y(n620) );
  BUFX2 U2097 ( .A(n8635), .Y(n621) );
  BUFX2 U2098 ( .A(n8658), .Y(n622) );
  BUFX2 U2099 ( .A(n8660), .Y(n623) );
  BUFX2 U2100 ( .A(n8666), .Y(n624) );
  BUFX2 U2101 ( .A(n8673), .Y(n625) );
  BUFX2 U2102 ( .A(n8711), .Y(n626) );
  BUFX2 U2103 ( .A(n8732), .Y(n627) );
  BUFX2 U2104 ( .A(n8752), .Y(n628) );
  BUFX2 U2105 ( .A(n8761), .Y(n629) );
  BUFX2 U2106 ( .A(n8773), .Y(n630) );
  BUFX2 U2107 ( .A(n8778), .Y(n631) );
  BUFX2 U2108 ( .A(n8788), .Y(n632) );
  BUFX2 U2109 ( .A(n8795), .Y(n633) );
  BUFX2 U2110 ( .A(n8800), .Y(n634) );
  BUFX2 U2111 ( .A(n8814), .Y(n635) );
  BUFX2 U2112 ( .A(n8823), .Y(n636) );
  BUFX2 U2113 ( .A(n8833), .Y(n637) );
  BUFX2 U2114 ( .A(n8840), .Y(n638) );
  BUFX2 U2115 ( .A(n8847), .Y(n639) );
  BUFX2 U2116 ( .A(n8852), .Y(n640) );
  BUFX2 U2117 ( .A(n8870), .Y(n641) );
  BUFX2 U2118 ( .A(n8885), .Y(n642) );
  BUFX2 U2119 ( .A(n8890), .Y(n643) );
  BUFX2 U2120 ( .A(n8903), .Y(n644) );
  BUFX2 U2121 ( .A(n8916), .Y(n645) );
  BUFX2 U2122 ( .A(n8918), .Y(n646) );
  BUFX2 U2123 ( .A(n8931), .Y(n647) );
  BUFX2 U2124 ( .A(n8980), .Y(n648) );
  BUFX2 U2125 ( .A(n8985), .Y(n649) );
  BUFX2 U2126 ( .A(n8998), .Y(n650) );
  BUFX2 U2127 ( .A(n9006), .Y(n651) );
  BUFX2 U2128 ( .A(n9016), .Y(n652) );
  BUFX2 U2129 ( .A(n9022), .Y(n653) );
  BUFX2 U2130 ( .A(n9029), .Y(n654) );
  BUFX2 U2131 ( .A(n9042), .Y(n655) );
  BUFX2 U2132 ( .A(n9048), .Y(n656) );
  BUFX2 U2133 ( .A(n9053), .Y(n657) );
  BUFX2 U2134 ( .A(n9061), .Y(n658) );
  BUFX2 U2135 ( .A(n9073), .Y(n659) );
  BUFX2 U2136 ( .A(n9080), .Y(n660) );
  BUFX2 U2137 ( .A(n9087), .Y(n661) );
  BUFX2 U2138 ( .A(n9141), .Y(n662) );
  BUFX2 U2139 ( .A(n9155), .Y(n663) );
  BUFX2 U2140 ( .A(n9162), .Y(n664) );
  BUFX2 U2141 ( .A(n9167), .Y(n665) );
  BUFX2 U2142 ( .A(n9197), .Y(n666) );
  BUFX2 U2143 ( .A(n9217), .Y(n667) );
  BUFX2 U2144 ( .A(n9229), .Y(n668) );
  BUFX2 U2145 ( .A(n9236), .Y(n669) );
  BUFX2 U2146 ( .A(n9246), .Y(n670) );
  BUFX2 U2147 ( .A(n9257), .Y(n671) );
  BUFX2 U2148 ( .A(n9277), .Y(n672) );
  BUFX2 U2149 ( .A(n9282), .Y(n673) );
  BUFX2 U2150 ( .A(n9291), .Y(n674) );
  BUFX2 U2151 ( .A(n9298), .Y(n675) );
  BUFX2 U2152 ( .A(n9303), .Y(n676) );
  BUFX2 U2153 ( .A(n9338), .Y(n677) );
  BUFX2 U2154 ( .A(n9343), .Y(n678) );
  BUFX2 U2155 ( .A(n9354), .Y(n679) );
  BUFX2 U2156 ( .A(n9361), .Y(n680) );
  BUFX2 U2157 ( .A(n9418), .Y(n937) );
  BUFX2 U2158 ( .A(n9432), .Y(n938) );
  BUFX2 U2159 ( .A(n9437), .Y(n939) );
  BUFX2 U2160 ( .A(n9449), .Y(n940) );
  BUFX2 U2161 ( .A(n9463), .Y(n941) );
  BUFX2 U2162 ( .A(n9488), .Y(n942) );
  BUFX2 U2163 ( .A(n9538), .Y(n943) );
  BUFX2 U2164 ( .A(n9545), .Y(n944) );
  BUFX2 U2165 ( .A(n9553), .Y(n945) );
  BUFX2 U2166 ( .A(n9560), .Y(n946) );
  BUFX2 U2167 ( .A(n9570), .Y(n947) );
  BUFX2 U2168 ( .A(n9567), .Y(n948) );
  BUFX2 U2169 ( .A(n9573), .Y(n949) );
  INVX1 U2170 ( .A(n9583), .Y(n950) );
  INVX1 U2171 ( .A(n950), .Y(n951) );
  BUFX2 U2172 ( .A(n9588), .Y(n952) );
  BUFX2 U2173 ( .A(n9590), .Y(n953) );
  BUFX2 U2174 ( .A(n9598), .Y(n954) );
  BUFX2 U2175 ( .A(n9605), .Y(n955) );
  BUFX2 U2176 ( .A(n9617), .Y(n956) );
  BUFX2 U2177 ( .A(n9637), .Y(n957) );
  BUFX2 U2178 ( .A(n9665), .Y(n958) );
  BUFX2 U2179 ( .A(n9676), .Y(n959) );
  BUFX2 U2180 ( .A(n9683), .Y(n960) );
  BUFX2 U2181 ( .A(n9754), .Y(n961) );
  BUFX2 U2182 ( .A(n9761), .Y(n962) );
  BUFX2 U2183 ( .A(n9781), .Y(n963) );
  BUFX2 U2184 ( .A(n9790), .Y(n964) );
  BUFX2 U2185 ( .A(n9807), .Y(n965) );
  BUFX2 U2186 ( .A(n9812), .Y(n966) );
  BUFX2 U2187 ( .A(n9822), .Y(n967) );
  BUFX2 U2188 ( .A(n9829), .Y(n968) );
  BUFX2 U2189 ( .A(n9834), .Y(n969) );
  BUFX2 U2190 ( .A(n9849), .Y(n970) );
  BUFX2 U2191 ( .A(n9859), .Y(n971) );
  BUFX2 U2192 ( .A(n9869), .Y(n972) );
  BUFX2 U2193 ( .A(n9876), .Y(n973) );
  BUFX2 U2194 ( .A(n9883), .Y(n974) );
  BUFX2 U2195 ( .A(n9888), .Y(n975) );
  BUFX2 U2196 ( .A(n9907), .Y(n976) );
  BUFX2 U2197 ( .A(n9924), .Y(n977) );
  BUFX2 U2198 ( .A(n9929), .Y(n978) );
  BUFX2 U2199 ( .A(n9942), .Y(n979) );
  BUFX2 U2200 ( .A(n9949), .Y(n980) );
  BUFX2 U2201 ( .A(n10006), .Y(n981) );
  BUFX2 U2202 ( .A(n10013), .Y(n982) );
  BUFX2 U2203 ( .A(n10019), .Y(n983) );
  BUFX2 U2204 ( .A(n10032), .Y(n984) );
  BUFX2 U2205 ( .A(n10041), .Y(n985) );
  BUFX2 U2206 ( .A(n10051), .Y(n986) );
  BUFX2 U2207 ( .A(n10057), .Y(n987) );
  BUFX2 U2208 ( .A(n10064), .Y(n988) );
  BUFX2 U2209 ( .A(n10078), .Y(n989) );
  BUFX2 U2210 ( .A(n10084), .Y(n990) );
  BUFX2 U2211 ( .A(n10091), .Y(n991) );
  BUFX2 U2212 ( .A(n10100), .Y(n992) );
  BUFX2 U2213 ( .A(n10113), .Y(n993) );
  BUFX2 U2214 ( .A(n10120), .Y(n994) );
  BUFX2 U2215 ( .A(n10127), .Y(n995) );
  BUFX2 U2216 ( .A(n10181), .Y(n996) );
  BUFX2 U2217 ( .A(n10195), .Y(n997) );
  BUFX2 U2218 ( .A(n10202), .Y(n998) );
  BUFX2 U2219 ( .A(n10207), .Y(n999) );
  BUFX2 U2220 ( .A(n10236), .Y(n1000) );
  BUFX2 U2221 ( .A(n10257), .Y(n1001) );
  BUFX2 U2222 ( .A(n10269), .Y(n1130) );
  BUFX2 U2223 ( .A(n10276), .Y(n1131) );
  BUFX2 U2224 ( .A(n10286), .Y(n1132) );
  BUFX2 U2225 ( .A(n10299), .Y(n1133) );
  BUFX2 U2226 ( .A(n10320), .Y(n1134) );
  BUFX2 U2227 ( .A(n10325), .Y(n1135) );
  BUFX2 U2228 ( .A(n10336), .Y(n1136) );
  BUFX2 U2229 ( .A(n10343), .Y(n1137) );
  BUFX2 U2230 ( .A(n10390), .Y(n1138) );
  BUFX2 U2231 ( .A(n10395), .Y(n1139) );
  BUFX2 U2232 ( .A(n10406), .Y(n1140) );
  BUFX2 U2233 ( .A(n10473), .Y(n1141) );
  BUFX2 U2234 ( .A(n10586), .Y(n1142) );
  BUFX2 U2235 ( .A(n10588), .Y(n1143) );
  BUFX2 U2236 ( .A(n6632), .Y(n1144) );
  BUFX2 U2237 ( .A(n6646), .Y(n1145) );
  BUFX2 U2238 ( .A(n6950), .Y(n1146) );
  BUFX2 U2239 ( .A(n7041), .Y(n1147) );
  BUFX2 U2240 ( .A(n7432), .Y(n1148) );
  BUFX2 U2241 ( .A(n7661), .Y(n1149) );
  BUFX2 U2242 ( .A(n7674), .Y(n1150) );
  BUFX2 U2243 ( .A(n8054), .Y(n1151) );
  BUFX2 U2244 ( .A(n8119), .Y(n1152) );
  BUFX2 U2245 ( .A(n8730), .Y(n1153) );
  BUFX2 U2246 ( .A(n8978), .Y(n1154) );
  BUFX2 U2247 ( .A(n9065), .Y(n1155) );
  BUFX2 U2248 ( .A(n9131), .Y(n1156) );
  BUFX2 U2249 ( .A(n9694), .Y(n1157) );
  BUFX2 U2250 ( .A(n9707), .Y(n1158) );
  BUFX2 U2251 ( .A(n10105), .Y(n1159) );
  BUFX2 U2252 ( .A(n10171), .Y(n1160) );
  AND2X1 U2253 ( .A(n6076), .B(n5276), .Y(n6437) );
  INVX1 U2254 ( .A(n6437), .Y(n1161) );
  AND2X1 U2255 ( .A(n6076), .B(n43), .Y(n6439) );
  INVX1 U2256 ( .A(n6439), .Y(n1162) );
  OR2X1 U2257 ( .A(n8690), .B(n2340), .Y(n8709) );
  INVX1 U2258 ( .A(n8709), .Y(n1163) );
  BUFX2 U2259 ( .A(n6367), .Y(n1164) );
  BUFX2 U2260 ( .A(n6369), .Y(n1165) );
  BUFX2 U2261 ( .A(n6371), .Y(n1166) );
  BUFX2 U2262 ( .A(n6373), .Y(n1167) );
  BUFX2 U2263 ( .A(n6375), .Y(n1168) );
  BUFX2 U2264 ( .A(n6377), .Y(n1169) );
  BUFX2 U2265 ( .A(n6379), .Y(n1170) );
  BUFX2 U2266 ( .A(n6381), .Y(n1171) );
  BUFX2 U2267 ( .A(n6383), .Y(n1172) );
  BUFX2 U2268 ( .A(n6385), .Y(n1173) );
  BUFX2 U2269 ( .A(n6387), .Y(n1174) );
  INVX1 U2270 ( .A(n6389), .Y(n1175) );
  INVX1 U2271 ( .A(n1175), .Y(n1176) );
  BUFX2 U2272 ( .A(n6391), .Y(n1177) );
  BUFX2 U2273 ( .A(n6395), .Y(n1178) );
  BUFX2 U2274 ( .A(n6397), .Y(n1179) );
  BUFX2 U2275 ( .A(n6399), .Y(n1180) );
  BUFX2 U2276 ( .A(n6403), .Y(n1181) );
  BUFX2 U2277 ( .A(n6405), .Y(n1182) );
  BUFX2 U2278 ( .A(n6407), .Y(n1183) );
  BUFX2 U2279 ( .A(n6409), .Y(n1184) );
  BUFX2 U2280 ( .A(n6411), .Y(n1185) );
  BUFX2 U2281 ( .A(n6413), .Y(n1186) );
  BUFX2 U2282 ( .A(n6415), .Y(n1187) );
  BUFX2 U2283 ( .A(n6417), .Y(n1188) );
  BUFX2 U2284 ( .A(n6419), .Y(n1189) );
  BUFX2 U2285 ( .A(n6421), .Y(n1190) );
  BUFX2 U2286 ( .A(n6423), .Y(n1191) );
  BUFX2 U2287 ( .A(n6425), .Y(n1192) );
  BUFX2 U2288 ( .A(n6481), .Y(n1193) );
  BUFX2 U2289 ( .A(n6491), .Y(n1194) );
  BUFX2 U2290 ( .A(n6500), .Y(n1195) );
  BUFX2 U2291 ( .A(n6503), .Y(n1196) );
  BUFX2 U2292 ( .A(n6511), .Y(n1197) );
  BUFX2 U2293 ( .A(n6527), .Y(n1198) );
  BUFX2 U2294 ( .A(n6529), .Y(n1199) );
  BUFX2 U2295 ( .A(n6553), .Y(n1200) );
  BUFX2 U2296 ( .A(n6573), .Y(n1201) );
  BUFX2 U2297 ( .A(n6601), .Y(n1202) );
  BUFX2 U2298 ( .A(n6645), .Y(n1203) );
  BUFX2 U2299 ( .A(n6717), .Y(n1204) );
  BUFX2 U2300 ( .A(n6728), .Y(n1205) );
  BUFX2 U2301 ( .A(n6770), .Y(n1206) );
  BUFX2 U2302 ( .A(n6784), .Y(n1207) );
  BUFX2 U2303 ( .A(n6796), .Y(n1208) );
  BUFX2 U2304 ( .A(n6806), .Y(n1209) );
  BUFX2 U2305 ( .A(n6826), .Y(n1210) );
  BUFX2 U2306 ( .A(n6844), .Y(n1211) );
  BUFX2 U2307 ( .A(n6859), .Y(n1212) );
  BUFX2 U2308 ( .A(n6864), .Y(n1213) );
  BUFX2 U2309 ( .A(n6891), .Y(n1214) );
  BUFX2 U2310 ( .A(n6904), .Y(n1215) );
  BUFX2 U2311 ( .A(n6956), .Y(n1216) );
  BUFX2 U2312 ( .A(n6969), .Y(n1217) );
  BUFX2 U2313 ( .A(n6980), .Y(n1218) );
  BUFX2 U2314 ( .A(n7017), .Y(n1219) );
  BUFX2 U2315 ( .A(n7023), .Y(n1220) );
  BUFX2 U2316 ( .A(n7028), .Y(n1221) );
  BUFX2 U2317 ( .A(n7036), .Y(n1222) );
  BUFX2 U2318 ( .A(n7136), .Y(n1223) );
  INVX1 U2319 ( .A(n7216), .Y(n1224) );
  INVX1 U2320 ( .A(n1224), .Y(n1225) );
  BUFX2 U2321 ( .A(n7223), .Y(n1226) );
  BUFX2 U2322 ( .A(n7231), .Y(n1227) );
  BUFX2 U2323 ( .A(n7248), .Y(n1228) );
  BUFX2 U2324 ( .A(n7258), .Y(n1229) );
  BUFX2 U2325 ( .A(n7277), .Y(n1230) );
  BUFX2 U2326 ( .A(n7311), .Y(n1231) );
  BUFX2 U2327 ( .A(n7316), .Y(n1232) );
  BUFX2 U2328 ( .A(n7479), .Y(n1233) );
  BUFX2 U2329 ( .A(n7499), .Y(n1234) );
  BUFX2 U2330 ( .A(n7525), .Y(n1235) );
  BUFX2 U2331 ( .A(n7532), .Y(n1236) );
  BUFX2 U2332 ( .A(n7539), .Y(n1237) );
  BUFX2 U2333 ( .A(n7542), .Y(n1238) );
  BUFX2 U2334 ( .A(n7545), .Y(n1239) );
  BUFX2 U2335 ( .A(n7560), .Y(n1240) );
  BUFX2 U2336 ( .A(n7562), .Y(n1241) );
  BUFX2 U2337 ( .A(n7588), .Y(n1242) );
  BUFX2 U2338 ( .A(n7605), .Y(n1243) );
  BUFX2 U2339 ( .A(n7632), .Y(n1244) );
  BUFX2 U2340 ( .A(n7673), .Y(n1245) );
  BUFX2 U2341 ( .A(n7744), .Y(n1246) );
  BUFX2 U2342 ( .A(n7753), .Y(n1247) );
  BUFX2 U2343 ( .A(n7770), .Y(n1248) );
  BUFX2 U2344 ( .A(n7792), .Y(n1249) );
  BUFX2 U2345 ( .A(n7806), .Y(n1250) );
  BUFX2 U2346 ( .A(n7815), .Y(n1251) );
  BUFX2 U2347 ( .A(n7825), .Y(n1252) );
  BUFX2 U2348 ( .A(n7843), .Y(n1253) );
  BUFX2 U2349 ( .A(n7862), .Y(n1254) );
  BUFX2 U2350 ( .A(n7878), .Y(n1255) );
  BUFX2 U2351 ( .A(n7883), .Y(n1256) );
  BUFX2 U2352 ( .A(n7972), .Y(n1257) );
  BUFX2 U2353 ( .A(n7986), .Y(n1258) );
  BUFX2 U2354 ( .A(n7994), .Y(n1387) );
  BUFX2 U2355 ( .A(n8004), .Y(n1388) );
  BUFX2 U2356 ( .A(n8030), .Y(n1389) );
  BUFX2 U2357 ( .A(n8036), .Y(n1390) );
  BUFX2 U2358 ( .A(n8041), .Y(n1391) );
  BUFX2 U2359 ( .A(n8049), .Y(n1392) );
  BUFX2 U2360 ( .A(n8061), .Y(n1393) );
  BUFX2 U2361 ( .A(n8118), .Y(n1394) );
  BUFX2 U2362 ( .A(n8128), .Y(n1395) );
  BUFX2 U2363 ( .A(n8154), .Y(n1396) );
  BUFX2 U2364 ( .A(n8185), .Y(n1397) );
  BUFX2 U2365 ( .A(n8205), .Y(n1398) );
  BUFX2 U2366 ( .A(n8233), .Y(n1399) );
  BUFX2 U2367 ( .A(n8245), .Y(n1400) );
  BUFX2 U2368 ( .A(n8270), .Y(n1401) );
  BUFX2 U2369 ( .A(n8292), .Y(n1402) );
  BUFX2 U2370 ( .A(n8327), .Y(n1403) );
  BUFX2 U2371 ( .A(n8332), .Y(n1404) );
  BUFX2 U2372 ( .A(n8416), .Y(n1405) );
  BUFX2 U2373 ( .A(n8427), .Y(n1406) );
  BUFX2 U2374 ( .A(n8445), .Y(n1407) );
  BUFX2 U2375 ( .A(n8461), .Y(n1408) );
  BUFX2 U2376 ( .A(n8487), .Y(n1409) );
  BUFX2 U2377 ( .A(n8529), .Y(n1410) );
  BUFX2 U2378 ( .A(n8536), .Y(n1411) );
  BUFX2 U2379 ( .A(n8543), .Y(n1412) );
  BUFX2 U2380 ( .A(n8546), .Y(n1413) );
  BUFX2 U2381 ( .A(n8549), .Y(n1414) );
  BUFX2 U2382 ( .A(n8564), .Y(n1415) );
  BUFX2 U2383 ( .A(n8566), .Y(n1416) );
  BUFX2 U2384 ( .A(n8590), .Y(n1417) );
  BUFX2 U2385 ( .A(n8607), .Y(n1418) );
  BUFX2 U2386 ( .A(n8634), .Y(n1419) );
  BUFX2 U2387 ( .A(n8751), .Y(n1420) );
  BUFX2 U2388 ( .A(n8760), .Y(n1421) );
  BUFX2 U2389 ( .A(n8799), .Y(n1422) );
  BUFX2 U2390 ( .A(n8813), .Y(n1423) );
  BUFX2 U2391 ( .A(n8822), .Y(n1424) );
  BUFX2 U2392 ( .A(n8851), .Y(n1425) );
  BUFX2 U2393 ( .A(n8869), .Y(n1426) );
  BUFX2 U2394 ( .A(n8884), .Y(n1427) );
  BUFX2 U2395 ( .A(n8889), .Y(n1428) );
  BUFX2 U2396 ( .A(n8917), .Y(n1429) );
  BUFX2 U2397 ( .A(n8930), .Y(n1430) );
  BUFX2 U2398 ( .A(n8984), .Y(n1431) );
  BUFX2 U2399 ( .A(n8997), .Y(n1432) );
  BUFX2 U2400 ( .A(n9005), .Y(n1433) );
  BUFX2 U2401 ( .A(n9041), .Y(n1434) );
  BUFX2 U2402 ( .A(n9047), .Y(n1435) );
  BUFX2 U2403 ( .A(n9052), .Y(n1436) );
  BUFX2 U2404 ( .A(n9060), .Y(n1437) );
  BUFX2 U2405 ( .A(n9130), .Y(n1438) );
  BUFX2 U2406 ( .A(n9140), .Y(n1439) );
  BUFX2 U2407 ( .A(n9166), .Y(n1440) );
  BUFX2 U2408 ( .A(n9196), .Y(n1441) );
  BUFX2 U2409 ( .A(n9245), .Y(n1442) );
  BUFX2 U2410 ( .A(n9256), .Y(n1443) );
  BUFX2 U2411 ( .A(n9281), .Y(n1444) );
  BUFX2 U2412 ( .A(n9302), .Y(n1445) );
  BUFX2 U2413 ( .A(n9337), .Y(n1446) );
  BUFX2 U2414 ( .A(n9342), .Y(n1447) );
  BUFX2 U2415 ( .A(n9431), .Y(n1448) );
  BUFX2 U2416 ( .A(n9462), .Y(n1449) );
  BUFX2 U2417 ( .A(n9552), .Y(n1450) );
  BUFX2 U2418 ( .A(n9559), .Y(n1451) );
  BUFX2 U2419 ( .A(n9566), .Y(n1452) );
  BUFX2 U2420 ( .A(n9569), .Y(n1453) );
  BUFX2 U2421 ( .A(n9572), .Y(n1454) );
  BUFX2 U2422 ( .A(n9587), .Y(n1455) );
  BUFX2 U2423 ( .A(n9589), .Y(n1456) );
  BUFX2 U2424 ( .A(n9616), .Y(n1457) );
  BUFX2 U2425 ( .A(n9636), .Y(n1458) );
  BUFX2 U2426 ( .A(n9664), .Y(n1459) );
  BUFX2 U2427 ( .A(n9706), .Y(n1460) );
  BUFX2 U2428 ( .A(n9780), .Y(n1461) );
  BUFX2 U2429 ( .A(n9789), .Y(n1462) );
  BUFX2 U2430 ( .A(n9811), .Y(n1463) );
  BUFX2 U2431 ( .A(n9833), .Y(n1464) );
  BUFX2 U2432 ( .A(n9848), .Y(n1465) );
  BUFX2 U2433 ( .A(n9858), .Y(n1466) );
  BUFX2 U2434 ( .A(n9868), .Y(n1467) );
  BUFX2 U2435 ( .A(n9887), .Y(n1468) );
  BUFX2 U2436 ( .A(n9906), .Y(n1469) );
  BUFX2 U2437 ( .A(n9923), .Y(n1470) );
  BUFX2 U2438 ( .A(n10018), .Y(n1471) );
  BUFX2 U2439 ( .A(n10031), .Y(n1472) );
  BUFX2 U2440 ( .A(n10040), .Y(n1473) );
  BUFX2 U2441 ( .A(n10050), .Y(n1474) );
  BUFX2 U2442 ( .A(n10083), .Y(n1475) );
  BUFX2 U2443 ( .A(n10090), .Y(n1476) );
  BUFX2 U2444 ( .A(n10099), .Y(n1477) );
  BUFX2 U2445 ( .A(n10170), .Y(n1478) );
  BUFX2 U2446 ( .A(n10180), .Y(n1479) );
  BUFX2 U2447 ( .A(n10206), .Y(n1480) );
  BUFX2 U2448 ( .A(n10235), .Y(n1481) );
  BUFX2 U2449 ( .A(n10285), .Y(n1482) );
  BUFX2 U2450 ( .A(n10298), .Y(n1483) );
  BUFX2 U2451 ( .A(n10324), .Y(n1484) );
  BUFX2 U2452 ( .A(n10389), .Y(n1485) );
  BUFX2 U2453 ( .A(n10394), .Y(n1486) );
  BUFX2 U2454 ( .A(n10587), .Y(n1487) );
  BUFX2 U2455 ( .A(n6743), .Y(n1488) );
  BUFX2 U2456 ( .A(n7431), .Y(n1489) );
  INVX1 U2457 ( .A(n7765), .Y(n1490) );
  INVX1 U2458 ( .A(n1490), .Y(n1491) );
  BUFX2 U2459 ( .A(n8772), .Y(n1492) );
  BUFX2 U2460 ( .A(n9276), .Y(n1493) );
  INVX1 U2461 ( .A(n9806), .Y(n1494) );
  INVX1 U2462 ( .A(n1494), .Y(n1495) );
  AND2X2 U2463 ( .A(n6275), .B(n5730), .Y(n6436) );
  INVX1 U2464 ( .A(n6436), .Y(n1496) );
  AND2X1 U2465 ( .A(n66), .B(n5730), .Y(n6438) );
  INVX1 U2466 ( .A(n6438), .Y(n1497) );
  AND2X1 U2467 ( .A(n520), .B(n6143), .Y(n6473) );
  INVX1 U2468 ( .A(n6473), .Y(n1498) );
  AND2X1 U2469 ( .A(n2198), .B(n5782), .Y(n6536) );
  INVX1 U2470 ( .A(n6536), .Y(n1499) );
  AND2X1 U2471 ( .A(n522), .B(n5773), .Y(n6619) );
  INVX1 U2472 ( .A(n6619), .Y(n1500) );
  AND2X1 U2473 ( .A(n2200), .B(n6113), .Y(n6690) );
  INVX1 U2474 ( .A(n6690), .Y(n1501) );
  AND2X1 U2475 ( .A(n523), .B(n6143), .Y(n6697) );
  INVX1 U2476 ( .A(n6697), .Y(n1502) );
  AND2X1 U2477 ( .A(n2201), .B(n6113), .Y(n6758) );
  INVX1 U2478 ( .A(n6758), .Y(n1503) );
  AND2X1 U2479 ( .A(n524), .B(n5773), .Y(n6765) );
  INVX1 U2480 ( .A(n6765), .Y(n1504) );
  AND2X1 U2481 ( .A(n2202), .B(n6113), .Y(n6814) );
  INVX1 U2482 ( .A(n6814), .Y(n1505) );
  AND2X1 U2483 ( .A(n525), .B(n5773), .Y(n6821) );
  INVX1 U2484 ( .A(n6821), .Y(n1506) );
  AND2X1 U2485 ( .A(n2203), .B(n6113), .Y(n6877) );
  INVX1 U2486 ( .A(n6877), .Y(n1507) );
  AND2X1 U2487 ( .A(n2236), .B(n5838), .Y(n6889) );
  INVX1 U2488 ( .A(n6889), .Y(n1508) );
  AND2X1 U2489 ( .A(n2525), .B(n5856), .Y(n6902) );
  INVX1 U2490 ( .A(n6902), .Y(n1509) );
  OR2X1 U2491 ( .A(n6929), .B(n6928), .Y(n6930) );
  INVX1 U2492 ( .A(n6930), .Y(n1510) );
  AND2X1 U2493 ( .A(n2205), .B(n6113), .Y(n6997) );
  INVX1 U2494 ( .A(n6997), .Y(n1511) );
  AND2X1 U2495 ( .A(n528), .B(n5773), .Y(n7004) );
  INVX1 U2496 ( .A(n7004), .Y(n1512) );
  AND2X1 U2497 ( .A(n2206), .B(n6113), .Y(n7054) );
  INVX1 U2498 ( .A(n7054), .Y(n1513) );
  AND2X1 U2499 ( .A(n529), .B(n5773), .Y(n7061) );
  INVX1 U2500 ( .A(n7061), .Y(n1514) );
  AND2X1 U2501 ( .A(n2207), .B(n5782), .Y(n7124) );
  INVX1 U2502 ( .A(n7124), .Y(n1515) );
  AND2X1 U2503 ( .A(n2208), .B(n6113), .Y(n7199) );
  INVX1 U2504 ( .A(n7199), .Y(n1517) );
  AND2X1 U2505 ( .A(n2209), .B(n5782), .Y(n7265) );
  INVX1 U2506 ( .A(n7265), .Y(n1533) );
  AND2X1 U2507 ( .A(n532), .B(n5773), .Y(n7272) );
  INVX1 U2508 ( .A(n7272), .Y(n1549) );
  AND2X1 U2509 ( .A(n2210), .B(n6113), .Y(n7327) );
  INVX1 U2510 ( .A(n7327), .Y(n1565) );
  AND2X1 U2511 ( .A(n533), .B(n5773), .Y(n7334) );
  INVX1 U2512 ( .A(n7334), .Y(n1581) );
  AND2X1 U2513 ( .A(n2211), .B(n5782), .Y(n7392) );
  INVX1 U2514 ( .A(n7392), .Y(n1613) );
  AND2X1 U2515 ( .A(n534), .B(n5773), .Y(n7399) );
  INVX1 U2516 ( .A(n7399), .Y(n1644) );
  AND2X1 U2517 ( .A(n2212), .B(n5782), .Y(n7458) );
  INVX1 U2518 ( .A(n7458), .Y(n1645) );
  AND2X1 U2519 ( .A(n535), .B(n6143), .Y(n7465) );
  INVX1 U2520 ( .A(n7465), .Y(n1646) );
  AND2X1 U2521 ( .A(n2213), .B(n5782), .Y(n7510) );
  INVX1 U2522 ( .A(n7510), .Y(n1647) );
  AND2X1 U2523 ( .A(n536), .B(n6143), .Y(n7517) );
  INVX1 U2524 ( .A(n7517), .Y(n1648) );
  AND2X1 U2525 ( .A(n2214), .B(n5782), .Y(n7569) );
  INVX1 U2526 ( .A(n7569), .Y(n1649) );
  AND2X1 U2527 ( .A(n537), .B(n6143), .Y(n7576) );
  INVX1 U2528 ( .A(n7576), .Y(n1650) );
  AND2X1 U2529 ( .A(n2215), .B(n5782), .Y(n7643) );
  INVX1 U2530 ( .A(n7643), .Y(n1651) );
  AND2X1 U2531 ( .A(n538), .B(n6143), .Y(n7650) );
  INVX1 U2532 ( .A(n7650), .Y(n1652) );
  AND2X1 U2533 ( .A(n2216), .B(n5782), .Y(n7718) );
  INVX1 U2534 ( .A(n7718), .Y(n1653) );
  AND2X1 U2535 ( .A(n539), .B(n6143), .Y(n7725) );
  INVX1 U2536 ( .A(n7725), .Y(n1654) );
  AND2X1 U2537 ( .A(n2217), .B(n5782), .Y(n7780) );
  INVX1 U2538 ( .A(n7780), .Y(n1655) );
  AND2X1 U2539 ( .A(n540), .B(n6143), .Y(n7787) );
  INVX1 U2540 ( .A(n7787), .Y(n1656) );
  AND2X1 U2541 ( .A(n2218), .B(n5782), .Y(n7831) );
  INVX1 U2542 ( .A(n7831), .Y(n1657) );
  AND2X1 U2543 ( .A(n541), .B(n6143), .Y(n7838) );
  INVX1 U2544 ( .A(n7838), .Y(n1658) );
  AND2X1 U2545 ( .A(n2219), .B(n5782), .Y(n7896) );
  INVX1 U2546 ( .A(n7896), .Y(n1659) );
  AND2X1 U2547 ( .A(n542), .B(n6143), .Y(n7903) );
  INVX1 U2548 ( .A(n7903), .Y(n1660) );
  AND2X1 U2549 ( .A(n1120), .B(n5826), .Y(n7921) );
  INVX1 U2550 ( .A(n7921), .Y(n1661) );
  AND2X1 U2551 ( .A(n2220), .B(n5782), .Y(n7959) );
  INVX1 U2552 ( .A(n7959), .Y(n1662) );
  AND2X1 U2553 ( .A(n543), .B(n6143), .Y(n7966) );
  INVX1 U2554 ( .A(n7966), .Y(n1663) );
  AND2X1 U2555 ( .A(n2221), .B(n5782), .Y(n8010) );
  INVX1 U2556 ( .A(n8010), .Y(n1664) );
  AND2X1 U2557 ( .A(n544), .B(n6143), .Y(n8017) );
  INVX1 U2558 ( .A(n8017), .Y(n1665) );
  AND2X1 U2559 ( .A(n2222), .B(n5782), .Y(n8067) );
  INVX1 U2560 ( .A(n8067), .Y(n1666) );
  AND2X1 U2561 ( .A(n545), .B(n6143), .Y(n8074) );
  INVX1 U2562 ( .A(n8074), .Y(n1667) );
  AND2X1 U2563 ( .A(n2223), .B(n5782), .Y(n8142) );
  INVX1 U2564 ( .A(n8142), .Y(n1668) );
  AND2X1 U2565 ( .A(n546), .B(n6143), .Y(n8149) );
  INVX1 U2566 ( .A(n8149), .Y(n1669) );
  AND2X1 U2567 ( .A(n2224), .B(n5782), .Y(n8216) );
  INVX1 U2568 ( .A(n8216), .Y(n1670) );
  AND2X1 U2569 ( .A(n547), .B(n6143), .Y(n8223) );
  INVX1 U2570 ( .A(n8223), .Y(n1671) );
  AND2X1 U2571 ( .A(n2225), .B(n5782), .Y(n8280) );
  INVX1 U2572 ( .A(n8280), .Y(n1672) );
  AND2X1 U2573 ( .A(n548), .B(n6143), .Y(n8287) );
  INVX1 U2574 ( .A(n8287), .Y(n1673) );
  AND2X1 U2575 ( .A(n2226), .B(n5782), .Y(n8343) );
  INVX1 U2576 ( .A(n8343), .Y(n1674) );
  AND2X1 U2577 ( .A(n2227), .B(n5782), .Y(n8406) );
  INVX1 U2578 ( .A(n8406), .Y(n1675) );
  AND2X1 U2579 ( .A(n470), .B(n5839), .Y(n8457) );
  INVX1 U2580 ( .A(n8457), .Y(n1676) );
  AND2X1 U2581 ( .A(n2582), .B(n5831), .Y(n8504) );
  INVX1 U2582 ( .A(n8504), .Y(n1677) );
  AND2X1 U2583 ( .A(n488), .B(n6143), .Y(n8521) );
  INVX1 U2584 ( .A(n8521), .Y(n1678) );
  AND2X1 U2585 ( .A(n2166), .B(n5782), .Y(n8573) );
  INVX1 U2586 ( .A(n8573), .Y(n1679) );
  AND2X1 U2587 ( .A(n2489), .B(n5856), .Y(n8670) );
  INVX1 U2588 ( .A(n8670), .Y(n1680) );
  OR2X1 U2589 ( .A(n8707), .B(n8706), .Y(n8708) );
  INVX1 U2590 ( .A(n8708), .Y(n1681) );
  AND2X1 U2591 ( .A(n491), .B(n6143), .Y(n8731) );
  INVX1 U2592 ( .A(n8731), .Y(n1682) );
  AND2X1 U2593 ( .A(n2169), .B(n5782), .Y(n8787) );
  INVX1 U2594 ( .A(n8787), .Y(n1683) );
  AND2X1 U2595 ( .A(n492), .B(n5773), .Y(n8794) );
  INVX1 U2596 ( .A(n8794), .Y(n1684) );
  AND2X1 U2597 ( .A(n2170), .B(n5782), .Y(n8839) );
  INVX1 U2598 ( .A(n8839), .Y(n1685) );
  AND2X1 U2599 ( .A(n493), .B(n6143), .Y(n8846) );
  INVX1 U2600 ( .A(n8846), .Y(n1686) );
  AND2X1 U2601 ( .A(n2171), .B(n5782), .Y(n8902) );
  INVX1 U2602 ( .A(n8902), .Y(n1687) );
  AND2X1 U2603 ( .A(n2268), .B(n5838), .Y(n8915) );
  INVX1 U2604 ( .A(n8915), .Y(n1688) );
  AND2X1 U2605 ( .A(n2493), .B(n5856), .Y(n8928) );
  INVX1 U2606 ( .A(n8928), .Y(n1689) );
  OR2X1 U2607 ( .A(n8956), .B(n8955), .Y(n8957) );
  INVX1 U2608 ( .A(n8957), .Y(n1690) );
  AND2X1 U2609 ( .A(n495), .B(n5773), .Y(n8979) );
  INVX1 U2610 ( .A(n8979), .Y(n1691) );
  AND2X1 U2611 ( .A(n2173), .B(n5782), .Y(n9021) );
  INVX1 U2612 ( .A(n9021), .Y(n1692) );
  AND2X1 U2613 ( .A(n496), .B(n5773), .Y(n9028) );
  INVX1 U2614 ( .A(n9028), .Y(n1693) );
  AND2X1 U2615 ( .A(n2174), .B(n5782), .Y(n9079) );
  INVX1 U2616 ( .A(n9079), .Y(n1694) );
  AND2X1 U2617 ( .A(n497), .B(n6143), .Y(n9086) );
  INVX1 U2618 ( .A(n9086), .Y(n1695) );
  AND2X1 U2619 ( .A(n2175), .B(n5782), .Y(n9154) );
  INVX1 U2620 ( .A(n9154), .Y(n1696) );
  AND2X1 U2621 ( .A(n498), .B(n5773), .Y(n9161) );
  INVX1 U2622 ( .A(n9161), .Y(n1697) );
  AND2X1 U2623 ( .A(n2176), .B(n5782), .Y(n9228) );
  INVX1 U2624 ( .A(n9228), .Y(n1698) );
  AND2X1 U2625 ( .A(n499), .B(n6143), .Y(n9235) );
  INVX1 U2626 ( .A(n9235), .Y(n1699) );
  AND2X1 U2627 ( .A(n2177), .B(n5782), .Y(n9290) );
  INVX1 U2628 ( .A(n9290), .Y(n1700) );
  AND2X1 U2629 ( .A(n500), .B(n6143), .Y(n9297) );
  INVX1 U2630 ( .A(n9297), .Y(n1701) );
  AND2X1 U2631 ( .A(n2178), .B(n5782), .Y(n9353) );
  INVX1 U2632 ( .A(n9353), .Y(n1702) );
  AND2X1 U2633 ( .A(n501), .B(n5773), .Y(n9360) );
  INVX1 U2634 ( .A(n9360), .Y(n1703) );
  AND2X1 U2635 ( .A(n2179), .B(n5782), .Y(n9417) );
  INVX1 U2636 ( .A(n9417), .Y(n1704) );
  AND2X1 U2637 ( .A(n502), .B(n5773), .Y(n9436) );
  INVX1 U2638 ( .A(n9436), .Y(n1705) );
  AND2X1 U2639 ( .A(n2180), .B(n6113), .Y(n9448) );
  INVX1 U2640 ( .A(n9448), .Y(n1706) );
  OR2X1 U2641 ( .A(n9465), .B(n2341), .Y(n9466) );
  INVX1 U2642 ( .A(n9466), .Y(n1707) );
  AND2X1 U2643 ( .A(n1546), .B(n6123), .Y(n9468) );
  INVX1 U2644 ( .A(n9468), .Y(n1708) );
  AND2X1 U2645 ( .A(n503), .B(n6143), .Y(n9487) );
  INVX1 U2646 ( .A(n9487), .Y(n1709) );
  AND2X1 U2647 ( .A(n2181), .B(n5782), .Y(n9537) );
  INVX1 U2648 ( .A(n9537), .Y(n1710) );
  AND2X1 U2649 ( .A(n504), .B(n5773), .Y(n9544) );
  INVX1 U2650 ( .A(n9544), .Y(n1711) );
  AND2X1 U2651 ( .A(n2182), .B(n5782), .Y(n9597) );
  INVX1 U2652 ( .A(n9597), .Y(n1712) );
  AND2X1 U2653 ( .A(n505), .B(n6143), .Y(n9604) );
  INVX1 U2654 ( .A(n9604), .Y(n1713) );
  AND2X1 U2655 ( .A(n2183), .B(n5782), .Y(n9675) );
  INVX1 U2656 ( .A(n9675), .Y(n1714) );
  AND2X1 U2657 ( .A(n506), .B(n5773), .Y(n9682) );
  INVX1 U2658 ( .A(n9682), .Y(n1715) );
  AND2X1 U2659 ( .A(n2184), .B(n5782), .Y(n9753) );
  INVX1 U2660 ( .A(n9753), .Y(n1716) );
  AND2X1 U2661 ( .A(n507), .B(n6143), .Y(n9760) );
  INVX1 U2662 ( .A(n9760), .Y(n1717) );
  AND2X1 U2663 ( .A(n2185), .B(n5782), .Y(n9821) );
  INVX1 U2664 ( .A(n9821), .Y(n1718) );
  AND2X1 U2665 ( .A(n508), .B(n5773), .Y(n9828) );
  INVX1 U2666 ( .A(n9828), .Y(n1719) );
  AND2X1 U2667 ( .A(n2186), .B(n5782), .Y(n9875) );
  INVX1 U2668 ( .A(n9875), .Y(n1720) );
  AND2X1 U2669 ( .A(n509), .B(n5773), .Y(n9882) );
  INVX1 U2670 ( .A(n9882), .Y(n1721) );
  AND2X1 U2671 ( .A(n2187), .B(n5782), .Y(n9941) );
  INVX1 U2672 ( .A(n9941), .Y(n1722) );
  AND2X1 U2673 ( .A(n510), .B(n6143), .Y(n9948) );
  INVX1 U2674 ( .A(n9948), .Y(n1723) );
  AND2X1 U2675 ( .A(n1088), .B(n6127), .Y(n9966) );
  INVX1 U2676 ( .A(n9966), .Y(n1724) );
  AND2X1 U2677 ( .A(n2188), .B(n5782), .Y(n10005) );
  INVX1 U2678 ( .A(n10005), .Y(n1725) );
  AND2X1 U2679 ( .A(n511), .B(n5773), .Y(n10012) );
  INVX1 U2680 ( .A(n10012), .Y(n1726) );
  AND2X1 U2681 ( .A(n2189), .B(n5782), .Y(n10056) );
  INVX1 U2682 ( .A(n10056), .Y(n1727) );
  AND2X1 U2683 ( .A(n512), .B(n6143), .Y(n10063) );
  INVX1 U2684 ( .A(n10063), .Y(n1728) );
  AND2X1 U2685 ( .A(n2190), .B(n5782), .Y(n10119) );
  INVX1 U2686 ( .A(n10119), .Y(n1729) );
  AND2X1 U2687 ( .A(n513), .B(n5773), .Y(n10126) );
  INVX1 U2688 ( .A(n10126), .Y(n1730) );
  AND2X1 U2689 ( .A(n2191), .B(n5782), .Y(n10194) );
  INVX1 U2690 ( .A(n10194), .Y(n1731) );
  AND2X1 U2691 ( .A(n514), .B(n6143), .Y(n10201) );
  INVX1 U2692 ( .A(n10201), .Y(n1732) );
  AND2X1 U2693 ( .A(n2192), .B(n5782), .Y(n10268) );
  INVX1 U2694 ( .A(n10268), .Y(n1733) );
  AND2X1 U2695 ( .A(n515), .B(n5773), .Y(n10275) );
  INVX1 U2696 ( .A(n10275), .Y(n1734) );
  AND2X1 U2697 ( .A(n2193), .B(n5782), .Y(n10335) );
  INVX1 U2698 ( .A(n10335), .Y(n1735) );
  AND2X1 U2699 ( .A(n516), .B(n6143), .Y(n10342) );
  INVX1 U2700 ( .A(n10342), .Y(n1736) );
  AND2X1 U2701 ( .A(n2194), .B(n5782), .Y(n10405) );
  INVX1 U2702 ( .A(n10405), .Y(n1737) );
  AND2X1 U2703 ( .A(n2195), .B(n6113), .Y(n10472) );
  INVX1 U2704 ( .A(n10472), .Y(n1738) );
  AND2X1 U2705 ( .A(n3160), .B(n5776), .Y(n10585) );
  INVX1 U2706 ( .A(n10585), .Y(n1739) );
  BUFX2 U2707 ( .A(n6484), .Y(n1740) );
  BUFX2 U2708 ( .A(n6624), .Y(n1742) );
  BUFX2 U2709 ( .A(n6711), .Y(n1758) );
  BUFX2 U2710 ( .A(n6912), .Y(n1774) );
  BUFX2 U2711 ( .A(n6919), .Y(n1790) );
  BUFX2 U2712 ( .A(n6927), .Y(n1806) );
  BUFX2 U2713 ( .A(n7074), .Y(n1838) );
  BUFX2 U2714 ( .A(n7406), .Y(n1869) );
  BUFX2 U2715 ( .A(n7423), .Y(n1870) );
  BUFX2 U2716 ( .A(n7477), .Y(n1871) );
  BUFX2 U2717 ( .A(n7528), .Y(n1872) );
  BUFX2 U2718 ( .A(n7655), .Y(n1873) );
  BUFX2 U2719 ( .A(n7738), .Y(n1874) );
  BUFX2 U2720 ( .A(n8484), .Y(n1875) );
  BUFX2 U2721 ( .A(n8532), .Y(n1876) );
  BUFX2 U2722 ( .A(n8680), .Y(n1877) );
  BUFX2 U2723 ( .A(n8682), .Y(n1878) );
  BUFX2 U2724 ( .A(n8699), .Y(n1879) );
  BUFX2 U2725 ( .A(n8705), .Y(n1880) );
  BUFX2 U2726 ( .A(n8745), .Y(n1881) );
  BUFX2 U2727 ( .A(n8938), .Y(n1882) );
  BUFX2 U2728 ( .A(n8945), .Y(n1883) );
  BUFX2 U2729 ( .A(n8953), .Y(n1884) );
  BUFX2 U2730 ( .A(n9451), .Y(n1885) );
  BUFX2 U2731 ( .A(n9459), .Y(n1886) );
  BUFX2 U2732 ( .A(n9499), .Y(n1887) );
  BUFX2 U2733 ( .A(n9555), .Y(n1888) );
  BUFX2 U2734 ( .A(n9687), .Y(n1889) );
  BUFX2 U2735 ( .A(n9773), .Y(n1890) );
  BUFX2 U2736 ( .A(n10496), .Y(n1891) );
  BUFX2 U2737 ( .A(n10501), .Y(n1892) );
  BUFX2 U2738 ( .A(n10562), .Y(n1893) );
  BUFX2 U2739 ( .A(n6642), .Y(n1894) );
  BUFX2 U2740 ( .A(n6651), .Y(n1895) );
  BUFX2 U2741 ( .A(n6914), .Y(n1896) );
  BUFX2 U2742 ( .A(n7072), .Y(n1897) );
  BUFX2 U2743 ( .A(n7082), .Y(n1898) );
  BUFX2 U2744 ( .A(n7088), .Y(n1899) );
  BUFX2 U2745 ( .A(n7426), .Y(n1900) );
  BUFX2 U2746 ( .A(n7670), .Y(n1901) );
  BUFX2 U2747 ( .A(n7679), .Y(n1902) );
  BUFX2 U2748 ( .A(n8098), .Y(n1903) );
  BUFX2 U2749 ( .A(n8099), .Y(n1904) );
  BUFX2 U2750 ( .A(n8132), .Y(n1905) );
  BUFX2 U2751 ( .A(n8719), .Y(n1906) );
  BUFX2 U2752 ( .A(n8940), .Y(n1907) );
  BUFX2 U2753 ( .A(n9110), .Y(n1908) );
  BUFX2 U2754 ( .A(n9111), .Y(n1909) );
  BUFX2 U2755 ( .A(n9144), .Y(n1910) );
  BUFX2 U2756 ( .A(n9453), .Y(n1911) );
  BUFX2 U2757 ( .A(n9702), .Y(n1912) );
  BUFX2 U2758 ( .A(n9712), .Y(n1913) );
  BUFX2 U2759 ( .A(n10150), .Y(n1914) );
  BUFX2 U2760 ( .A(n10151), .Y(n1915) );
  BUFX2 U2761 ( .A(n10184), .Y(n1916) );
  AND2X1 U2762 ( .A(n6076), .B(n6024), .Y(n6450) );
  INVX1 U2763 ( .A(n6450), .Y(n1917) );
  AND2X1 U2764 ( .A(n6790), .B(n6080), .Y(n6507) );
  INVX1 U2765 ( .A(n6507), .Y(n1918) );
  AND2X1 U2766 ( .A(n6790), .B(n6081), .Y(n6508) );
  INVX1 U2767 ( .A(n6508), .Y(n1919) );
  AND2X1 U2768 ( .A(n6790), .B(n6077), .Y(n6509) );
  INVX1 U2769 ( .A(n6509), .Y(n1920) );
  AND2X1 U2770 ( .A(n7490), .B(n7362), .Y(n6566) );
  INVX1 U2771 ( .A(n6566), .Y(n1921) );
  AND2X1 U2772 ( .A(n1958), .B(n6142), .Y(n6612) );
  INVX1 U2773 ( .A(n6612), .Y(n1922) );
  AND2X1 U2774 ( .A(n10487), .B(n6659), .Y(n6660) );
  INVX1 U2775 ( .A(n6660), .Y(n1923) );
  AND2X1 U2776 ( .A(n847), .B(n5857), .Y(n6884) );
  INVX1 U2777 ( .A(n6884), .Y(n1924) );
  AND2X1 U2778 ( .A(n6791), .B(n6939), .Y(n6940) );
  INVX1 U2779 ( .A(n6940), .Y(n1925) );
  AND2X1 U2780 ( .A(n5515), .B(n10505), .Y(n7149) );
  INVX1 U2781 ( .A(n7149), .Y(n1926) );
  AND2X1 U2782 ( .A(n7490), .B(n8378), .Y(n7599) );
  INVX1 U2783 ( .A(n7599), .Y(n1927) );
  AND2X1 U2784 ( .A(n10487), .B(n7688), .Y(n7689) );
  INVX1 U2785 ( .A(n7689), .Y(n1928) );
  AND2X1 U2786 ( .A(n8172), .B(n10491), .Y(n8173) );
  INVX1 U2787 ( .A(n8173), .Y(n1929) );
  AND2X1 U2788 ( .A(n7490), .B(n9388), .Y(n8601) );
  INVX1 U2789 ( .A(n8601), .Y(n1930) );
  AND2X1 U2790 ( .A(n1960), .B(n6142), .Y(n8645) );
  INVX1 U2791 ( .A(n8645), .Y(n1931) );
  AND2X1 U2792 ( .A(n10487), .B(n8693), .Y(n8694) );
  INVX1 U2793 ( .A(n8694), .Y(n1932) );
  AND2X1 U2794 ( .A(n3548), .B(n6092), .Y(n8720) );
  INVX1 U2795 ( .A(n8720), .Y(n1933) );
  AND2X1 U2796 ( .A(n815), .B(n5857), .Y(n8909) );
  INVX1 U2797 ( .A(n8909), .Y(n1934) );
  AND2X1 U2798 ( .A(n6791), .B(n8966), .Y(n8967) );
  INVX1 U2799 ( .A(n8967), .Y(n1935) );
  AND2X1 U2800 ( .A(n9046), .B(n4852), .Y(n9476) );
  INVX1 U2801 ( .A(n9476), .Y(n1936) );
  AND2X1 U2802 ( .A(n9460), .B(n5053), .Y(n9497) );
  INVX1 U2803 ( .A(n9497), .Y(n1937) );
  AND2X1 U2804 ( .A(n7490), .B(n10440), .Y(n9628) );
  INVX1 U2805 ( .A(n9628), .Y(n1938) );
  AND2X1 U2806 ( .A(n10487), .B(n9722), .Y(n9723) );
  INVX1 U2807 ( .A(n9723), .Y(n1939) );
  AND2X1 U2808 ( .A(n10222), .B(n10491), .Y(n10223) );
  INVX1 U2809 ( .A(n10223), .Y(n1940) );
  AND2X1 U2810 ( .A(n6054), .B(n5220), .Y(n10563) );
  INVX1 U2811 ( .A(n10563), .Y(n1941) );
  BUFX2 U2812 ( .A(n6365), .Y(n1942) );
  BUFX2 U2813 ( .A(n6427), .Y(n1943) );
  BUFX2 U2814 ( .A(n7486), .Y(n1944) );
  AND2X1 U2815 ( .A(n1770), .B(n5777), .Y(n9409) );
  INVX1 U2816 ( .A(n9409), .Y(n1945) );
  AND2X1 U2817 ( .A(n454), .B(n5839), .Y(n9427) );
  INVX1 U2818 ( .A(n9427), .Y(n1946) );
  AND2X1 U2819 ( .A(n1270), .B(n5785), .Y(n10327) );
  INVX1 U2820 ( .A(n10327), .Y(n1947) );
  AND2X1 U2821 ( .A(n1754), .B(n5777), .Y(n10463) );
  INVX1 U2822 ( .A(n10463), .Y(n1948) );
  BUFX2 U2823 ( .A(n6366), .Y(n1949) );
  INVX1 U2824 ( .A(n6428), .Y(n1950) );
  INVX1 U2825 ( .A(n1950), .Y(n1951) );
  BUFX2 U2826 ( .A(n9410), .Y(n1952) );
  BUFX2 U2827 ( .A(n10328), .Y(n1953) );
  INVX1 U2828 ( .A(n10326), .Y(n1954) );
  INVX1 U2829 ( .A(n1954), .Y(n1955) );
  BUFX2 U2830 ( .A(n10464), .Y(n1956) );
  BUFX2 U2831 ( .A(n10462), .Y(n1957) );
  BUFX2 U2832 ( .A(n6611), .Y(n1958) );
  BUFX2 U2833 ( .A(n7485), .Y(n1959) );
  BUFX2 U2834 ( .A(n8644), .Y(n1960) );
  BUFX2 U2835 ( .A(n9426), .Y(n1961) );
  BUFX2 U2836 ( .A(n6575), .Y(n1962) );
  BUFX2 U2837 ( .A(n7607), .Y(n1963) );
  BUFX2 U2838 ( .A(n8612), .Y(n1964) );
  BUFX2 U2839 ( .A(n9641), .Y(n1965) );
  BUFX2 U2840 ( .A(n6542), .Y(n1966) );
  BUFX2 U2841 ( .A(n6618), .Y(n1967) );
  BUFX2 U2842 ( .A(n6600), .Y(n1968) );
  BUFX2 U2843 ( .A(n6696), .Y(n1969) );
  BUFX2 U2844 ( .A(n6648), .Y(n1970) );
  BUFX2 U2845 ( .A(n6667), .Y(n1971) );
  BUFX2 U2846 ( .A(n6677), .Y(n1972) );
  BUFX2 U2847 ( .A(n6764), .Y(n1973) );
  BUFX2 U2848 ( .A(n6820), .Y(n1974) );
  BUFX2 U2849 ( .A(n6883), .Y(n1975) );
  BUFX2 U2850 ( .A(n6842), .Y(n1976) );
  BUFX2 U2851 ( .A(n7003), .Y(n1977) );
  BUFX2 U2852 ( .A(n7060), .Y(n1978) );
  BUFX2 U2853 ( .A(n7130), .Y(n1979) );
  BUFX2 U2854 ( .A(n7101), .Y(n1980) );
  BUFX2 U2855 ( .A(n7112), .Y(n1981) );
  BUFX2 U2856 ( .A(n7205), .Y(n1982) );
  BUFX2 U2857 ( .A(n7177), .Y(n1983) );
  BUFX2 U2858 ( .A(n7187), .Y(n1984) );
  BUFX2 U2859 ( .A(n7271), .Y(n1985) );
  BUFX2 U2860 ( .A(n7333), .Y(n1986) );
  BUFX2 U2861 ( .A(n7295), .Y(n1987) );
  BUFX2 U2862 ( .A(n7398), .Y(n1988) );
  BUFX2 U2863 ( .A(n7350), .Y(n1989) );
  BUFX2 U2864 ( .A(n7368), .Y(n1990) );
  BUFX2 U2865 ( .A(n7380), .Y(n1991) );
  BUFX2 U2866 ( .A(n7464), .Y(n1992) );
  BUFX2 U2867 ( .A(n7516), .Y(n1993) );
  BUFX2 U2868 ( .A(n7575), .Y(n1994) );
  BUFX2 U2869 ( .A(n7649), .Y(n1995) );
  BUFX2 U2870 ( .A(n7631), .Y(n1996) );
  BUFX2 U2871 ( .A(n7724), .Y(n1997) );
  BUFX2 U2872 ( .A(n7676), .Y(n1998) );
  BUFX2 U2873 ( .A(n7696), .Y(n1999) );
  BUFX2 U2874 ( .A(n7706), .Y(n2000) );
  BUFX2 U2875 ( .A(n7786), .Y(n2001) );
  BUFX2 U2876 ( .A(n7837), .Y(n2002) );
  BUFX2 U2877 ( .A(n7902), .Y(n2003) );
  BUFX2 U2878 ( .A(n7859), .Y(n2004) );
  BUFX2 U2879 ( .A(n7965), .Y(n2005) );
  BUFX2 U2880 ( .A(n7915), .Y(n2006) );
  BUFX2 U2881 ( .A(n7938), .Y(n2007) );
  BUFX2 U2882 ( .A(n8016), .Y(n2008) );
  BUFX2 U2883 ( .A(n8073), .Y(n2009) );
  BUFX2 U2884 ( .A(n8148), .Y(n2010) );
  BUFX2 U2885 ( .A(n8086), .Y(n2011) );
  BUFX2 U2886 ( .A(n8096), .Y(n2012) );
  BUFX2 U2887 ( .A(n8222), .Y(n2013) );
  BUFX2 U2888 ( .A(n8286), .Y(n2014) );
  BUFX2 U2889 ( .A(n8349), .Y(n2015) );
  BUFX2 U2890 ( .A(n8367), .Y(n2016) );
  BUFX2 U2891 ( .A(n8384), .Y(n2017) );
  BUFX2 U2892 ( .A(n8444), .Y(n2018) );
  BUFX2 U2893 ( .A(n8579), .Y(n2019) );
  BUFX2 U2894 ( .A(n8651), .Y(n2020) );
  BUFX2 U2895 ( .A(n8633), .Y(n2021) );
  BUFX2 U2896 ( .A(n8793), .Y(n2022) );
  BUFX2 U2897 ( .A(n8845), .Y(n2023) );
  BUFX2 U2898 ( .A(n8908), .Y(n2024) );
  BUFX2 U2899 ( .A(n8867), .Y(n2025) );
  BUFX2 U2900 ( .A(n9027), .Y(n2026) );
  BUFX2 U2901 ( .A(n9085), .Y(n2027) );
  BUFX2 U2902 ( .A(n9160), .Y(n2028) );
  BUFX2 U2903 ( .A(n9098), .Y(n2029) );
  BUFX2 U2904 ( .A(n9108), .Y(n2030) );
  BUFX2 U2905 ( .A(n9234), .Y(n2031) );
  BUFX2 U2906 ( .A(n9215), .Y(n2032) );
  BUFX2 U2907 ( .A(n9296), .Y(n2033) );
  BUFX2 U2908 ( .A(n9359), .Y(n2034) );
  BUFX2 U2909 ( .A(n9321), .Y(n2035) );
  BUFX2 U2910 ( .A(n9423), .Y(n2036) );
  BUFX2 U2911 ( .A(n9377), .Y(n2037) );
  BUFX2 U2912 ( .A(n9394), .Y(n2038) );
  BUFX2 U2913 ( .A(n9404), .Y(n2039) );
  BUFX2 U2914 ( .A(n9543), .Y(n2040) );
  BUFX2 U2915 ( .A(n9603), .Y(n2041) );
  BUFX2 U2916 ( .A(n9681), .Y(n2042) );
  BUFX2 U2917 ( .A(n9663), .Y(n2043) );
  BUFX2 U2918 ( .A(n9759), .Y(n2044) );
  BUFX2 U2919 ( .A(n9709), .Y(n2045) );
  BUFX2 U2920 ( .A(n9730), .Y(n2046) );
  BUFX2 U2921 ( .A(n9741), .Y(n2047) );
  BUFX2 U2922 ( .A(n9827), .Y(n2048) );
  BUFX2 U2923 ( .A(n9881), .Y(n2049) );
  BUFX2 U2924 ( .A(n9947), .Y(n2050) );
  BUFX2 U2925 ( .A(n9903), .Y(n2051) );
  BUFX2 U2926 ( .A(n10011), .Y(n2052) );
  BUFX2 U2927 ( .A(n9960), .Y(n2053) );
  BUFX2 U2928 ( .A(n9984), .Y(n2054) );
  BUFX2 U2929 ( .A(n10062), .Y(n2055) );
  BUFX2 U2930 ( .A(n10125), .Y(n2056) );
  BUFX2 U2931 ( .A(n10200), .Y(n2057) );
  BUFX2 U2932 ( .A(n10138), .Y(n2058) );
  BUFX2 U2933 ( .A(n10148), .Y(n2059) );
  BUFX2 U2934 ( .A(n10274), .Y(n2060) );
  BUFX2 U2935 ( .A(n10255), .Y(n2061) );
  BUFX2 U2936 ( .A(n10341), .Y(n2062) );
  BUFX2 U2937 ( .A(n10411), .Y(n2063) );
  BUFX2 U2938 ( .A(n10366), .Y(n2064) );
  BUFX2 U2939 ( .A(n10429), .Y(n2065) );
  BUFX2 U2940 ( .A(n10446), .Y(n2066) );
  INVX1 U2941 ( .A(n6563), .Y(n2067) );
  INVX1 U2942 ( .A(n6589), .Y(n2068) );
  INVX1 U2943 ( .A(n6832), .Y(n2069) );
  INVX1 U2944 ( .A(n7283), .Y(n2070) );
  INVX1 U2945 ( .A(n7596), .Y(n2071) );
  INVX1 U2946 ( .A(n7621), .Y(n2072) );
  INVX1 U2947 ( .A(n7849), .Y(n2073) );
  INVX1 U2948 ( .A(n8194), .Y(n2074) );
  INVX1 U2949 ( .A(n8298), .Y(n2075) );
  INVX1 U2950 ( .A(n8424), .Y(n2076) );
  INVX1 U2951 ( .A(n8598), .Y(n2077) );
  INVX1 U2952 ( .A(n8623), .Y(n2078) );
  INVX1 U2953 ( .A(n8857), .Y(n2079) );
  INVX1 U2954 ( .A(n9205), .Y(n2080) );
  INVX1 U2955 ( .A(n9308), .Y(n2081) );
  INVX1 U2956 ( .A(n9624), .Y(n2082) );
  INVX1 U2957 ( .A(n9653), .Y(n2083) );
  INVX1 U2958 ( .A(n9893), .Y(n2084) );
  INVX1 U2959 ( .A(n10245), .Y(n2085) );
  INVX1 U2960 ( .A(n10590), .Y(n2086) );
  BUFX2 U2961 ( .A(n6541), .Y(n2087) );
  BUFX2 U2962 ( .A(n6562), .Y(n2088) );
  BUFX2 U2963 ( .A(n6588), .Y(n2089) );
  BUFX2 U2964 ( .A(n6599), .Y(n2090) );
  BUFX2 U2965 ( .A(n6617), .Y(n2091) );
  BUFX2 U2966 ( .A(n6666), .Y(n2092) );
  BUFX2 U2967 ( .A(n6676), .Y(n2093) );
  BUFX2 U2968 ( .A(n6695), .Y(n2094) );
  BUFX2 U2969 ( .A(n6763), .Y(n2095) );
  BUFX2 U2970 ( .A(n6819), .Y(n2096) );
  BUFX2 U2971 ( .A(n6831), .Y(n2097) );
  BUFX2 U2972 ( .A(n6841), .Y(n2098) );
  BUFX2 U2973 ( .A(n6882), .Y(n2099) );
  BUFX2 U2974 ( .A(n7002), .Y(n2100) );
  BUFX2 U2975 ( .A(n7059), .Y(n2101) );
  BUFX2 U2976 ( .A(n7100), .Y(n2102) );
  BUFX2 U2977 ( .A(n7111), .Y(n2103) );
  BUFX2 U2978 ( .A(n7129), .Y(n2104) );
  BUFX2 U2979 ( .A(n7176), .Y(n2105) );
  BUFX2 U2980 ( .A(n7186), .Y(n2106) );
  BUFX2 U2981 ( .A(n7204), .Y(n2107) );
  BUFX2 U2982 ( .A(n7270), .Y(n2108) );
  BUFX2 U2983 ( .A(n7282), .Y(n2109) );
  BUFX2 U2984 ( .A(n7294), .Y(n2110) );
  BUFX2 U2985 ( .A(n7332), .Y(n2111) );
  BUFX2 U2986 ( .A(n7349), .Y(n2112) );
  BUFX2 U2987 ( .A(n7367), .Y(n2113) );
  BUFX2 U2988 ( .A(n7379), .Y(n2114) );
  INVX1 U2989 ( .A(n7574), .Y(n2115) );
  INVX1 U2990 ( .A(n2115), .Y(n2116) );
  BUFX2 U2991 ( .A(n7595), .Y(n2117) );
  BUFX2 U2992 ( .A(n7620), .Y(n2118) );
  BUFX2 U2993 ( .A(n7630), .Y(n2119) );
  BUFX2 U2994 ( .A(n7648), .Y(n2120) );
  BUFX2 U2995 ( .A(n7695), .Y(n2121) );
  BUFX2 U2996 ( .A(n7705), .Y(n2122) );
  BUFX2 U2997 ( .A(n7723), .Y(n2123) );
  BUFX2 U2998 ( .A(n7785), .Y(n2124) );
  INVX1 U2999 ( .A(n7836), .Y(n2125) );
  INVX1 U3000 ( .A(n2125), .Y(n2126) );
  BUFX2 U3001 ( .A(n7848), .Y(n2127) );
  BUFX2 U3002 ( .A(n7858), .Y(n2128) );
  BUFX2 U3003 ( .A(n7901), .Y(n2129) );
  BUFX2 U3004 ( .A(n7914), .Y(n2130) );
  BUFX2 U3005 ( .A(n7937), .Y(n2131) );
  BUFX2 U3006 ( .A(n7964), .Y(n2132) );
  BUFX2 U3007 ( .A(n8072), .Y(n2133) );
  BUFX2 U3008 ( .A(n8085), .Y(n2134) );
  BUFX2 U3009 ( .A(n8095), .Y(n2135) );
  BUFX2 U3010 ( .A(n8147), .Y(n2136) );
  BUFX2 U3011 ( .A(n8193), .Y(n2137) );
  BUFX2 U3012 ( .A(n8203), .Y(n2138) );
  BUFX2 U3013 ( .A(n8221), .Y(n2139) );
  BUFX2 U3014 ( .A(n8297), .Y(n2140) );
  BUFX2 U3015 ( .A(n8310), .Y(n2141) );
  INVX1 U3016 ( .A(n8348), .Y(n2142) );
  INVX1 U3017 ( .A(n2142), .Y(n2143) );
  BUFX2 U3018 ( .A(n8366), .Y(n2144) );
  BUFX2 U3019 ( .A(n8383), .Y(n2145) );
  BUFX2 U3020 ( .A(n8393), .Y(n2146) );
  BUFX2 U3021 ( .A(n8423), .Y(n2147) );
  BUFX2 U3022 ( .A(n8443), .Y(n2148) );
  BUFX2 U3023 ( .A(n8578), .Y(n2149) );
  BUFX2 U3024 ( .A(n8597), .Y(n2150) );
  BUFX2 U3025 ( .A(n8622), .Y(n2151) );
  BUFX2 U3026 ( .A(n8632), .Y(n2152) );
  BUFX2 U3027 ( .A(n8650), .Y(n2153) );
  BUFX2 U3028 ( .A(n8792), .Y(n2154) );
  BUFX2 U3029 ( .A(n8844), .Y(n2155) );
  BUFX2 U3030 ( .A(n8856), .Y(n2156) );
  BUFX2 U3031 ( .A(n8866), .Y(n2157) );
  BUFX2 U3032 ( .A(n8907), .Y(n2158) );
  BUFX2 U3033 ( .A(n9026), .Y(n2159) );
  BUFX2 U3034 ( .A(n9084), .Y(n2160) );
  BUFX2 U3035 ( .A(n9097), .Y(n2161) );
  BUFX2 U3036 ( .A(n9107), .Y(n2162) );
  BUFX2 U3037 ( .A(n9159), .Y(n2163) );
  BUFX2 U3038 ( .A(n9204), .Y(n2164) );
  BUFX2 U3039 ( .A(n9214), .Y(n2165) );
  BUFX2 U3040 ( .A(n9233), .Y(n2294) );
  INVX1 U3041 ( .A(n9295), .Y(n2295) );
  INVX1 U3042 ( .A(n2295), .Y(n2296) );
  BUFX2 U3043 ( .A(n9358), .Y(n2297) );
  BUFX2 U3044 ( .A(n9376), .Y(n2298) );
  BUFX2 U3045 ( .A(n9393), .Y(n2299) );
  INVX1 U3046 ( .A(n9403), .Y(n2300) );
  INVX1 U3047 ( .A(n2300), .Y(n2301) );
  BUFX2 U3048 ( .A(n9602), .Y(n2302) );
  BUFX2 U3049 ( .A(n9623), .Y(n2303) );
  BUFX2 U3050 ( .A(n9652), .Y(n2304) );
  BUFX2 U3051 ( .A(n9662), .Y(n2305) );
  BUFX2 U3052 ( .A(n9680), .Y(n2306) );
  BUFX2 U3053 ( .A(n9729), .Y(n2307) );
  BUFX2 U3054 ( .A(n9740), .Y(n2308) );
  BUFX2 U3055 ( .A(n9758), .Y(n2309) );
  BUFX2 U3056 ( .A(n9826), .Y(n2310) );
  INVX1 U3057 ( .A(n9880), .Y(n2311) );
  INVX1 U3058 ( .A(n2311), .Y(n2312) );
  BUFX2 U3059 ( .A(n9892), .Y(n2313) );
  BUFX2 U3060 ( .A(n9902), .Y(n2314) );
  BUFX2 U3061 ( .A(n9946), .Y(n2315) );
  BUFX2 U3062 ( .A(n9959), .Y(n2316) );
  BUFX2 U3063 ( .A(n9983), .Y(n2317) );
  BUFX2 U3064 ( .A(n10010), .Y(n2318) );
  BUFX2 U3065 ( .A(n10124), .Y(n2319) );
  BUFX2 U3066 ( .A(n10137), .Y(n2320) );
  BUFX2 U3067 ( .A(n10147), .Y(n2321) );
  BUFX2 U3068 ( .A(n10199), .Y(n2322) );
  BUFX2 U3069 ( .A(n10244), .Y(n2323) );
  BUFX2 U3070 ( .A(n10254), .Y(n2324) );
  INVX1 U3071 ( .A(n10273), .Y(n2325) );
  INVX1 U3072 ( .A(n2325), .Y(n2326) );
  INVX1 U3073 ( .A(n10340), .Y(n2327) );
  INVX1 U3074 ( .A(n2327), .Y(n2328) );
  BUFX2 U3075 ( .A(n10352), .Y(n2329) );
  BUFX2 U3076 ( .A(n10365), .Y(n2330) );
  BUFX2 U3077 ( .A(n10428), .Y(n2331) );
  BUFX2 U3078 ( .A(n10445), .Y(n2332) );
  BUFX2 U3079 ( .A(n10457), .Y(n2333) );
  BUFX2 U3080 ( .A(n10526), .Y(n2334) );
  INVX1 U3081 ( .A(n6647), .Y(n2335) );
  INVX1 U3082 ( .A(n7675), .Y(n2336) );
  INVX1 U3083 ( .A(n8459), .Y(n2337) );
  INVX1 U3084 ( .A(n9708), .Y(n2338) );
  AND2X2 U3085 ( .A(n1143), .B(n1487), .Y(n10589) );
  INVX1 U3086 ( .A(n10589), .Y(n2339) );
  BUFX2 U3087 ( .A(n8689), .Y(n2340) );
  INVX1 U3088 ( .A(n9464), .Y(n2341) );
  BUFX2 U3089 ( .A(n7170), .Y(n2342) );
  BUFX2 U3090 ( .A(n7441), .Y(n2343) );
  BUFX2 U3091 ( .A(n7445), .Y(n2344) );
  BUFX2 U3092 ( .A(n7449), .Y(n2345) );
  BUFX2 U3093 ( .A(n8166), .Y(n2346) );
  INVX1 U3094 ( .A(n2348), .Y(n2347) );
  BUFX2 U3095 ( .A(n8476), .Y(n2348) );
  BUFX2 U3096 ( .A(n9178), .Y(n2349) );
  BUFX2 U3097 ( .A(n9517), .Y(n2350) );
  BUFX2 U3098 ( .A(n9521), .Y(n2351) );
  BUFX2 U3099 ( .A(n9525), .Y(n2352) );
  BUFX2 U3100 ( .A(n9529), .Y(n2353) );
  BUFX2 U3101 ( .A(n10485), .Y(n2354) );
  BUFX2 U3102 ( .A(n10494), .Y(n2355) );
  BUFX2 U3103 ( .A(n10516), .Y(n2356) );
  BUFX2 U3104 ( .A(n10531), .Y(n2357) );
  BUFX2 U3105 ( .A(n10535), .Y(n2358) );
  BUFX2 U3106 ( .A(n10573), .Y(n2359) );
  BUFX2 U3107 ( .A(n10584), .Y(n2360) );
  BUFX2 U3108 ( .A(n10594), .Y(n2361) );
  INVX1 U3109 ( .A(n10598), .Y(n2362) );
  INVX1 U3110 ( .A(n6549), .Y(n2363) );
  OR2X1 U3111 ( .A(n6282), .B(n6153), .Y(n6568) );
  INVX1 U3112 ( .A(n6568), .Y(n2364) );
  OR2X1 U3113 ( .A(n5948), .B(n6172), .Y(n7066) );
  INVX1 U3114 ( .A(n7066), .Y(n2365) );
  INVX1 U3115 ( .A(n7420), .Y(n2366) );
  INVX1 U3116 ( .A(n7433), .Y(n2367) );
  OR2X1 U3117 ( .A(n6297), .B(n6188), .Y(n7584) );
  INVX1 U3118 ( .A(n7584), .Y(n2368) );
  OR2X1 U3119 ( .A(n6297), .B(n6153), .Y(n7601) );
  INVX1 U3120 ( .A(n7601), .Y(n2369) );
  INVX1 U3121 ( .A(n8101), .Y(n2370) );
  OR2X1 U3122 ( .A(n6325), .B(n6218), .Y(n8586) );
  INVX1 U3123 ( .A(n8586), .Y(n2371) );
  OR2X1 U3124 ( .A(n6325), .B(n6153), .Y(n8603) );
  INVX1 U3125 ( .A(n8603), .Y(n2372) );
  OR2X1 U3126 ( .A(n6024), .B(n6231), .Y(n9113) );
  INVX1 U3127 ( .A(n9113), .Y(n2373) );
  OR2X1 U3128 ( .A(n6345), .B(n6244), .Y(n9612) );
  INVX1 U3129 ( .A(n9612), .Y(n2374) );
  OR2X1 U3130 ( .A(n6064), .B(n6355), .Y(n9625) );
  INVX1 U3131 ( .A(n9625), .Y(n2375) );
  OR2X1 U3132 ( .A(n6345), .B(n6153), .Y(n9631) );
  INVX1 U3133 ( .A(n9631), .Y(n2376) );
  INVX1 U3134 ( .A(n10153), .Y(n2377) );
  BUFX2 U3135 ( .A(n6477), .Y(n2378) );
  BUFX2 U3136 ( .A(n6540), .Y(n2379) );
  BUFX2 U3137 ( .A(n6616), .Y(n2380) );
  BUFX2 U3138 ( .A(n6561), .Y(n2381) );
  BUFX2 U3139 ( .A(n6587), .Y(n2382) );
  BUFX2 U3140 ( .A(n6598), .Y(n2383) );
  BUFX2 U3141 ( .A(n6623), .Y(n2384) );
  BUFX2 U3142 ( .A(n6639), .Y(n2385) );
  BUFX2 U3143 ( .A(n6654), .Y(n2386) );
  BUFX2 U3144 ( .A(n6665), .Y(n2387) );
  BUFX2 U3145 ( .A(n6675), .Y(n2388) );
  BUFX2 U3146 ( .A(n6694), .Y(n2389) );
  BUFX2 U3147 ( .A(n6701), .Y(n2390) );
  BUFX2 U3148 ( .A(n6752), .Y(n2391) );
  BUFX2 U3149 ( .A(n6762), .Y(n2392) );
  BUFX2 U3150 ( .A(n6800), .Y(n2393) );
  BUFX2 U3151 ( .A(n6818), .Y(n2394) );
  BUFX2 U3152 ( .A(n6830), .Y(n2395) );
  BUFX2 U3153 ( .A(n6840), .Y(n2396) );
  BUFX2 U3154 ( .A(n6881), .Y(n2397) );
  BUFX2 U3155 ( .A(n7001), .Y(n2398) );
  BUFX2 U3156 ( .A(n7008), .Y(n2399) );
  BUFX2 U3157 ( .A(n7058), .Y(n2400) );
  BUFX2 U3158 ( .A(n7065), .Y(n2401) );
  BUFX2 U3159 ( .A(n7096), .Y(n2402) );
  BUFX2 U3160 ( .A(n7099), .Y(n2403) );
  BUFX2 U3161 ( .A(n7107), .Y(n2404) );
  BUFX2 U3162 ( .A(n7110), .Y(n2405) );
  BUFX2 U3163 ( .A(n7128), .Y(n2406) );
  BUFX2 U3164 ( .A(n7166), .Y(n2407) );
  BUFX2 U3165 ( .A(n7175), .Y(n2408) );
  BUFX2 U3166 ( .A(n7185), .Y(n2409) );
  BUFX2 U3167 ( .A(n7203), .Y(n2410) );
  BUFX2 U3168 ( .A(n7269), .Y(n2411) );
  BUFX2 U3169 ( .A(n7293), .Y(n2412) );
  BUFX2 U3170 ( .A(n7331), .Y(n2413) );
  BUFX2 U3171 ( .A(n7344), .Y(n2414) );
  BUFX2 U3172 ( .A(n7357), .Y(n2415) );
  BUFX2 U3173 ( .A(n7366), .Y(n2416) );
  BUFX2 U3174 ( .A(n7378), .Y(n2417) );
  INVX1 U3175 ( .A(n7396), .Y(n2418) );
  INVX1 U3176 ( .A(n2418), .Y(n2419) );
  BUFX2 U3177 ( .A(n7444), .Y(n2420) );
  BUFX2 U3178 ( .A(n7462), .Y(n2421) );
  BUFX2 U3179 ( .A(n7508), .Y(n2422) );
  BUFX2 U3180 ( .A(n7521), .Y(n2423) );
  INVX1 U3181 ( .A(n7573), .Y(n2424) );
  INVX1 U3182 ( .A(n2424), .Y(n2425) );
  BUFX2 U3183 ( .A(n7580), .Y(n2426) );
  BUFX2 U3184 ( .A(n7594), .Y(n2427) );
  BUFX2 U3185 ( .A(n7619), .Y(n2428) );
  BUFX2 U3186 ( .A(n7629), .Y(n2429) );
  BUFX2 U3187 ( .A(n7647), .Y(n2430) );
  BUFX2 U3188 ( .A(n7654), .Y(n2431) );
  BUFX2 U3189 ( .A(n7667), .Y(n2432) );
  BUFX2 U3190 ( .A(n7682), .Y(n2433) );
  BUFX2 U3191 ( .A(n7694), .Y(n2434) );
  BUFX2 U3192 ( .A(n7704), .Y(n2435) );
  BUFX2 U3193 ( .A(n7722), .Y(n2436) );
  BUFX2 U3194 ( .A(n7729), .Y(n2437) );
  BUFX2 U3195 ( .A(n7784), .Y(n2438) );
  BUFX2 U3196 ( .A(n7791), .Y(n2439) );
  BUFX2 U3197 ( .A(n7835), .Y(n2440) );
  BUFX2 U3198 ( .A(n7842), .Y(n2441) );
  BUFX2 U3199 ( .A(n7847), .Y(n2442) );
  BUFX2 U3200 ( .A(n7857), .Y(n2443) );
  BUFX2 U3201 ( .A(n7900), .Y(n2444) );
  BUFX2 U3202 ( .A(n7907), .Y(n2445) );
  BUFX2 U3203 ( .A(n7910), .Y(n2446) );
  BUFX2 U3204 ( .A(n7929), .Y(n2447) );
  BUFX2 U3205 ( .A(n7936), .Y(n2448) );
  BUFX2 U3206 ( .A(n7963), .Y(n2449) );
  BUFX2 U3207 ( .A(n7970), .Y(n2450) );
  BUFX2 U3208 ( .A(n8021), .Y(n2451) );
  BUFX2 U3209 ( .A(n8071), .Y(n2452) );
  BUFX2 U3210 ( .A(n8078), .Y(n2453) );
  BUFX2 U3211 ( .A(n8081), .Y(n2454) );
  BUFX2 U3212 ( .A(n8084), .Y(n2455) );
  BUFX2 U3213 ( .A(n8094), .Y(n2456) );
  BUFX2 U3214 ( .A(n8146), .Y(n2457) );
  BUFX2 U3215 ( .A(n8153), .Y(n2458) );
  BUFX2 U3216 ( .A(n8192), .Y(n2459) );
  BUFX2 U3217 ( .A(n8202), .Y(n2460) );
  BUFX2 U3218 ( .A(n8220), .Y(n2461) );
  BUFX2 U3219 ( .A(n8227), .Y(n2462) );
  BUFX2 U3220 ( .A(n8269), .Y(n2463) );
  INVX1 U3221 ( .A(n8284), .Y(n2464) );
  INVX1 U3222 ( .A(n2464), .Y(n2465) );
  BUFX2 U3223 ( .A(n8291), .Y(n2466) );
  BUFX2 U3224 ( .A(n8296), .Y(n2467) );
  BUFX2 U3225 ( .A(n8309), .Y(n2468) );
  BUFX2 U3226 ( .A(n8347), .Y(n2469) );
  BUFX2 U3227 ( .A(n8354), .Y(n2470) );
  BUFX2 U3228 ( .A(n8360), .Y(n2471) );
  BUFX2 U3229 ( .A(n8373), .Y(n2472) );
  BUFX2 U3230 ( .A(n8382), .Y(n2473) );
  BUFX2 U3231 ( .A(n8392), .Y(n2474) );
  BUFX2 U3232 ( .A(n8422), .Y(n2475) );
  BUFX2 U3233 ( .A(n8442), .Y(n2476) );
  BUFX2 U3234 ( .A(n8450), .Y(n2477) );
  BUFX2 U3235 ( .A(n8520), .Y(n2478) );
  BUFX2 U3236 ( .A(n8475), .Y(n2479) );
  BUFX2 U3237 ( .A(n8514), .Y(n2480) );
  BUFX2 U3238 ( .A(n8525), .Y(n2481) );
  BUFX2 U3239 ( .A(n8577), .Y(n2482) );
  BUFX2 U3240 ( .A(n8582), .Y(n2483) );
  BUFX2 U3241 ( .A(n8649), .Y(n2484) );
  BUFX2 U3242 ( .A(n8596), .Y(n2485) );
  BUFX2 U3243 ( .A(n8621), .Y(n2486) );
  BUFX2 U3244 ( .A(n8631), .Y(n2615) );
  BUFX2 U3245 ( .A(n8735), .Y(n2616) );
  BUFX2 U3246 ( .A(n8791), .Y(n2617) );
  BUFX2 U3247 ( .A(n8798), .Y(n2618) );
  BUFX2 U3248 ( .A(n8826), .Y(n2619) );
  BUFX2 U3249 ( .A(n8843), .Y(n2620) );
  BUFX2 U3250 ( .A(n8850), .Y(n2621) );
  BUFX2 U3251 ( .A(n8855), .Y(n2622) );
  BUFX2 U3252 ( .A(n8865), .Y(n2623) );
  BUFX2 U3253 ( .A(n8906), .Y(n2624) );
  BUFX2 U3254 ( .A(n8983), .Y(n2625) );
  BUFX2 U3255 ( .A(n9025), .Y(n2626) );
  BUFX2 U3256 ( .A(n9064), .Y(n2627) );
  BUFX2 U3257 ( .A(n9083), .Y(n2628) );
  BUFX2 U3258 ( .A(n9106), .Y(n2629) );
  BUFX2 U3259 ( .A(n9158), .Y(n2630) );
  BUFX2 U3260 ( .A(n9203), .Y(n2631) );
  BUFX2 U3261 ( .A(n9213), .Y(n2632) );
  BUFX2 U3262 ( .A(n9220), .Y(n2633) );
  BUFX2 U3263 ( .A(n9232), .Y(n2634) );
  BUFX2 U3264 ( .A(n9294), .Y(n2635) );
  BUFX2 U3265 ( .A(n9319), .Y(n2636) );
  BUFX2 U3266 ( .A(n9357), .Y(n2637) );
  BUFX2 U3267 ( .A(n9370), .Y(n2638) );
  BUFX2 U3268 ( .A(n9383), .Y(n2639) );
  BUFX2 U3269 ( .A(n9392), .Y(n2640) );
  BUFX2 U3270 ( .A(n9402), .Y(n2641) );
  BUFX2 U3271 ( .A(n9472), .Y(n2642) );
  BUFX2 U3272 ( .A(n9520), .Y(n2643) );
  BUFX2 U3273 ( .A(n9548), .Y(n2644) );
  BUFX2 U3274 ( .A(n9601), .Y(n2645) );
  BUFX2 U3275 ( .A(n9608), .Y(n2646) );
  BUFX2 U3276 ( .A(n9622), .Y(n2647) );
  BUFX2 U3277 ( .A(n9651), .Y(n2648) );
  BUFX2 U3278 ( .A(n9661), .Y(n2649) );
  BUFX2 U3279 ( .A(n9679), .Y(n2650) );
  BUFX2 U3280 ( .A(n9686), .Y(n2651) );
  BUFX2 U3281 ( .A(n9699), .Y(n2652) );
  BUFX2 U3282 ( .A(n9715), .Y(n2653) );
  BUFX2 U3283 ( .A(n9728), .Y(n2654) );
  BUFX2 U3284 ( .A(n9739), .Y(n2655) );
  BUFX2 U3285 ( .A(n9757), .Y(n2656) );
  BUFX2 U3286 ( .A(n9764), .Y(n2657) );
  BUFX2 U3287 ( .A(n9825), .Y(n2658) );
  BUFX2 U3288 ( .A(n9832), .Y(n2659) );
  BUFX2 U3289 ( .A(n9879), .Y(n2660) );
  BUFX2 U3290 ( .A(n9886), .Y(n2661) );
  BUFX2 U3291 ( .A(n9891), .Y(n2662) );
  BUFX2 U3292 ( .A(n9901), .Y(n2663) );
  BUFX2 U3293 ( .A(n9945), .Y(n2664) );
  BUFX2 U3294 ( .A(n9952), .Y(n2665) );
  BUFX2 U3295 ( .A(n9955), .Y(n2666) );
  BUFX2 U3296 ( .A(n9958), .Y(n2667) );
  BUFX2 U3297 ( .A(n9975), .Y(n2668) );
  BUFX2 U3298 ( .A(n9982), .Y(n2669) );
  BUFX2 U3299 ( .A(n10009), .Y(n2670) );
  BUFX2 U3300 ( .A(n10016), .Y(n2671) );
  BUFX2 U3301 ( .A(n10123), .Y(n2672) );
  BUFX2 U3302 ( .A(n10130), .Y(n2673) );
  BUFX2 U3303 ( .A(n10133), .Y(n2674) );
  BUFX2 U3304 ( .A(n10136), .Y(n2675) );
  BUFX2 U3305 ( .A(n10146), .Y(n2676) );
  BUFX2 U3306 ( .A(n10198), .Y(n2677) );
  BUFX2 U3307 ( .A(n10205), .Y(n2678) );
  BUFX2 U3308 ( .A(n10243), .Y(n2679) );
  BUFX2 U3309 ( .A(n10253), .Y(n2680) );
  BUFX2 U3310 ( .A(n10260), .Y(n2681) );
  BUFX2 U3311 ( .A(n10272), .Y(n2682) );
  BUFX2 U3312 ( .A(n10279), .Y(n2683) );
  INVX1 U3313 ( .A(n10339), .Y(n2684) );
  INVX1 U3314 ( .A(n2684), .Y(n2685) );
  BUFX2 U3315 ( .A(n10346), .Y(n2686) );
  BUFX2 U3316 ( .A(n10351), .Y(n2687) );
  BUFX2 U3317 ( .A(n10364), .Y(n2688) );
  BUFX2 U3318 ( .A(n10416), .Y(n2689) );
  BUFX2 U3319 ( .A(n10422), .Y(n2690) );
  BUFX2 U3320 ( .A(n10435), .Y(n2691) );
  BUFX2 U3321 ( .A(n10444), .Y(n2692) );
  BUFX2 U3322 ( .A(n10456), .Y(n2693) );
  BUFX2 U3323 ( .A(n10484), .Y(n2694) );
  BUFX2 U3324 ( .A(n10546), .Y(n2695) );
  BUFX2 U3325 ( .A(n10515), .Y(n2696) );
  BUFX2 U3326 ( .A(n10525), .Y(n2697) );
  BUFX2 U3327 ( .A(n6985), .Y(n2698) );
  BUFX2 U3328 ( .A(n7227), .Y(n2699) );
  BUFX2 U3329 ( .A(n7448), .Y(n2700) );
  BUFX2 U3330 ( .A(n7452), .Y(n2701) );
  BUFX2 U3331 ( .A(n7456), .Y(n2702) );
  BUFX2 U3332 ( .A(n7495), .Y(n2703) );
  BUFX2 U3333 ( .A(n8500), .Y(n2704) );
  BUFX2 U3334 ( .A(n9512), .Y(n2705) );
  BUFX2 U3335 ( .A(n9524), .Y(n2706) );
  BUFX2 U3336 ( .A(n9528), .Y(n2707) );
  BUFX2 U3337 ( .A(n9532), .Y(n2708) );
  INVX1 U3338 ( .A(n10550), .Y(n2709) );
  INVX1 U3339 ( .A(n2709), .Y(n2710) );
  BUFX2 U3340 ( .A(n10530), .Y(n2711) );
  BUFX2 U3341 ( .A(n10534), .Y(n2712) );
  BUFX2 U3342 ( .A(n10538), .Y(n2713) );
  BUFX2 U3343 ( .A(n10560), .Y(n2714) );
  BUFX2 U3344 ( .A(n10572), .Y(n2715) );
  BUFX2 U3345 ( .A(n10593), .Y(n2716) );
  BUFX2 U3346 ( .A(n10597), .Y(n2717) );
  INVX1 U3347 ( .A(n6610), .Y(n2718) );
  INVX1 U3348 ( .A(n6688), .Y(n2719) );
  INVX1 U3349 ( .A(n6875), .Y(n2720) );
  AND2X1 U3350 ( .A(n6169), .B(n6285), .Y(n7169) );
  INVX1 U3351 ( .A(n7169), .Y(n2721) );
  AND2X1 U3352 ( .A(n7070), .B(n6288), .Y(n7242) );
  INVX1 U3353 ( .A(n7242), .Y(n2722) );
  INVX1 U3354 ( .A(n7325), .Y(n2723) );
  INVX1 U3355 ( .A(n7390), .Y(n2724) );
  INVX1 U3356 ( .A(n7641), .Y(n2725) );
  INVX1 U3357 ( .A(n7716), .Y(n2726) );
  AND2X1 U3358 ( .A(n6730), .B(n5989), .Y(n7810) );
  INVX1 U3359 ( .A(n7810), .Y(n2727) );
  INVX1 U3360 ( .A(n7894), .Y(n2728) );
  INVX1 U3361 ( .A(n7957), .Y(n2729) );
  INVX1 U3362 ( .A(n8140), .Y(n2730) );
  AND2X1 U3363 ( .A(n10290), .B(n8413), .Y(n8160) );
  INVX1 U3364 ( .A(n8160), .Y(n2731) );
  AND2X1 U3365 ( .A(n6201), .B(n6300), .Y(n8165) );
  INVX1 U3366 ( .A(n8165), .Y(n2732) );
  AND2X1 U3367 ( .A(n8115), .B(n8238), .Y(n8240) );
  INVX1 U3368 ( .A(n8240), .Y(n2733) );
  AND2X1 U3369 ( .A(n8102), .B(n6305), .Y(n8256) );
  INVX1 U3370 ( .A(n8256), .Y(n2734) );
  INVX1 U3371 ( .A(n8341), .Y(n2735) );
  INVX1 U3372 ( .A(n8404), .Y(n2736) );
  INVX1 U3373 ( .A(n8643), .Y(n2737) );
  AND2X1 U3374 ( .A(n6319), .B(n9793), .Y(n8688) );
  INVX1 U3375 ( .A(n8688), .Y(n2738) );
  INVX1 U3376 ( .A(n8900), .Y(n2739) );
  INVX1 U3377 ( .A(n9152), .Y(n2740) );
  AND2X1 U3378 ( .A(n10290), .B(n9473), .Y(n9172) );
  INVX1 U3379 ( .A(n9172), .Y(n2741) );
  INVX1 U3380 ( .A(n9177), .Y(n2742) );
  AND2X1 U3381 ( .A(n9127), .B(n9250), .Y(n9251) );
  INVX1 U3382 ( .A(n9251), .Y(n2743) );
  AND2X1 U3383 ( .A(n9114), .B(n5286), .Y(n9267) );
  INVX1 U3384 ( .A(n9267), .Y(n2744) );
  INVX1 U3385 ( .A(n9351), .Y(n2745) );
  INVX1 U3386 ( .A(n9415), .Y(n2746) );
  INVX1 U3387 ( .A(n9673), .Y(n2747) );
  INVX1 U3388 ( .A(n9751), .Y(n2748) );
  AND2X1 U3389 ( .A(n6730), .B(n6061), .Y(n9852) );
  INVX1 U3390 ( .A(n9852), .Y(n2749) );
  INVX1 U3391 ( .A(n9939), .Y(n2750) );
  INVX1 U3392 ( .A(n10003), .Y(n2751) );
  INVX1 U3393 ( .A(n10192), .Y(n2752) );
  AND2X1 U3394 ( .A(n10290), .B(n10495), .Y(n10212) );
  INVX1 U3395 ( .A(n10212), .Y(n2753) );
  AND2X1 U3396 ( .A(n10167), .B(n10292), .Y(n10293) );
  INVX1 U3397 ( .A(n10293), .Y(n2754) );
  AND2X1 U3398 ( .A(n6054), .B(n10154), .Y(n10309) );
  INVX1 U3399 ( .A(n10309), .Y(n2755) );
  INVX1 U3400 ( .A(n10403), .Y(n2756) );
  INVX1 U3401 ( .A(n10470), .Y(n2757) );
  INVX1 U3402 ( .A(n10583), .Y(n2758) );
  BUFX2 U3403 ( .A(n6915), .Y(n2759) );
  BUFX2 U3404 ( .A(n7083), .Y(n2760) );
  BUFX2 U3405 ( .A(n8941), .Y(n2761) );
  BUFX2 U3406 ( .A(n9452), .Y(n2762) );
  BUFX2 U3407 ( .A(n6479), .Y(n2763) );
  BUFX2 U3408 ( .A(n7030), .Y(n2764) );
  BUFX2 U3409 ( .A(n7523), .Y(n2765) );
  BUFX2 U3410 ( .A(n8043), .Y(n2766) );
  BUFX2 U3411 ( .A(n8108), .Y(n2767) );
  BUFX2 U3412 ( .A(n8527), .Y(n2768) );
  BUFX2 U3413 ( .A(n9054), .Y(n2769) );
  BUFX2 U3414 ( .A(n9120), .Y(n2770) );
  BUFX2 U3415 ( .A(n9550), .Y(n2771) );
  BUFX2 U3416 ( .A(n10092), .Y(n2772) );
  BUFX2 U3417 ( .A(n10160), .Y(n2773) );
  BUFX2 U3418 ( .A(n7228), .Y(n2774) );
  AND2X1 U3419 ( .A(n5741), .B(n5631), .Y(n6727) );
  INVX1 U3420 ( .A(n6727), .Y(n2775) );
  AND2X1 U3421 ( .A(n10383), .B(n5563), .Y(n7307) );
  INVX1 U3422 ( .A(n7307), .Y(n2776) );
  AND2X1 U3423 ( .A(n5741), .B(n5630), .Y(n7752) );
  INVX1 U3424 ( .A(n7752), .Y(n2777) );
  AND2X1 U3425 ( .A(n10383), .B(n4700), .Y(n8323) );
  INVX1 U3426 ( .A(n8323), .Y(n2778) );
  AND2X1 U3427 ( .A(n5741), .B(n5711), .Y(n8759) );
  INVX1 U3428 ( .A(n8759), .Y(n2779) );
  AND2X1 U3429 ( .A(n10383), .B(n4701), .Y(n9333) );
  INVX1 U3430 ( .A(n9333), .Y(n2780) );
  AND2X1 U3431 ( .A(n5741), .B(n4702), .Y(n9788) );
  INVX1 U3432 ( .A(n9788), .Y(n2781) );
  AND2X1 U3433 ( .A(n10383), .B(n4703), .Y(n10385) );
  INVX1 U3434 ( .A(n10385), .Y(n2782) );
  BUFX2 U3435 ( .A(n8107), .Y(n2783) );
  BUFX2 U3436 ( .A(n9119), .Y(n2784) );
  BUFX2 U3437 ( .A(n10159), .Y(n2785) );
  BUFX2 U3438 ( .A(n6521), .Y(n2786) );
  BUFX2 U3439 ( .A(n7044), .Y(n2787) );
  BUFX2 U3440 ( .A(n7287), .Y(n2788) );
  BUFX2 U3441 ( .A(n7372), .Y(n2789) );
  BUFX2 U3442 ( .A(n7496), .Y(n2790) );
  BUFX2 U3443 ( .A(n7554), .Y(n2791) );
  BUFX2 U3444 ( .A(n8057), .Y(n2792) );
  BUFX2 U3445 ( .A(n8303), .Y(n2793) );
  BUFX2 U3446 ( .A(n8386), .Y(n2794) );
  BUFX2 U3447 ( .A(n8436), .Y(n2795) );
  BUFX2 U3448 ( .A(n8501), .Y(n2796) );
  BUFX2 U3449 ( .A(n8558), .Y(n2797) );
  BUFX2 U3450 ( .A(n8664), .Y(n2798) );
  BUFX2 U3451 ( .A(n9068), .Y(n2799) );
  BUFX2 U3452 ( .A(n9313), .Y(n2800) );
  BUFX2 U3453 ( .A(n9396), .Y(n2801) );
  BUFX2 U3454 ( .A(n9444), .Y(n2802) );
  BUFX2 U3455 ( .A(n9513), .Y(n2803) );
  BUFX2 U3456 ( .A(n9581), .Y(n2804) );
  BUFX2 U3457 ( .A(n10108), .Y(n2805) );
  BUFX2 U3458 ( .A(n10358), .Y(n2806) );
  BUFX2 U3459 ( .A(n10450), .Y(n2807) );
  BUFX2 U3460 ( .A(n10561), .Y(n2936) );
  AND2X1 U3461 ( .A(n5264), .B(n6986), .Y(n6987) );
  INVX1 U3462 ( .A(n6987), .Y(n2937) );
  AND2X1 U3463 ( .A(n5264), .B(n7999), .Y(n8000) );
  INVX1 U3464 ( .A(n8000), .Y(n2938) );
  OR2X1 U3465 ( .A(n8262), .B(n10315), .Y(n8263) );
  INVX1 U3466 ( .A(n8263), .Y(n2939) );
  AND2X1 U3467 ( .A(n5264), .B(n9010), .Y(n9011) );
  INVX1 U3468 ( .A(n9011), .Y(n2940) );
  AND2X1 U3469 ( .A(n5264), .B(n10045), .Y(n10046) );
  INVX1 U3470 ( .A(n10046), .Y(n2941) );
  BUFX2 U3471 ( .A(n6689), .Y(n2942) );
  BUFX2 U3472 ( .A(n6876), .Y(n2943) );
  BUFX2 U3473 ( .A(n7123), .Y(n2944) );
  BUFX2 U3474 ( .A(n7198), .Y(n2945) );
  BUFX2 U3475 ( .A(n7326), .Y(n2946) );
  INVX1 U3476 ( .A(n7391), .Y(n2947) );
  INVX1 U3477 ( .A(n2947), .Y(n2948) );
  BUFX2 U3478 ( .A(n7457), .Y(n2949) );
  INVX1 U3479 ( .A(n7509), .Y(n2950) );
  INVX1 U3480 ( .A(n2950), .Y(n2951) );
  BUFX2 U3481 ( .A(n7642), .Y(n2952) );
  BUFX2 U3482 ( .A(n7717), .Y(n2953) );
  BUFX2 U3483 ( .A(n7895), .Y(n2954) );
  BUFX2 U3484 ( .A(n7958), .Y(n2955) );
  BUFX2 U3485 ( .A(n8141), .Y(n2956) );
  BUFX2 U3486 ( .A(n8215), .Y(n2957) );
  BUFX2 U3487 ( .A(n8342), .Y(n2958) );
  BUFX2 U3488 ( .A(n8704), .Y(n2959) );
  BUFX2 U3489 ( .A(n8901), .Y(n2960) );
  BUFX2 U3490 ( .A(n9153), .Y(n2961) );
  BUFX2 U3491 ( .A(n9227), .Y(n2962) );
  BUFX2 U3492 ( .A(n9352), .Y(n2963) );
  BUFX2 U3493 ( .A(n9674), .Y(n2964) );
  BUFX2 U3494 ( .A(n9752), .Y(n2965) );
  BUFX2 U3495 ( .A(n9940), .Y(n2966) );
  BUFX2 U3496 ( .A(n10004), .Y(n2967) );
  BUFX2 U3497 ( .A(n10193), .Y(n2968) );
  BUFX2 U3498 ( .A(n10267), .Y(n2969) );
  INVX1 U3499 ( .A(n10404), .Y(n2970) );
  INVX1 U3500 ( .A(n2970), .Y(n2971) );
  AND2X1 U3501 ( .A(n6534), .B(n6533), .Y(n6535) );
  INVX1 U3502 ( .A(n6535), .Y(n2972) );
  AND2X1 U3503 ( .A(n6756), .B(n6755), .Y(n6757) );
  INVX1 U3504 ( .A(n6757), .Y(n2973) );
  AND2X1 U3505 ( .A(n6812), .B(n6811), .Y(n6813) );
  INVX1 U3506 ( .A(n6813), .Y(n2974) );
  AND2X1 U3507 ( .A(n6995), .B(n6994), .Y(n6996) );
  INVX1 U3508 ( .A(n6996), .Y(n2975) );
  AND2X1 U3509 ( .A(n7052), .B(n7051), .Y(n7053) );
  INVX1 U3510 ( .A(n7053), .Y(n2976) );
  AND2X1 U3511 ( .A(n7263), .B(n7262), .Y(n7264) );
  INVX1 U3512 ( .A(n7264), .Y(n2977) );
  AND2X1 U3513 ( .A(n7567), .B(n7566), .Y(n7568) );
  INVX1 U3514 ( .A(n7568), .Y(n2978) );
  AND2X1 U3515 ( .A(n7778), .B(n7777), .Y(n7779) );
  INVX1 U3516 ( .A(n7779), .Y(n2979) );
  AND2X1 U3517 ( .A(n7829), .B(n7828), .Y(n7830) );
  INVX1 U3518 ( .A(n7830), .Y(n2980) );
  INVX1 U3519 ( .A(n8009), .Y(n2981) );
  AND2X1 U3520 ( .A(n8065), .B(n8064), .Y(n8066) );
  INVX1 U3521 ( .A(n8066), .Y(n2982) );
  INVX1 U3522 ( .A(n8162), .Y(n2983) );
  AND2X1 U3523 ( .A(n8278), .B(n8277), .Y(n8279) );
  INVX1 U3524 ( .A(n8279), .Y(n2984) );
  AND2X1 U3525 ( .A(n8571), .B(n8570), .Y(n8572) );
  INVX1 U3526 ( .A(n8572), .Y(n2985) );
  AND2X1 U3527 ( .A(n8785), .B(n8784), .Y(n8786) );
  INVX1 U3528 ( .A(n8786), .Y(n2986) );
  AND2X1 U3529 ( .A(n8837), .B(n8836), .Y(n8838) );
  INVX1 U3530 ( .A(n8838), .Y(n2987) );
  AND2X1 U3531 ( .A(n9019), .B(n9018), .Y(n9020) );
  INVX1 U3532 ( .A(n9020), .Y(n2988) );
  AND2X1 U3533 ( .A(n9077), .B(n9076), .Y(n9078) );
  INVX1 U3534 ( .A(n9078), .Y(n2989) );
  INVX1 U3535 ( .A(n9174), .Y(n2990) );
  AND2X1 U3536 ( .A(n9288), .B(n9287), .Y(n9289) );
  INVX1 U3537 ( .A(n9289), .Y(n2991) );
  AND2X1 U3538 ( .A(n9595), .B(n9594), .Y(n9596) );
  INVX1 U3539 ( .A(n9596), .Y(n2992) );
  AND2X1 U3540 ( .A(n9819), .B(n9818), .Y(n9820) );
  INVX1 U3541 ( .A(n9820), .Y(n2993) );
  AND2X1 U3542 ( .A(n9873), .B(n9872), .Y(n9874) );
  INVX1 U3543 ( .A(n9874), .Y(n2994) );
  INVX1 U3544 ( .A(n10055), .Y(n2995) );
  AND2X1 U3545 ( .A(n10117), .B(n10116), .Y(n10118) );
  INVX1 U3546 ( .A(n10118), .Y(n2996) );
  INVX1 U3547 ( .A(n10214), .Y(n2997) );
  AND2X1 U3548 ( .A(n10333), .B(n10332), .Y(n10334) );
  INVX1 U3549 ( .A(n10334), .Y(n2998) );
  BUFX2 U3550 ( .A(n6539), .Y(n2999) );
  BUFX2 U3551 ( .A(n6693), .Y(n3000) );
  BUFX2 U3552 ( .A(n6761), .Y(n3001) );
  BUFX2 U3553 ( .A(n7057), .Y(n3002) );
  BUFX2 U3554 ( .A(n7127), .Y(n3003) );
  BUFX2 U3555 ( .A(n7202), .Y(n3004) );
  BUFX2 U3556 ( .A(n7268), .Y(n3005) );
  BUFX2 U3557 ( .A(n7330), .Y(n3006) );
  BUFX2 U3558 ( .A(n7395), .Y(n3007) );
  BUFX2 U3559 ( .A(n7461), .Y(n3008) );
  BUFX2 U3560 ( .A(n7646), .Y(n3009) );
  BUFX2 U3561 ( .A(n7721), .Y(n3010) );
  BUFX2 U3562 ( .A(n7783), .Y(n3011) );
  BUFX2 U3563 ( .A(n7834), .Y(n3012) );
  BUFX2 U3564 ( .A(n7899), .Y(n3013) );
  BUFX2 U3565 ( .A(n7962), .Y(n3014) );
  BUFX2 U3566 ( .A(n8013), .Y(n3015) );
  BUFX2 U3567 ( .A(n8070), .Y(n3016) );
  BUFX2 U3568 ( .A(n8121), .Y(n3017) );
  BUFX2 U3569 ( .A(n8145), .Y(n3018) );
  BUFX2 U3570 ( .A(n8219), .Y(n3019) );
  BUFX2 U3571 ( .A(n8268), .Y(n3020) );
  BUFX2 U3572 ( .A(n8283), .Y(n3021) );
  BUFX2 U3573 ( .A(n8346), .Y(n3022) );
  INVX1 U3574 ( .A(n8409), .Y(n3023) );
  INVX1 U3575 ( .A(n3023), .Y(n3024) );
  BUFX2 U3576 ( .A(n8464), .Y(n3025) );
  BUFX2 U3577 ( .A(n8474), .Y(n3026) );
  BUFX2 U3578 ( .A(n8576), .Y(n3027) );
  BUFX2 U3579 ( .A(n8790), .Y(n3028) );
  BUFX2 U3580 ( .A(n8842), .Y(n3029) );
  BUFX2 U3581 ( .A(n8905), .Y(n3030) );
  BUFX2 U3582 ( .A(n9024), .Y(n3031) );
  BUFX2 U3583 ( .A(n9082), .Y(n3032) );
  BUFX2 U3584 ( .A(n9133), .Y(n3033) );
  BUFX2 U3585 ( .A(n9157), .Y(n3034) );
  BUFX2 U3586 ( .A(n9356), .Y(n3035) );
  BUFX2 U3587 ( .A(n9420), .Y(n3036) );
  BUFX2 U3588 ( .A(n9585), .Y(n3037) );
  BUFX2 U3589 ( .A(n9678), .Y(n3038) );
  BUFX2 U3590 ( .A(n9824), .Y(n3039) );
  BUFX2 U3591 ( .A(n9878), .Y(n3040) );
  BUFX2 U3592 ( .A(n9944), .Y(n3041) );
  BUFX2 U3593 ( .A(n10059), .Y(n3042) );
  BUFX2 U3594 ( .A(n10173), .Y(n3043) );
  BUFX2 U3595 ( .A(n10197), .Y(n3044) );
  BUFX2 U3596 ( .A(n10338), .Y(n3045) );
  BUFX2 U3597 ( .A(n10408), .Y(n3046) );
  INVX1 U3598 ( .A(n10475), .Y(n3047) );
  INVX1 U3599 ( .A(n3047), .Y(n3048) );
  BUFX2 U3600 ( .A(n10483), .Y(n3049) );
  BUFX2 U3601 ( .A(n10533), .Y(n3050) );
  BUFX2 U3602 ( .A(n10571), .Y(n3051) );
  BUFX2 U3603 ( .A(n7348), .Y(n3052) );
  BUFX2 U3604 ( .A(n7443), .Y(n3053) );
  BUFX2 U3605 ( .A(n8365), .Y(n3054) );
  BUFX2 U3606 ( .A(n8687), .Y(n3055) );
  BUFX2 U3607 ( .A(n9374), .Y(n3056) );
  BUFX2 U3608 ( .A(n9519), .Y(n3057) );
  BUFX2 U3609 ( .A(n10427), .Y(n3058) );
  BUFX2 U3610 ( .A(n10493), .Y(n3059) );
  BUFX2 U3611 ( .A(n10514), .Y(n3060) );
  AND2X1 U3612 ( .A(n5918), .B(n6066), .Y(n6560) );
  INVX1 U3613 ( .A(n6560), .Y(n3061) );
  AND2X1 U3614 ( .A(n6858), .B(n6721), .Y(n6586) );
  INVX1 U3615 ( .A(n6586), .Y(n3062) );
  INVX1 U3616 ( .A(n6609), .Y(n3063) );
  AND2X1 U3617 ( .A(n1099), .B(n5826), .Y(n6594) );
  INVX1 U3618 ( .A(n6594), .Y(n3064) );
  AND2X1 U3619 ( .A(n2552), .B(n6102), .Y(n6597) );
  INVX1 U3620 ( .A(n6597), .Y(n3065) );
  INVX1 U3621 ( .A(n6638), .Y(n3066) );
  AND2X1 U3622 ( .A(n8968), .B(n6939), .Y(n6653) );
  INVX1 U3623 ( .A(n6653), .Y(n3067) );
  AND2X1 U3624 ( .A(n5903), .B(n7171), .Y(n6664) );
  INVX1 U3625 ( .A(n6664), .Y(n3068) );
  INVX1 U3626 ( .A(n6687), .Y(n3069) );
  AND2X1 U3627 ( .A(n1100), .B(n6127), .Y(n6671) );
  INVX1 U3628 ( .A(n6671), .Y(n3070) );
  INVX1 U3629 ( .A(n6674), .Y(n3071) );
  AND2X1 U3630 ( .A(n6315), .B(n10502), .Y(n6679) );
  INVX1 U3631 ( .A(n6679), .Y(n3072) );
  AND2X1 U3632 ( .A(n2556), .B(n6102), .Y(n6839) );
  INVX1 U3633 ( .A(n6839), .Y(n3073) );
  INVX1 U3634 ( .A(n6874), .Y(n3074) );
  AND2X1 U3635 ( .A(n10500), .B(n4699), .Y(n7095) );
  INVX1 U3636 ( .A(n7095), .Y(n3075) );
  AND2X1 U3637 ( .A(n7022), .B(n4849), .Y(n7098) );
  INVX1 U3638 ( .A(n7098), .Y(n3076) );
  INVX1 U3639 ( .A(n7121), .Y(n3077) );
  INVX1 U3640 ( .A(n7106), .Y(n3078) );
  INVX1 U3641 ( .A(n7109), .Y(n3079) );
  AND2X1 U3642 ( .A(n6627), .B(n4860), .Y(n7165) );
  INVX1 U3643 ( .A(n7165), .Y(n3080) );
  INVX1 U3644 ( .A(n7168), .Y(n3081) );
  AND2X1 U3645 ( .A(n7172), .B(n7417), .Y(n7174) );
  INVX1 U3646 ( .A(n7174), .Y(n3082) );
  INVX1 U3647 ( .A(n7196), .Y(n3083) );
  AND2X1 U3648 ( .A(n1108), .B(n5826), .Y(n7181) );
  INVX1 U3649 ( .A(n7181), .Y(n3084) );
  AND2X1 U3650 ( .A(n2561), .B(n5831), .Y(n7184) );
  INVX1 U3651 ( .A(n7184), .Y(n3085) );
  AND2X1 U3652 ( .A(n5764), .B(n7284), .Y(n7226) );
  INVX1 U3653 ( .A(n7226), .Y(n3086) );
  AND2X1 U3654 ( .A(n2563), .B(n5831), .Y(n7292) );
  INVX1 U3655 ( .A(n7292), .Y(n3087) );
  INVX1 U3656 ( .A(n7324), .Y(n3088) );
  AND2X1 U3657 ( .A(n7222), .B(n7353), .Y(n7356) );
  INVX1 U3658 ( .A(n7356), .Y(n3089) );
  AND2X1 U3659 ( .A(n7361), .B(n7138), .Y(n7365) );
  INVX1 U3660 ( .A(n7365), .Y(n3090) );
  INVX1 U3661 ( .A(n7389), .Y(n3091) );
  AND2X1 U3662 ( .A(n1111), .B(n5826), .Y(n7374) );
  INVX1 U3663 ( .A(n7374), .Y(n3092) );
  AND2X1 U3664 ( .A(n2564), .B(n6102), .Y(n7377) );
  INVX1 U3665 ( .A(n7377), .Y(n3093) );
  AND2X1 U3666 ( .A(n2565), .B(n5831), .Y(n7439) );
  INVX1 U3667 ( .A(n7439), .Y(n3094) );
  AND2X1 U3668 ( .A(n414), .B(n6117), .Y(n7447) );
  INVX1 U3669 ( .A(n7447), .Y(n3095) );
  AND2X1 U3670 ( .A(n1803), .B(n5777), .Y(n7451) );
  INVX1 U3671 ( .A(n7451), .Y(n3096) );
  AND2X1 U3672 ( .A(n1321), .B(n5785), .Y(n7455) );
  INVX1 U3673 ( .A(n7455), .Y(n3097) );
  AND2X1 U3674 ( .A(n5958), .B(n6066), .Y(n7593) );
  INVX1 U3675 ( .A(n7593), .Y(n3098) );
  AND2X1 U3676 ( .A(n7877), .B(n6721), .Y(n7618) );
  INVX1 U3677 ( .A(n7618), .Y(n3099) );
  INVX1 U3678 ( .A(n7640), .Y(n3100) );
  AND2X1 U3679 ( .A(n1115), .B(n5826), .Y(n7625) );
  INVX1 U3680 ( .A(n7625), .Y(n3101) );
  AND2X1 U3681 ( .A(n2568), .B(n6102), .Y(n7628) );
  INVX1 U3682 ( .A(n7628), .Y(n3102) );
  INVX1 U3683 ( .A(n7666), .Y(n3103) );
  AND2X1 U3684 ( .A(n8968), .B(n7926), .Y(n7681) );
  INVX1 U3685 ( .A(n7681), .Y(n3104) );
  AND2X1 U3686 ( .A(n6191), .B(n8167), .Y(n7693) );
  INVX1 U3687 ( .A(n7693), .Y(n3105) );
  INVX1 U3688 ( .A(n7715), .Y(n3106) );
  AND2X1 U3689 ( .A(n1116), .B(n5826), .Y(n7700) );
  INVX1 U3690 ( .A(n7700), .Y(n3107) );
  AND2X1 U3691 ( .A(n2569), .B(n5831), .Y(n7703) );
  INVX1 U3692 ( .A(n7703), .Y(n3108) );
  AND2X2 U3693 ( .A(n3181), .B(n5776), .Y(n7790) );
  INVX1 U3694 ( .A(n7790), .Y(n3109) );
  AND2X2 U3695 ( .A(n3182), .B(n5776), .Y(n7841) );
  INVX1 U3696 ( .A(n7841), .Y(n3110) );
  AND2X1 U3697 ( .A(n2572), .B(n5831), .Y(n7856) );
  INVX1 U3698 ( .A(n7856), .Y(n3111) );
  INVX1 U3699 ( .A(n7893), .Y(n3112) );
  AND2X2 U3700 ( .A(n3183), .B(n5776), .Y(n7906) );
  INVX1 U3701 ( .A(n7906), .Y(n3113) );
  AND2X1 U3702 ( .A(n5957), .B(n9500), .Y(n7909) );
  INVX1 U3703 ( .A(n7909), .Y(n3114) );
  AND2X1 U3704 ( .A(n6791), .B(n7926), .Y(n7928) );
  INVX1 U3705 ( .A(n7928), .Y(n3115) );
  AND2X1 U3706 ( .A(n7873), .B(n7931), .Y(n7935) );
  INVX1 U3707 ( .A(n7935), .Y(n3116) );
  AND2X2 U3708 ( .A(n3184), .B(n5776), .Y(n7969) );
  INVX1 U3709 ( .A(n7969), .Y(n3117) );
  AND2X2 U3710 ( .A(n3186), .B(n5776), .Y(n8077) );
  INVX1 U3711 ( .A(n8077), .Y(n3118) );
  AND2X1 U3712 ( .A(n6347), .B(n10502), .Y(n8080) );
  INVX1 U3713 ( .A(n8080), .Y(n3119) );
  AND2X1 U3714 ( .A(n1123), .B(n5826), .Y(n8090) );
  INVX1 U3715 ( .A(n8090), .Y(n3120) );
  AND2X1 U3716 ( .A(n2576), .B(n5831), .Y(n8093) );
  INVX1 U3717 ( .A(n8093), .Y(n3121) );
  INVX1 U3718 ( .A(n8139), .Y(n3122) );
  AND2X2 U3719 ( .A(n3187), .B(n5776), .Y(n8152) );
  INVX1 U3720 ( .A(n8152), .Y(n3123) );
  AND2X1 U3721 ( .A(n6203), .B(n6299), .Y(n8164) );
  INVX1 U3722 ( .A(n8164), .Y(n3124) );
  AND2X1 U3723 ( .A(n8415), .B(n6626), .Y(n8191) );
  INVX1 U3724 ( .A(n8191), .Y(n3125) );
  INVX1 U3725 ( .A(n8213), .Y(n3126) );
  AND2X1 U3726 ( .A(n1124), .B(n5826), .Y(n8198) );
  INVX1 U3727 ( .A(n8198), .Y(n3127) );
  AND2X1 U3728 ( .A(n2577), .B(n5831), .Y(n8201) );
  INVX1 U3729 ( .A(n8201), .Y(n3128) );
  AND2X2 U3730 ( .A(n3188), .B(n5776), .Y(n8226) );
  INVX1 U3731 ( .A(n8226), .Y(n3257) );
  AND2X2 U3732 ( .A(n3189), .B(n5776), .Y(n8290) );
  INVX1 U3733 ( .A(n8290), .Y(n3258) );
  AND2X1 U3734 ( .A(n1046), .B(n6129), .Y(n8295) );
  INVX1 U3735 ( .A(n8295), .Y(n3259) );
  AND2X1 U3736 ( .A(n1126), .B(n5826), .Y(n8305) );
  INVX1 U3737 ( .A(n8305), .Y(n3260) );
  AND2X1 U3738 ( .A(n2579), .B(n5831), .Y(n8308) );
  INVX1 U3739 ( .A(n8308), .Y(n3261) );
  INVX1 U3740 ( .A(n8340), .Y(n3262) );
  AND2X2 U3741 ( .A(n3190), .B(n5776), .Y(n8353) );
  INVX1 U3742 ( .A(n8353), .Y(n3263) );
  AND2X1 U3743 ( .A(n7222), .B(n8369), .Y(n8372) );
  INVX1 U3744 ( .A(n8372), .Y(n3264) );
  AND2X1 U3745 ( .A(n8377), .B(n8156), .Y(n8381) );
  INVX1 U3746 ( .A(n8381), .Y(n3265) );
  INVX1 U3747 ( .A(n8403), .Y(n3266) );
  AND2X1 U3748 ( .A(n1127), .B(n5826), .Y(n8388) );
  INVX1 U3749 ( .A(n8388), .Y(n3267) );
  AND2X1 U3750 ( .A(n2580), .B(n5831), .Y(n8391) );
  INVX1 U3751 ( .A(n8391), .Y(n3268) );
  AND2X1 U3752 ( .A(n8485), .B(n8418), .Y(n8421) );
  INVX1 U3753 ( .A(n8421), .Y(n3269) );
  AND2X1 U3754 ( .A(n6296), .B(n9969), .Y(n8438) );
  INVX1 U3755 ( .A(n8438), .Y(n3270) );
  AND2X1 U3756 ( .A(n582), .B(n5823), .Y(n8441) );
  INVX1 U3757 ( .A(n8441), .Y(n3271) );
  AND2X1 U3758 ( .A(n1129), .B(n5826), .Y(n8513) );
  INVX1 U3759 ( .A(n8513), .Y(n3272) );
  AND2X1 U3760 ( .A(n1324), .B(n6139), .Y(n8581) );
  INVX1 U3761 ( .A(n8581), .Y(n3273) );
  AND2X1 U3762 ( .A(n6315), .B(n6066), .Y(n8595) );
  INVX1 U3763 ( .A(n8595), .Y(n3274) );
  AND2X1 U3764 ( .A(n8883), .B(n6721), .Y(n8620) );
  INVX1 U3765 ( .A(n8620), .Y(n3275) );
  INVX1 U3766 ( .A(n8642), .Y(n3276) );
  AND2X1 U3767 ( .A(n1067), .B(n5826), .Y(n8627) );
  INVX1 U3768 ( .A(n8627), .Y(n3277) );
  AND2X1 U3769 ( .A(n2584), .B(n5831), .Y(n8630) );
  INVX1 U3770 ( .A(n8630), .Y(n3278) );
  AND2X1 U3771 ( .A(n1071), .B(n6127), .Y(n8861) );
  INVX1 U3772 ( .A(n8861), .Y(n3279) );
  AND2X1 U3773 ( .A(n2588), .B(n5831), .Y(n8864) );
  INVX1 U3774 ( .A(n8864), .Y(n3280) );
  INVX1 U3775 ( .A(n8899), .Y(n3281) );
  AND2X1 U3776 ( .A(n5934), .B(n10502), .Y(n9092) );
  INVX1 U3777 ( .A(n9092), .Y(n3282) );
  AND2X1 U3778 ( .A(n1075), .B(n6127), .Y(n9102) );
  INVX1 U3779 ( .A(n9102), .Y(n3283) );
  AND2X1 U3780 ( .A(n2592), .B(n5831), .Y(n9105) );
  INVX1 U3781 ( .A(n9105), .Y(n3284) );
  INVX1 U3782 ( .A(n9151), .Y(n3285) );
  INVX1 U3783 ( .A(n9176), .Y(n3286) );
  AND2X1 U3784 ( .A(n152), .B(n6626), .Y(n9202) );
  INVX1 U3785 ( .A(n9202), .Y(n3287) );
  INVX1 U3786 ( .A(n9225), .Y(n3288) );
  AND2X1 U3787 ( .A(n1076), .B(n6127), .Y(n9209) );
  INVX1 U3788 ( .A(n9209), .Y(n3289) );
  AND2X1 U3789 ( .A(n2593), .B(n5831), .Y(n9212) );
  INVX1 U3790 ( .A(n9212), .Y(n3290) );
  AND2X1 U3791 ( .A(n2595), .B(n6102), .Y(n9318) );
  INVX1 U3792 ( .A(n9318), .Y(n3291) );
  INVX1 U3793 ( .A(n9350), .Y(n3292) );
  AND2X1 U3794 ( .A(n7222), .B(n9379), .Y(n9382) );
  INVX1 U3795 ( .A(n9382), .Y(n3293) );
  AND2X1 U3796 ( .A(n9387), .B(n9168), .Y(n9391) );
  INVX1 U3797 ( .A(n9391), .Y(n3294) );
  INVX1 U3798 ( .A(n9414), .Y(n3295) );
  AND2X1 U3799 ( .A(n1079), .B(n6127), .Y(n9398) );
  INVX1 U3800 ( .A(n9398), .Y(n3296) );
  AND2X1 U3801 ( .A(n2596), .B(n5831), .Y(n9401) );
  INVX1 U3802 ( .A(n9401), .Y(n3297) );
  AND2X1 U3803 ( .A(n1771), .B(n5777), .Y(n9471) );
  INVX1 U3804 ( .A(n9471), .Y(n3298) );
  AND2X1 U3805 ( .A(n920), .B(n5824), .Y(n9523) );
  INVX1 U3806 ( .A(n9523), .Y(n3299) );
  AND2X1 U3807 ( .A(n1081), .B(n5826), .Y(n9527) );
  INVX1 U3808 ( .A(n9527), .Y(n3300) );
  AND2X1 U3809 ( .A(n6029), .B(n6066), .Y(n9621) );
  INVX1 U3810 ( .A(n9621), .Y(n3301) );
  AND2X1 U3811 ( .A(n9922), .B(n6721), .Y(n9650) );
  INVX1 U3812 ( .A(n9650), .Y(n3302) );
  INVX1 U3813 ( .A(n9672), .Y(n3303) );
  AND2X1 U3814 ( .A(n1083), .B(n6127), .Y(n9657) );
  INVX1 U3815 ( .A(n9657), .Y(n3304) );
  AND2X1 U3816 ( .A(n2600), .B(n5831), .Y(n9660) );
  INVX1 U3817 ( .A(n9660), .Y(n3305) );
  INVX1 U3818 ( .A(n9698), .Y(n3306) );
  AND2X1 U3819 ( .A(n8968), .B(n9972), .Y(n9714) );
  INVX1 U3820 ( .A(n9714), .Y(n3307) );
  INVX1 U3821 ( .A(n9727), .Y(n3308) );
  INVX1 U3822 ( .A(n9750), .Y(n3309) );
  AND2X1 U3823 ( .A(n1084), .B(n6127), .Y(n9735) );
  INVX1 U3824 ( .A(n9735), .Y(n3310) );
  AND2X1 U3825 ( .A(n2601), .B(n5831), .Y(n9738) );
  INVX1 U3826 ( .A(n9738), .Y(n3311) );
  AND2X2 U3827 ( .A(n3149), .B(n5776), .Y(n9831) );
  INVX1 U3828 ( .A(n9831), .Y(n3312) );
  AND2X2 U3829 ( .A(n3150), .B(n5776), .Y(n9885) );
  INVX1 U3830 ( .A(n9885), .Y(n3313) );
  AND2X1 U3831 ( .A(n2604), .B(n5831), .Y(n9900) );
  INVX1 U3832 ( .A(n9900), .Y(n3314) );
  INVX1 U3833 ( .A(n9938), .Y(n3315) );
  AND2X2 U3834 ( .A(n3151), .B(n5776), .Y(n9951) );
  INVX1 U3835 ( .A(n9951), .Y(n3316) );
  AND2X1 U3836 ( .A(n9500), .B(n6342), .Y(n9954) );
  INVX1 U3837 ( .A(n9954), .Y(n3317) );
  AND2X1 U3838 ( .A(n6791), .B(n9972), .Y(n9974) );
  INVX1 U3839 ( .A(n9974), .Y(n3318) );
  AND2X1 U3840 ( .A(n9725), .B(n9918), .Y(n9981) );
  INVX1 U3841 ( .A(n9981), .Y(n3319) );
  AND2X2 U3842 ( .A(n3152), .B(n5776), .Y(n10015) );
  INVX1 U3843 ( .A(n10015), .Y(n3320) );
  AND2X2 U3844 ( .A(n3154), .B(n5776), .Y(n10129) );
  INVX1 U3845 ( .A(n10129), .Y(n3321) );
  AND2X1 U3846 ( .A(n5976), .B(n10502), .Y(n10132) );
  INVX1 U3847 ( .A(n10132), .Y(n3322) );
  AND2X1 U3848 ( .A(n2608), .B(n5831), .Y(n10145) );
  INVX1 U3849 ( .A(n10145), .Y(n3323) );
  INVX1 U3850 ( .A(n10191), .Y(n3324) );
  AND2X2 U3851 ( .A(n3155), .B(n5776), .Y(n10204) );
  INVX1 U3852 ( .A(n10204), .Y(n3325) );
  AND2X1 U3853 ( .A(n153), .B(n6626), .Y(n10242) );
  INVX1 U3854 ( .A(n10242), .Y(n3326) );
  INVX1 U3855 ( .A(n10265), .Y(n3327) );
  AND2X1 U3856 ( .A(n1092), .B(n6127), .Y(n10249) );
  INVX1 U3857 ( .A(n10249), .Y(n3328) );
  AND2X1 U3858 ( .A(n2609), .B(n6102), .Y(n10252) );
  INVX1 U3859 ( .A(n10252), .Y(n3330) );
  AND2X2 U3860 ( .A(n3156), .B(n5776), .Y(n10278) );
  INVX1 U3861 ( .A(n10278), .Y(n3331) );
  AND2X2 U3862 ( .A(n3157), .B(n5776), .Y(n10345) );
  INVX1 U3863 ( .A(n10345), .Y(n3332) );
  AND2X1 U3864 ( .A(n1014), .B(n5786), .Y(n10350) );
  INVX1 U3865 ( .A(n10350), .Y(n3333) );
  AND2X1 U3866 ( .A(n1094), .B(n6127), .Y(n10360) );
  INVX1 U3867 ( .A(n10360), .Y(n3334) );
  AND2X1 U3868 ( .A(n2611), .B(n5831), .Y(n10363) );
  INVX1 U3869 ( .A(n10363), .Y(n3335) );
  INVX1 U3870 ( .A(n10402), .Y(n3336) );
  AND2X2 U3871 ( .A(n3158), .B(n5776), .Y(n10415) );
  INVX1 U3872 ( .A(n10415), .Y(n3338) );
  AND2X1 U3873 ( .A(n7222), .B(n10431), .Y(n10434) );
  INVX1 U3874 ( .A(n10434), .Y(n3339) );
  AND2X1 U3875 ( .A(n10439), .B(n10208), .Y(n10443) );
  INVX1 U3876 ( .A(n10443), .Y(n3340) );
  INVX1 U3877 ( .A(n10469), .Y(n3341) );
  AND2X1 U3878 ( .A(n1095), .B(n6127), .Y(n10452) );
  AND2X1 U3879 ( .A(n2612), .B(n6102), .Y(n10455) );
  INVX1 U3880 ( .A(n10455), .Y(n3342) );
  AND2X1 U3881 ( .A(oprA[34]), .B(n10502), .Y(n10460) );
  INVX1 U3882 ( .A(n10460), .Y(n3343) );
  AND2X1 U3883 ( .A(n614), .B(n5823), .Y(n10545) );
  INVX1 U3884 ( .A(n10545), .Y(n3344) );
  AND2X1 U3885 ( .A(n6054), .B(n5175), .Y(n10524) );
  INVX1 U3886 ( .A(n10524), .Y(n3346) );
  INVX1 U3887 ( .A(n10529), .Y(n3347) );
  AND2X1 U3888 ( .A(n687), .B(n5790), .Y(n10537) );
  INVX1 U3889 ( .A(n10537), .Y(n3348) );
  AND2X1 U3890 ( .A(n1096), .B(n6127), .Y(n10541) );
  INVX1 U3891 ( .A(n10541), .Y(n3349) );
  AND2X1 U3892 ( .A(n2293), .B(n5838), .Y(n10592) );
  INVX1 U3893 ( .A(n10592), .Y(n3350) );
  AND2X1 U3894 ( .A(n688), .B(n5790), .Y(n10596) );
  INVX1 U3895 ( .A(n10596), .Y(n3351) );
  BUFX2 U3896 ( .A(n6577), .Y(n3352) );
  BUFX2 U3897 ( .A(n7609), .Y(n3354) );
  BUFX2 U3898 ( .A(n8614), .Y(n3355) );
  BUFX2 U3899 ( .A(n9643), .Y(n3356) );
  BUFX2 U3900 ( .A(n6548), .Y(n3357) );
  BUFX2 U3901 ( .A(n6726), .Y(n3358) );
  BUFX2 U3902 ( .A(n7243), .Y(n3359) );
  BUFX2 U3903 ( .A(n7583), .Y(n3360) );
  BUFX2 U3904 ( .A(n7751), .Y(n3362) );
  BUFX2 U3905 ( .A(n8257), .Y(n3363) );
  BUFX2 U3906 ( .A(n8585), .Y(n3364) );
  BUFX2 U3907 ( .A(n8758), .Y(n3365) );
  BUFX2 U3908 ( .A(n9268), .Y(n3366) );
  BUFX2 U3909 ( .A(n9611), .Y(n3367) );
  BUFX2 U3910 ( .A(n9787), .Y(n3368) );
  BUFX2 U3911 ( .A(n10310), .Y(n3370) );
  INVX1 U3912 ( .A(n7139), .Y(n3371) );
  BUFX2 U3913 ( .A(n8161), .Y(n3372) );
  BUFX2 U3914 ( .A(n8241), .Y(n3373) );
  BUFX2 U3915 ( .A(n9173), .Y(n3374) );
  BUFX2 U3916 ( .A(n9252), .Y(n3375) );
  BUFX2 U3917 ( .A(n10213), .Y(n3376) );
  BUFX2 U3918 ( .A(n10294), .Y(n3378) );
  BUFX2 U3919 ( .A(n6559), .Y(n3379) );
  BUFX2 U3920 ( .A(n6585), .Y(n3380) );
  BUFX2 U3921 ( .A(n6593), .Y(n3381) );
  BUFX2 U3922 ( .A(n6596), .Y(n3382) );
  BUFX2 U3923 ( .A(n6637), .Y(n3383) );
  BUFX2 U3924 ( .A(n6652), .Y(n3384) );
  BUFX2 U3925 ( .A(n6663), .Y(n3386) );
  BUFX2 U3926 ( .A(n6670), .Y(n3387) );
  BUFX2 U3927 ( .A(n6673), .Y(n3388) );
  BUFX2 U3928 ( .A(n6803), .Y(n3389) );
  BUFX2 U3929 ( .A(n6835), .Y(n3390) );
  BUFX2 U3930 ( .A(n6838), .Y(n3391) );
  BUFX2 U3931 ( .A(n7094), .Y(n3392) );
  BUFX2 U3932 ( .A(n7097), .Y(n3393) );
  BUFX2 U3933 ( .A(n7108), .Y(n3394) );
  BUFX2 U3934 ( .A(n7164), .Y(n3395) );
  BUFX2 U3935 ( .A(n7173), .Y(n3396) );
  BUFX2 U3936 ( .A(n7180), .Y(n3397) );
  BUFX2 U3937 ( .A(n7183), .Y(n3398) );
  BUFX2 U3938 ( .A(n7240), .Y(n3399) );
  BUFX2 U3939 ( .A(n7291), .Y(n3400) );
  BUFX2 U3940 ( .A(n7342), .Y(n3401) );
  BUFX2 U3941 ( .A(n7347), .Y(n3402) );
  BUFX2 U3942 ( .A(n7355), .Y(n3403) );
  BUFX2 U3943 ( .A(n7364), .Y(n3404) );
  BUFX2 U3944 ( .A(n7373), .Y(n3405) );
  BUFX2 U3945 ( .A(n7376), .Y(n3406) );
  BUFX2 U3946 ( .A(n7438), .Y(n3407) );
  BUFX2 U3947 ( .A(n7454), .Y(n3408) );
  BUFX2 U3948 ( .A(n7592), .Y(n3409) );
  BUFX2 U3949 ( .A(n7617), .Y(n3410) );
  BUFX2 U3950 ( .A(n7624), .Y(n3411) );
  BUFX2 U3951 ( .A(n7627), .Y(n3412) );
  BUFX2 U3952 ( .A(n7665), .Y(n3413) );
  BUFX2 U3953 ( .A(n7680), .Y(n3414) );
  BUFX2 U3954 ( .A(n7692), .Y(n3415) );
  BUFX2 U3955 ( .A(n7699), .Y(n3416) );
  BUFX2 U3956 ( .A(n7702), .Y(n3417) );
  BUFX2 U3957 ( .A(n7845), .Y(n3418) );
  BUFX2 U3958 ( .A(n7852), .Y(n3419) );
  BUFX2 U3959 ( .A(n7855), .Y(n3420) );
  BUFX2 U3960 ( .A(n7908), .Y(n3421) );
  BUFX2 U3961 ( .A(n7927), .Y(n3422) );
  BUFX2 U3962 ( .A(n7934), .Y(n3423) );
  BUFX2 U3963 ( .A(n8079), .Y(n3424) );
  BUFX2 U3964 ( .A(n8089), .Y(n3425) );
  BUFX2 U3965 ( .A(n8092), .Y(n3426) );
  BUFX2 U3966 ( .A(n8159), .Y(n3427) );
  BUFX2 U3967 ( .A(n8190), .Y(n3428) );
  BUFX2 U3968 ( .A(n8197), .Y(n3429) );
  BUFX2 U3969 ( .A(n8200), .Y(n3430) );
  BUFX2 U3970 ( .A(n8254), .Y(n3431) );
  BUFX2 U3971 ( .A(n8294), .Y(n3432) );
  BUFX2 U3972 ( .A(n8304), .Y(n3433) );
  BUFX2 U3973 ( .A(n8307), .Y(n3434) );
  BUFX2 U3974 ( .A(n8315), .Y(n3435) );
  BUFX2 U3975 ( .A(n8358), .Y(n3436) );
  BUFX2 U3976 ( .A(n8364), .Y(n3437) );
  BUFX2 U3977 ( .A(n8371), .Y(n3438) );
  BUFX2 U3978 ( .A(n8380), .Y(n3439) );
  BUFX2 U3979 ( .A(n8387), .Y(n3440) );
  BUFX2 U3980 ( .A(n8390), .Y(n3441) );
  BUFX2 U3981 ( .A(n8420), .Y(n3442) );
  BUFX2 U3982 ( .A(n8437), .Y(n3443) );
  BUFX2 U3983 ( .A(n8440), .Y(n3444) );
  BUFX2 U3984 ( .A(n8580), .Y(n3445) );
  BUFX2 U3985 ( .A(n8594), .Y(n3446) );
  BUFX2 U3986 ( .A(n8619), .Y(n3447) );
  BUFX2 U3987 ( .A(n8626), .Y(n3448) );
  BUFX2 U3988 ( .A(n8629), .Y(n3449) );
  BUFX2 U3989 ( .A(n8686), .Y(n3578) );
  BUFX2 U3990 ( .A(n8853), .Y(n3579) );
  BUFX2 U3991 ( .A(n8860), .Y(n3580) );
  BUFX2 U3992 ( .A(n9091), .Y(n3581) );
  BUFX2 U3993 ( .A(n9101), .Y(n3582) );
  BUFX2 U3994 ( .A(n9104), .Y(n3583) );
  BUFX2 U3995 ( .A(n9171), .Y(n3584) );
  BUFX2 U3996 ( .A(n9201), .Y(n3585) );
  BUFX2 U3997 ( .A(n9208), .Y(n3586) );
  BUFX2 U3998 ( .A(n9211), .Y(n3587) );
  BUFX2 U3999 ( .A(n9265), .Y(n3588) );
  BUFX2 U4000 ( .A(n9317), .Y(n3589) );
  BUFX2 U4001 ( .A(n9325), .Y(n3590) );
  BUFX2 U4002 ( .A(n9368), .Y(n3591) );
  BUFX2 U4003 ( .A(n9373), .Y(n3592) );
  BUFX2 U4004 ( .A(n9381), .Y(n3593) );
  BUFX2 U4005 ( .A(n9390), .Y(n3594) );
  BUFX2 U4006 ( .A(n9397), .Y(n3595) );
  INVX1 U4007 ( .A(n9400), .Y(n3596) );
  INVX1 U4008 ( .A(n3596), .Y(n3597) );
  BUFX2 U4009 ( .A(n9518), .Y(n3598) );
  BUFX2 U4010 ( .A(n9620), .Y(n3599) );
  BUFX2 U4011 ( .A(n9649), .Y(n3600) );
  BUFX2 U4012 ( .A(n9656), .Y(n3601) );
  BUFX2 U4013 ( .A(n9659), .Y(n3602) );
  BUFX2 U4014 ( .A(n9697), .Y(n3603) );
  BUFX2 U4015 ( .A(n9713), .Y(n3604) );
  BUFX2 U4016 ( .A(n9726), .Y(n3605) );
  BUFX2 U4017 ( .A(n9734), .Y(n3606) );
  BUFX2 U4018 ( .A(n9737), .Y(n3607) );
  BUFX2 U4019 ( .A(n9889), .Y(n3608) );
  BUFX2 U4020 ( .A(n9899), .Y(n3609) );
  BUFX2 U4021 ( .A(n9953), .Y(n3610) );
  BUFX2 U4022 ( .A(n9956), .Y(n3611) );
  BUFX2 U4023 ( .A(n9973), .Y(n3612) );
  BUFX2 U4024 ( .A(n9980), .Y(n3613) );
  BUFX2 U4025 ( .A(n10131), .Y(n3614) );
  BUFX2 U4026 ( .A(n10144), .Y(n3615) );
  BUFX2 U4027 ( .A(n10211), .Y(n3616) );
  BUFX2 U4028 ( .A(n10241), .Y(n3617) );
  BUFX2 U4029 ( .A(n10248), .Y(n3618) );
  BUFX2 U4030 ( .A(n10251), .Y(n3619) );
  BUFX2 U4031 ( .A(n10307), .Y(n3620) );
  BUFX2 U4032 ( .A(n10349), .Y(n3621) );
  BUFX2 U4033 ( .A(n10359), .Y(n3622) );
  BUFX2 U4034 ( .A(n10362), .Y(n3623) );
  BUFX2 U4035 ( .A(n10420), .Y(n3624) );
  BUFX2 U4036 ( .A(n10426), .Y(n3625) );
  BUFX2 U4037 ( .A(n10433), .Y(n3626) );
  BUFX2 U4038 ( .A(n10442), .Y(n3627) );
  BUFX2 U4039 ( .A(n10454), .Y(n3628) );
  INVX1 U4040 ( .A(n10459), .Y(n3629) );
  INVX1 U4041 ( .A(n3629), .Y(n3630) );
  BUFX2 U4042 ( .A(n10523), .Y(n3631) );
  BUFX2 U4043 ( .A(n10540), .Y(n3632) );
  BUFX2 U4044 ( .A(n10570), .Y(n3633) );
  BUFX2 U4045 ( .A(n6547), .Y(n3634) );
  BUFX2 U4046 ( .A(n6614), .Y(n3635) );
  BUFX2 U4047 ( .A(n7043), .Y(n3636) );
  BUFX2 U4048 ( .A(n7105), .Y(n3637) );
  BUFX2 U4049 ( .A(n7489), .Y(n3638) );
  INVX1 U4050 ( .A(n30), .Y(n3639) );
  BUFX2 U4051 ( .A(n7582), .Y(n3640) );
  BUFX2 U4052 ( .A(n8056), .Y(n3641) );
  BUFX2 U4053 ( .A(n8473), .Y(n3642) );
  BUFX2 U4054 ( .A(n8512), .Y(n3643) );
  BUFX2 U4055 ( .A(n8584), .Y(n3644) );
  BUFX2 U4056 ( .A(n8647), .Y(n3645) );
  BUFX2 U4057 ( .A(n9067), .Y(n3646) );
  BUFX2 U4058 ( .A(n9610), .Y(n3647) );
  BUFX2 U4059 ( .A(n10107), .Y(n3648) );
  BUFX2 U4060 ( .A(n10482), .Y(n3649) );
  OR2X1 U4061 ( .A(n6519), .B(n6518), .Y(n6520) );
  INVX1 U4062 ( .A(n6520), .Y(n3650) );
  AND2X1 U4063 ( .A(n9), .B(n6281), .Y(n6550) );
  INVX1 U4064 ( .A(n6550), .Y(n3651) );
  AND2X1 U4065 ( .A(n5887), .B(n6281), .Y(n6571) );
  INVX1 U4066 ( .A(n6571), .Y(n3652) );
  OR2X1 U4067 ( .A(n6630), .B(n6781), .Y(n6631) );
  INVX1 U4068 ( .A(n6631), .Y(n3653) );
  OR2X1 U4069 ( .A(n6724), .B(n5807), .Y(n6725) );
  INVX1 U4070 ( .A(n6725), .Y(n3654) );
  AND2X1 U4071 ( .A(n6971), .B(n5833), .Y(n6972) );
  INVX1 U4072 ( .A(n6972), .Y(n3655) );
  AND2X1 U4073 ( .A(n6169), .B(n6291), .Y(n7067) );
  INVX1 U4074 ( .A(n7067), .Y(n3656) );
  AND2X1 U4075 ( .A(n566), .B(n5823), .Y(n7442) );
  INVX1 U4076 ( .A(n7442), .Y(n3657) );
  AND2X1 U4077 ( .A(n735), .B(n6119), .Y(n7446) );
  INVX1 U4078 ( .A(n7446), .Y(n3658) );
  OR2X1 U4079 ( .A(n7552), .B(n7551), .Y(n7553) );
  INVX1 U4080 ( .A(n7553), .Y(n3659) );
  INVX1 U4081 ( .A(n7585), .Y(n3660) );
  AND2X1 U4082 ( .A(n5886), .B(n5967), .Y(n7603) );
  INVX1 U4083 ( .A(n7603), .Y(n3661) );
  OR2X1 U4084 ( .A(n7659), .B(n7803), .Y(n7660) );
  INVX1 U4085 ( .A(n7660), .Y(n3662) );
  OR2X1 U4086 ( .A(n7749), .B(n5810), .Y(n7750) );
  INVX1 U4087 ( .A(n7750), .Y(n3663) );
  AND2X1 U4088 ( .A(n6201), .B(n6310), .Y(n8104) );
  INVX1 U4089 ( .A(n8104), .Y(n3664) );
  AND2X1 U4090 ( .A(n1049), .B(n6129), .Y(n8508) );
  INVX1 U4091 ( .A(n8508), .Y(n3665) );
  OR2X1 U4092 ( .A(n8556), .B(n8555), .Y(n8557) );
  INVX1 U4093 ( .A(n8557), .Y(n3666) );
  INVX1 U4094 ( .A(n8587), .Y(n3667) );
  AND2X1 U4095 ( .A(n5887), .B(n6324), .Y(n8605) );
  INVX1 U4096 ( .A(n8605), .Y(n3668) );
  OR2X1 U4097 ( .A(n8701), .B(n8810), .Y(n8702) );
  INVX1 U4098 ( .A(n8702), .Y(n3669) );
  OR2X1 U4099 ( .A(n8756), .B(n5809), .Y(n8757) );
  INVX1 U4100 ( .A(n8757), .Y(n3670) );
  INVX1 U4101 ( .A(n9116), .Y(n3671) );
  AND2X1 U4102 ( .A(n3240), .B(n5827), .Y(n9514) );
  INVX1 U4103 ( .A(n9514), .Y(n3672) );
  AND2X1 U4104 ( .A(n383), .B(n5778), .Y(n9522) );
  INVX1 U4105 ( .A(n9522), .Y(n3673) );
  AND2X1 U4106 ( .A(n1772), .B(n6121), .Y(n9526) );
  INVX1 U4107 ( .A(n9526), .Y(n3674) );
  AND2X1 U4108 ( .A(n455), .B(n5839), .Y(n9530) );
  INVX1 U4109 ( .A(n9530), .Y(n3675) );
  OR2X1 U4110 ( .A(n9579), .B(n9578), .Y(n9580) );
  INVX1 U4111 ( .A(n9580), .Y(n3676) );
  INVX1 U4112 ( .A(n9613), .Y(n3677) );
  INVX1 U4113 ( .A(n9634), .Y(n3678) );
  OR2X1 U4114 ( .A(n9692), .B(n9844), .Y(n9693) );
  INVX1 U4115 ( .A(n9693), .Y(n3679) );
  OR2X1 U4116 ( .A(n9785), .B(n5811), .Y(n9786) );
  INVX1 U4117 ( .A(n9786), .Y(n3680) );
  INVX1 U4118 ( .A(n10156), .Y(n3681) );
  AND2X1 U4119 ( .A(n5865), .B(n10491), .Y(n10492) );
  INVX1 U4120 ( .A(n10492), .Y(n3682) );
  INVX1 U4121 ( .A(n10528), .Y(n3683) );
  AND2X1 U4122 ( .A(n2292), .B(n5838), .Y(n10532) );
  INVX1 U4123 ( .A(n10532), .Y(n3684) );
  AND2X1 U4124 ( .A(n1755), .B(n5777), .Y(n10536) );
  INVX1 U4125 ( .A(n10536), .Y(n3685) );
  AND2X1 U4126 ( .A(n518), .B(n6143), .Y(n10548) );
  INVX1 U4127 ( .A(n10548), .Y(n3686) );
  INVX1 U4128 ( .A(n10591), .Y(n3687) );
  AND2X1 U4129 ( .A(n1756), .B(n5777), .Y(n10595) );
  INVX1 U4130 ( .A(n10595), .Y(n3688) );
  INVX1 U4131 ( .A(n6493), .Y(n3690) );
  INVX1 U4132 ( .A(n6494), .Y(n3691) );
  INVX1 U4133 ( .A(n6495), .Y(n3692) );
  INVX1 U4134 ( .A(n6524), .Y(n3695) );
  INVX1 U4135 ( .A(n6525), .Y(n3696) );
  INVX1 U4136 ( .A(n6526), .Y(n3697) );
  INVX1 U4137 ( .A(n6715), .Y(n3700) );
  INVX1 U4138 ( .A(n6716), .Y(n3701) );
  INVX1 U4139 ( .A(n6745), .Y(n3704) );
  INVX1 U4140 ( .A(n6746), .Y(n3705) );
  INVX1 U4141 ( .A(n6747), .Y(n3706) );
  INVX1 U4142 ( .A(n6772), .Y(n3709) );
  INVX1 U4143 ( .A(n6773), .Y(n3710) );
  INVX1 U4144 ( .A(n6774), .Y(n3711) );
  BUFX2 U4145 ( .A(n6810), .Y(n3713) );
  INVX1 U4146 ( .A(n6861), .Y(n3715) );
  INVX1 U4147 ( .A(n6862), .Y(n3716) );
  INVX1 U4148 ( .A(n6863), .Y(n3717) );
  INVX1 U4149 ( .A(n6886), .Y(n3720) );
  INVX1 U4150 ( .A(n6888), .Y(n3721) );
  BUFX2 U4151 ( .A(n6908), .Y(n3723) );
  INVX1 U4152 ( .A(n6958), .Y(n3725) );
  INVX1 U4153 ( .A(n6959), .Y(n3726) );
  INVX1 U4154 ( .A(n6960), .Y(n3727) );
  INVX1 U4155 ( .A(n6982), .Y(n3730) );
  INVX1 U4156 ( .A(n6983), .Y(n3731) );
  INVX1 U4157 ( .A(n6984), .Y(n3732) );
  INVX1 U4158 ( .A(n7019), .Y(n3735) );
  INVX1 U4159 ( .A(n7020), .Y(n3736) );
  INVX1 U4160 ( .A(n7021), .Y(n3737) );
  INVX1 U4161 ( .A(n7038), .Y(n3740) );
  INVX1 U4162 ( .A(n7039), .Y(n3741) );
  INVX1 U4163 ( .A(n7040), .Y(n3742) );
  INVX1 U4164 ( .A(n7077), .Y(n3745) );
  INVX1 U4165 ( .A(n7079), .Y(n3746) );
  INVX1 U4166 ( .A(n7143), .Y(n3749) );
  INVX1 U4167 ( .A(n7145), .Y(n3750) );
  INVX1 U4168 ( .A(n7218), .Y(n3753) );
  INVX1 U4169 ( .A(n7219), .Y(n3754) );
  INVX1 U4170 ( .A(n7220), .Y(n3755) );
  BUFX2 U4171 ( .A(n7261), .Y(n3757) );
  INVX1 U4172 ( .A(n7313), .Y(n3759) );
  INVX1 U4173 ( .A(n7314), .Y(n3760) );
  INVX1 U4174 ( .A(n7315), .Y(n3761) );
  INVX1 U4175 ( .A(n7410), .Y(n3764) );
  INVX1 U4176 ( .A(n7411), .Y(n3765) );
  INVX1 U4177 ( .A(n7412), .Y(n3766) );
  INVX1 U4178 ( .A(n7472), .Y(n3769) );
  INVX1 U4179 ( .A(n7473), .Y(n3770) );
  INVX1 U4180 ( .A(n7474), .Y(n3899) );
  INVX1 U4181 ( .A(n7534), .Y(n3903) );
  INVX1 U4182 ( .A(n7535), .Y(n3904) );
  INVX1 U4183 ( .A(n7536), .Y(n3905) );
  INVX1 U4184 ( .A(n7557), .Y(n3908) );
  INVX1 U4185 ( .A(n7558), .Y(n3909) );
  INVX1 U4186 ( .A(n7559), .Y(n3910) );
  INVX1 U4187 ( .A(n7742), .Y(n3913) );
  INVX1 U4188 ( .A(n7743), .Y(n3914) );
  BUFX2 U4189 ( .A(n7776), .Y(n3916) );
  INVX1 U4190 ( .A(n7794), .Y(n3918) );
  INVX1 U4191 ( .A(n7795), .Y(n3919) );
  INVX1 U4192 ( .A(n7796), .Y(n3920) );
  INVX1 U4193 ( .A(n7817), .Y(n3923) );
  INVX1 U4194 ( .A(n7818), .Y(n3924) );
  INVX1 U4195 ( .A(n7819), .Y(n3925) );
  INVX1 U4196 ( .A(n7880), .Y(n3928) );
  INVX1 U4197 ( .A(n7881), .Y(n3929) );
  INVX1 U4198 ( .A(n7882), .Y(n3930) );
  INVX1 U4199 ( .A(n7916), .Y(n3933) );
  INVX1 U4200 ( .A(n7918), .Y(n3934) );
  INVX1 U4201 ( .A(n7974), .Y(n3937) );
  INVX1 U4202 ( .A(n7975), .Y(n3938) );
  INVX1 U4203 ( .A(n7976), .Y(n3939) );
  INVX1 U4204 ( .A(n7996), .Y(n3942) );
  INVX1 U4205 ( .A(n7997), .Y(n3943) );
  INVX1 U4206 ( .A(n7998), .Y(n3944) );
  INVX1 U4207 ( .A(n8032), .Y(n3947) );
  INVX1 U4208 ( .A(n8033), .Y(n3948) );
  INVX1 U4209 ( .A(n8034), .Y(n3949) );
  INVX1 U4210 ( .A(n8051), .Y(n3952) );
  INVX1 U4211 ( .A(n8052), .Y(n3953) );
  INVX1 U4212 ( .A(n8053), .Y(n3954) );
  BUFX2 U4213 ( .A(n8137), .Y(n3956) );
  INVX1 U4214 ( .A(n8168), .Y(n3958) );
  INVX1 U4215 ( .A(n8170), .Y(n3959) );
  INVX1 U4216 ( .A(n8235), .Y(n3962) );
  INVX1 U4217 ( .A(n8236), .Y(n3963) );
  INVX1 U4218 ( .A(n8237), .Y(n3964) );
  BUFX2 U4219 ( .A(n8276), .Y(n3966) );
  INVX1 U4220 ( .A(n8329), .Y(n3968) );
  INVX1 U4221 ( .A(n8330), .Y(n3969) );
  INVX1 U4222 ( .A(n8331), .Y(n3970) );
  INVX1 U4223 ( .A(n8479), .Y(n3973) );
  INVX1 U4224 ( .A(n8480), .Y(n3974) );
  INVX1 U4225 ( .A(n8481), .Y(n3975) );
  INVX1 U4226 ( .A(n8493), .Y(n3978) );
  INVX1 U4227 ( .A(n8494), .Y(n3979) );
  INVX1 U4228 ( .A(n8495), .Y(n3980) );
  INVX1 U4229 ( .A(n8538), .Y(n3983) );
  INVX1 U4230 ( .A(n8539), .Y(n3984) );
  INVX1 U4231 ( .A(n8540), .Y(n3985) );
  INVX1 U4232 ( .A(n8561), .Y(n3988) );
  INVX1 U4233 ( .A(n8562), .Y(n3989) );
  INVX1 U4234 ( .A(n8563), .Y(n3990) );
  INVX1 U4235 ( .A(n8654), .Y(n3993) );
  INVX1 U4236 ( .A(n8656), .Y(n3994) );
  BUFX2 U4237 ( .A(n8676), .Y(n3996) );
  INVX1 U4238 ( .A(n8749), .Y(n3998) );
  INVX1 U4239 ( .A(n8750), .Y(n3999) );
  BUFX2 U4240 ( .A(n8783), .Y(n4001) );
  INVX1 U4241 ( .A(n8801), .Y(n4003) );
  INVX1 U4242 ( .A(n8802), .Y(n4004) );
  INVX1 U4243 ( .A(n8803), .Y(n4005) );
  BUFX2 U4244 ( .A(n8835), .Y(n4007) );
  INVX1 U4245 ( .A(n8886), .Y(n4009) );
  INVX1 U4246 ( .A(n8887), .Y(n4010) );
  INVX1 U4247 ( .A(n8888), .Y(n4011) );
  INVX1 U4248 ( .A(n8912), .Y(n4014) );
  INVX1 U4249 ( .A(n8914), .Y(n4015) );
  BUFX2 U4250 ( .A(n8934), .Y(n4017) );
  INVX1 U4251 ( .A(n8986), .Y(n4019) );
  INVX1 U4252 ( .A(n8987), .Y(n4020) );
  INVX1 U4253 ( .A(n8988), .Y(n4021) );
  INVX1 U4254 ( .A(n9007), .Y(n4024) );
  INVX1 U4255 ( .A(n9008), .Y(n4025) );
  INVX1 U4256 ( .A(n9009), .Y(n4026) );
  INVX1 U4257 ( .A(n9043), .Y(n4029) );
  INVX1 U4258 ( .A(n9044), .Y(n4030) );
  INVX1 U4259 ( .A(n9045), .Y(n4031) );
  BUFX2 U4260 ( .A(n9075), .Y(n4033) );
  BUFX2 U4261 ( .A(n9149), .Y(n4034) );
  INVX1 U4262 ( .A(n9180), .Y(n4036) );
  INVX1 U4263 ( .A(n9182), .Y(n4037) );
  INVX1 U4264 ( .A(n9247), .Y(n4040) );
  INVX1 U4265 ( .A(n9248), .Y(n4041) );
  INVX1 U4266 ( .A(n9249), .Y(n4042) );
  INVX1 U4267 ( .A(n9278), .Y(n4045) );
  INVX1 U4268 ( .A(n9279), .Y(n4046) );
  INVX1 U4269 ( .A(n9280), .Y(n4047) );
  INVX1 U4270 ( .A(n9339), .Y(n4050) );
  INVX1 U4271 ( .A(n9340), .Y(n4051) );
  INVX1 U4272 ( .A(n9341), .Y(n4052) );
  INVX1 U4273 ( .A(n9438), .Y(n4056) );
  INVX1 U4274 ( .A(n9440), .Y(n4057) );
  INVX1 U4275 ( .A(n9493), .Y(n4060) );
  INVX1 U4276 ( .A(n9495), .Y(n4061) );
  INVX1 U4277 ( .A(n9561), .Y(n4064) );
  INVX1 U4278 ( .A(n9562), .Y(n4065) );
  INVX1 U4279 ( .A(n9563), .Y(n4066) );
  BUFX2 U4280 ( .A(n9593), .Y(n4068) );
  INVX1 U4281 ( .A(n5488), .Y(n4070) );
  INVX1 U4282 ( .A(n9779), .Y(n4071) );
  BUFX2 U4283 ( .A(n9817), .Y(n4073) );
  INVX1 U4284 ( .A(n9835), .Y(n4075) );
  INVX1 U4285 ( .A(n9836), .Y(n4076) );
  INVX1 U4286 ( .A(n9837), .Y(n4077) );
  BUFX2 U4287 ( .A(n9871), .Y(n4079) );
  INVX1 U4288 ( .A(n9925), .Y(n4081) );
  INVX1 U4289 ( .A(n9926), .Y(n4082) );
  INVX1 U4290 ( .A(n9927), .Y(n4083) );
  INVX1 U4291 ( .A(n9961), .Y(n4086) );
  INVX1 U4292 ( .A(n9963), .Y(n4087) );
  INVX1 U4293 ( .A(n10020), .Y(n4090) );
  INVX1 U4294 ( .A(n10021), .Y(n4091) );
  INVX1 U4295 ( .A(n10022), .Y(n4092) );
  INVX1 U4296 ( .A(n10042), .Y(n4095) );
  INVX1 U4297 ( .A(n10043), .Y(n4096) );
  INVX1 U4298 ( .A(n10044), .Y(n4097) );
  INVX1 U4299 ( .A(n10079), .Y(n4100) );
  INVX1 U4300 ( .A(n10080), .Y(n4101) );
  INVX1 U4301 ( .A(n10081), .Y(n4102) );
  BUFX2 U4302 ( .A(n10115), .Y(n4104) );
  BUFX2 U4303 ( .A(n10189), .Y(n4105) );
  INVX1 U4304 ( .A(n10219), .Y(n4107) );
  INVX1 U4305 ( .A(n10221), .Y(n4108) );
  INVX1 U4306 ( .A(n10287), .Y(n4111) );
  INVX1 U4307 ( .A(n10288), .Y(n4112) );
  INVX1 U4308 ( .A(n10289), .Y(n4113) );
  BUFX2 U4309 ( .A(n10331), .Y(n4115) );
  INVX1 U4310 ( .A(n10391), .Y(n4117) );
  INVX1 U4311 ( .A(n10392), .Y(n4118) );
  INVX1 U4312 ( .A(n10393), .Y(n4119) );
  INVX1 U4313 ( .A(n6946), .Y(n4121) );
  OR2X1 U4314 ( .A(n4713), .B(n4715), .Y(n8110) );
  INVX1 U4315 ( .A(n8110), .Y(n4122) );
  INVX1 U4316 ( .A(n8726), .Y(n4123) );
  INVX1 U4317 ( .A(n8974), .Y(n4124) );
  OR2X1 U4318 ( .A(n5632), .B(n5565), .Y(n9122) );
  INVX1 U4319 ( .A(n9122), .Y(n4125) );
  INVX1 U4320 ( .A(n9482), .Y(n4126) );
  OR2X1 U4321 ( .A(n4714), .B(n4716), .Y(n10162) );
  INVX1 U4322 ( .A(n10162), .Y(n4127) );
  BUFX2 U4323 ( .A(n6684), .Y(n4128) );
  BUFX2 U4324 ( .A(n6809), .Y(n4129) );
  BUFX2 U4325 ( .A(n6945), .Y(n4130) );
  INVX1 U4326 ( .A(n6988), .Y(n4132) );
  INVX1 U4327 ( .A(n6990), .Y(n4133) );
  INVX1 U4328 ( .A(n7045), .Y(n4136) );
  INVX1 U4329 ( .A(n7047), .Y(n4137) );
  INVX1 U4330 ( .A(n7113), .Y(n4140) );
  INVX1 U4331 ( .A(n5342), .Y(n4141) );
  INVX1 U4332 ( .A(n7188), .Y(n4144) );
  INVX1 U4333 ( .A(n7190), .Y(n4145) );
  INVX1 U4334 ( .A(n7255), .Y(n4148) );
  INVX1 U4335 ( .A(n7257), .Y(n4149) );
  INVX1 U4336 ( .A(n7381), .Y(n4152) );
  INVX1 U4337 ( .A(n7383), .Y(n4153) );
  INVX1 U4338 ( .A(n7707), .Y(n4156) );
  INVX1 U4339 ( .A(n7709), .Y(n4157) );
  INVX1 U4340 ( .A(n7822), .Y(n4160) );
  INVX1 U4341 ( .A(n7824), .Y(n4161) );
  INVX1 U4342 ( .A(n7947), .Y(n4164) );
  INVX1 U4343 ( .A(n7949), .Y(n4165) );
  INVX1 U4344 ( .A(n8001), .Y(n4168) );
  INVX1 U4345 ( .A(n8003), .Y(n4169) );
  INVX1 U4346 ( .A(n8058), .Y(n4172) );
  INVX1 U4347 ( .A(n8060), .Y(n4173) );
  INVX1 U4348 ( .A(n8395), .Y(n4176) );
  INVX1 U4349 ( .A(n8397), .Y(n4177) );
  INVX1 U4350 ( .A(n8712), .Y(n4180) );
  INVX1 U4351 ( .A(n8714), .Y(n4181) );
  INVX1 U4352 ( .A(n8829), .Y(n4184) );
  INVX1 U4353 ( .A(n8831), .Y(n4185) );
  BUFX2 U4354 ( .A(n8973), .Y(n4187) );
  INVX1 U4355 ( .A(n9012), .Y(n4189) );
  INVX1 U4356 ( .A(n9014), .Y(n4190) );
  INVX1 U4357 ( .A(n9069), .Y(n4193) );
  INVX1 U4358 ( .A(n9071), .Y(n4194) );
  INVX1 U4359 ( .A(n9405), .Y(n4197) );
  INVX1 U4360 ( .A(n9407), .Y(n4198) );
  INVX1 U4361 ( .A(n9445), .Y(n4201) );
  INVX1 U4362 ( .A(n9447), .Y(n4202) );
  INVX1 U4363 ( .A(n9742), .Y(n4205) );
  INVX1 U4364 ( .A(n9744), .Y(n4206) );
  INVX1 U4365 ( .A(n9865), .Y(n4209) );
  INVX1 U4366 ( .A(n9867), .Y(n4210) );
  INVX1 U4367 ( .A(n9993), .Y(n4213) );
  INVX1 U4368 ( .A(n9995), .Y(n4214) );
  INVX1 U4369 ( .A(n10047), .Y(n4217) );
  INVX1 U4370 ( .A(n10049), .Y(n4218) );
  INVX1 U4371 ( .A(n10109), .Y(n4221) );
  INVX1 U4372 ( .A(n10111), .Y(n4222) );
  INVX1 U4373 ( .A(n6514), .Y(n4224) );
  INVX1 U4374 ( .A(n6532), .Y(n4225) );
  INVX1 U4375 ( .A(n6606), .Y(n4226) );
  INVX1 U4376 ( .A(n6739), .Y(n4227) );
  INVX1 U4377 ( .A(n6754), .Y(n4228) );
  INVX1 U4378 ( .A(n6795), .Y(n4229) );
  INVX1 U4379 ( .A(n6872), .Y(n4230) );
  INVX1 U4380 ( .A(n6894), .Y(n4231) );
  INVX1 U4381 ( .A(n6907), .Y(n4232) );
  INVX1 U4382 ( .A(n6979), .Y(n4233) );
  INVX1 U4383 ( .A(n7035), .Y(n4234) );
  INVX1 U4384 ( .A(n7247), .Y(n4235) );
  INVX1 U4385 ( .A(n7322), .Y(n4236) );
  INVX1 U4386 ( .A(n7502), .Y(n4237) );
  INVX1 U4387 ( .A(n7548), .Y(n4238) );
  INVX1 U4388 ( .A(n7565), .Y(n4239) );
  INVX1 U4389 ( .A(n7637), .Y(n4240) );
  INVX1 U4390 ( .A(n7761), .Y(n4241) );
  INVX1 U4391 ( .A(n7775), .Y(n4242) );
  INVX1 U4392 ( .A(n7814), .Y(n4243) );
  INVX1 U4393 ( .A(n7891), .Y(n4244) );
  INVX1 U4394 ( .A(n7925), .Y(n4245) );
  INVX1 U4395 ( .A(n7993), .Y(n4246) );
  INVX1 U4396 ( .A(n8048), .Y(n4247) );
  INVX1 U4397 ( .A(n8136), .Y(n4248) );
  INVX1 U4398 ( .A(n8210), .Y(n4249) );
  INVX1 U4399 ( .A(n8261), .Y(n4250) );
  INVX1 U4400 ( .A(n8275), .Y(n4251) );
  INVX1 U4401 ( .A(n8338), .Y(n4252) );
  INVX1 U4402 ( .A(n8431), .Y(n4253) );
  INVX1 U4403 ( .A(n8452), .Y(n4254) );
  INVX1 U4404 ( .A(n8507), .Y(n4255) );
  INVX1 U4405 ( .A(n8552), .Y(n4256) );
  INVX1 U4406 ( .A(n8569), .Y(n4257) );
  INVX1 U4407 ( .A(n8639), .Y(n4258) );
  INVX1 U4408 ( .A(n8662), .Y(n4259) );
  INVX1 U4409 ( .A(n8675), .Y(n4260) );
  INVX1 U4410 ( .A(n8768), .Y(n4261) );
  INVX1 U4411 ( .A(n8782), .Y(n4262) );
  INVX1 U4412 ( .A(n8821), .Y(n4263) );
  INVX1 U4413 ( .A(n8897), .Y(n4264) );
  INVX1 U4414 ( .A(n8920), .Y(n4265) );
  INVX1 U4415 ( .A(n8933), .Y(n4266) );
  INVX1 U4416 ( .A(n9004), .Y(n4267) );
  INVX1 U4417 ( .A(n9059), .Y(n4268) );
  INVX1 U4418 ( .A(n9148), .Y(n4269) );
  INVX1 U4419 ( .A(n9222), .Y(n4270) );
  INVX1 U4420 ( .A(n9272), .Y(n4271) );
  INVX1 U4421 ( .A(n9286), .Y(n4272) );
  INVX1 U4422 ( .A(n9348), .Y(n4273) );
  AND2X1 U4423 ( .A(n5691), .B(n5600), .Y(n9434) );
  INVX1 U4424 ( .A(n9434), .Y(n4274) );
  INVX1 U4425 ( .A(n9575), .Y(n4275) );
  INVX1 U4426 ( .A(n9592), .Y(n4276) );
  INVX1 U4427 ( .A(n9669), .Y(n4277) );
  INVX1 U4428 ( .A(n9801), .Y(n4278) );
  INVX1 U4429 ( .A(n9816), .Y(n4279) );
  INVX1 U4430 ( .A(n9857), .Y(n4280) );
  INVX1 U4431 ( .A(n9936), .Y(n4281) );
  INVX1 U4432 ( .A(n9971), .Y(n4282) );
  INVX1 U4433 ( .A(n10039), .Y(n4283) );
  INVX1 U4434 ( .A(n10098), .Y(n4284) );
  INVX1 U4435 ( .A(n10188), .Y(n4289) );
  INVX1 U4436 ( .A(n10262), .Y(n4290) );
  INVX1 U4437 ( .A(n10314), .Y(n4291) );
  INVX1 U4438 ( .A(n10330), .Y(n4292) );
  INVX1 U4439 ( .A(n10400), .Y(n4293) );
  OR2X1 U4440 ( .A(n10499), .B(n5721), .Y(n10511) );
  INVX1 U4441 ( .A(n10511), .Y(n4294) );
  INVX1 U4442 ( .A(n6603), .Y(n4296) );
  INVX1 U4443 ( .A(n6605), .Y(n4297) );
  INVX1 U4444 ( .A(n6681), .Y(n4300) );
  INVX1 U4445 ( .A(n6683), .Y(n4304) );
  INVX1 U4446 ( .A(n6736), .Y(n4307) );
  INVX1 U4447 ( .A(n6738), .Y(n4308) );
  BUFX2 U4448 ( .A(n6753), .Y(n4310) );
  INVX1 U4449 ( .A(n6793), .Y(n4312) );
  INVX1 U4450 ( .A(n6869), .Y(n4315) );
  INVX1 U4451 ( .A(n6871), .Y(n4319) );
  INVX1 U4452 ( .A(n6942), .Y(n4322) );
  INVX1 U4453 ( .A(n6943), .Y(n4323) );
  INVX1 U4454 ( .A(n6944), .Y(n4324) );
  INVX1 U4455 ( .A(n6977), .Y(n4327) );
  INVX1 U4456 ( .A(n7032), .Y(n4330) );
  INVX1 U4457 ( .A(n7034), .Y(n4334) );
  INVX1 U4458 ( .A(n7116), .Y(n4337) );
  INVX1 U4459 ( .A(n7118), .Y(n4338) );
  INVX1 U4460 ( .A(n7154), .Y(n4341) );
  INVX1 U4461 ( .A(n7191), .Y(n4344) );
  INVX1 U4462 ( .A(n7193), .Y(n4345) );
  INVX1 U4463 ( .A(n7244), .Y(n4378) );
  INVX1 U4464 ( .A(n7246), .Y(n4379) );
  INVX1 U4465 ( .A(n7319), .Y(n4382) );
  INVX1 U4466 ( .A(n7321), .Y(n4383) );
  INVX1 U4467 ( .A(n7384), .Y(n4386) );
  INVX1 U4468 ( .A(n7386), .Y(n4387) );
  INVX1 U4469 ( .A(n7434), .Y(n4390) );
  INVX1 U4470 ( .A(n7435), .Y(n4391) );
  INVX1 U4471 ( .A(n7436), .Y(n4392) );
  INVX1 U4472 ( .A(n7634), .Y(n4395) );
  INVX1 U4473 ( .A(n7636), .Y(n4396) );
  INVX1 U4474 ( .A(n7710), .Y(n4399) );
  INVX1 U4475 ( .A(n7712), .Y(n4400) );
  INVX1 U4476 ( .A(n7758), .Y(n4403) );
  INVX1 U4477 ( .A(n7760), .Y(n4404) );
  INVX1 U4478 ( .A(n7772), .Y(n4407) );
  INVX1 U4479 ( .A(n7774), .Y(n4408) );
  INVX1 U4480 ( .A(n7812), .Y(n4411) );
  INVX1 U4481 ( .A(n7888), .Y(n4414) );
  INVX1 U4482 ( .A(n7890), .Y(n4415) );
  INVX1 U4483 ( .A(n7952), .Y(n4418) );
  INVX1 U4484 ( .A(n7953), .Y(n4419) );
  INVX1 U4485 ( .A(n7991), .Y(n4422) );
  INVX1 U4486 ( .A(n8045), .Y(n4425) );
  INVX1 U4487 ( .A(n8047), .Y(n4426) );
  INVX1 U4488 ( .A(n8133), .Y(n4429) );
  INVX1 U4489 ( .A(n8135), .Y(n4430) );
  INVX1 U4490 ( .A(n8178), .Y(n4433) );
  INVX1 U4491 ( .A(n8207), .Y(n4436) );
  INVX1 U4492 ( .A(n8209), .Y(n4437) );
  INVX1 U4493 ( .A(n8258), .Y(n4440) );
  INVX1 U4494 ( .A(n8260), .Y(n4441) );
  INVX1 U4495 ( .A(n8272), .Y(n4444) );
  INVX1 U4496 ( .A(n8274), .Y(n4445) );
  INVX1 U4497 ( .A(n8335), .Y(n4448) );
  INVX1 U4498 ( .A(n8337), .Y(n4449) );
  INVX1 U4499 ( .A(n8398), .Y(n4452) );
  INVX1 U4500 ( .A(n8400), .Y(n4453) );
  INVX1 U4501 ( .A(n8429), .Y(n4456) );
  INVX1 U4502 ( .A(n8430), .Y(n4457) );
  BUFX2 U4503 ( .A(n8451), .Y(n4459) );
  INVX1 U4504 ( .A(n5433), .Y(n4461) );
  INVX1 U4505 ( .A(n8638), .Y(n4462) );
  INVX1 U4506 ( .A(n8723), .Y(n4465) );
  INVX1 U4507 ( .A(n8724), .Y(n4466) );
  INVX1 U4508 ( .A(n8725), .Y(n4467) );
  INVX1 U4509 ( .A(n8765), .Y(n4470) );
  INVX1 U4510 ( .A(n8767), .Y(n4471) );
  INVX1 U4511 ( .A(n8779), .Y(n4474) );
  INVX1 U4512 ( .A(n8781), .Y(n4475) );
  INVX1 U4513 ( .A(n8819), .Y(n4478) );
  INVX1 U4514 ( .A(n8894), .Y(n4481) );
  INVX1 U4515 ( .A(n8896), .Y(n4482) );
  INVX1 U4516 ( .A(n8970), .Y(n4485) );
  INVX1 U4517 ( .A(n8971), .Y(n4486) );
  INVX1 U4518 ( .A(n8972), .Y(n4487) );
  INVX1 U4519 ( .A(n9002), .Y(n4490) );
  INVX1 U4520 ( .A(n9056), .Y(n4493) );
  INVX1 U4521 ( .A(n9058), .Y(n4494) );
  INVX1 U4522 ( .A(n9145), .Y(n4497) );
  INVX1 U4523 ( .A(n9147), .Y(n4498) );
  INVX1 U4524 ( .A(n9189), .Y(n4501) );
  BUFX2 U4525 ( .A(n9221), .Y(n4503) );
  INVX1 U4526 ( .A(n9269), .Y(n4505) );
  INVX1 U4527 ( .A(n9271), .Y(n4506) );
  INVX1 U4528 ( .A(n9283), .Y(n4509) );
  INVX1 U4529 ( .A(n9285), .Y(n4510) );
  INVX1 U4530 ( .A(n9345), .Y(n4513) );
  INVX1 U4531 ( .A(n9347), .Y(n4514) );
  INVX1 U4532 ( .A(n9478), .Y(n4518) );
  INVX1 U4533 ( .A(n9479), .Y(n4519) );
  INVX1 U4534 ( .A(n9480), .Y(n4520) );
  INVX1 U4535 ( .A(n9505), .Y(n4523) );
  INVX1 U4536 ( .A(n9506), .Y(n4524) );
  INVX1 U4537 ( .A(n9666), .Y(n4527) );
  INVX1 U4538 ( .A(n9668), .Y(n4528) );
  INVX1 U4539 ( .A(n9745), .Y(n4531) );
  INVX1 U4540 ( .A(n9747), .Y(n4532) );
  INVX1 U4541 ( .A(n9798), .Y(n4535) );
  INVX1 U4542 ( .A(n9800), .Y(n4536) );
  INVX1 U4543 ( .A(n9813), .Y(n4539) );
  INVX1 U4544 ( .A(n9815), .Y(n4540) );
  INVX1 U4545 ( .A(n9855), .Y(n4543) );
  INVX1 U4546 ( .A(n9933), .Y(n4546) );
  INVX1 U4547 ( .A(n9935), .Y(n4547) );
  INVX1 U4548 ( .A(n9998), .Y(n4550) );
  INVX1 U4549 ( .A(n9999), .Y(n4551) );
  INVX1 U4550 ( .A(n10037), .Y(n4554) );
  INVX1 U4551 ( .A(n10095), .Y(n4557) );
  INVX1 U4552 ( .A(n10097), .Y(n4558) );
  INVX1 U4553 ( .A(n10185), .Y(n4561) );
  INVX1 U4554 ( .A(n10187), .Y(n4562) );
  INVX1 U4555 ( .A(n10228), .Y(n4565) );
  BUFX2 U4556 ( .A(n10261), .Y(n4567) );
  INVX1 U4557 ( .A(n10311), .Y(n4569) );
  INVX1 U4558 ( .A(n10313), .Y(n4570) );
  INVX1 U4559 ( .A(n10397), .Y(n4574) );
  INVX1 U4560 ( .A(n10399), .Y(n4575) );
  INVX1 U4561 ( .A(n10508), .Y(n4579) );
  INVX1 U4562 ( .A(n10510), .Y(n4580) );
  INVX1 U4563 ( .A(n10576), .Y(n4583) );
  INVX1 U4564 ( .A(n10578), .Y(n4584) );
  INVX1 U4565 ( .A(n6513), .Y(n4586) );
  INVX1 U4566 ( .A(n6531), .Y(n4587) );
  INVX1 U4567 ( .A(n6808), .Y(n4588) );
  INVX1 U4568 ( .A(n6893), .Y(n4589) );
  INVX1 U4569 ( .A(n6906), .Y(n4590) );
  AND2X1 U4570 ( .A(n5487), .B(n5423), .Y(n6993) );
  INVX1 U4571 ( .A(n6993), .Y(n4591) );
  INVX1 U4572 ( .A(n7050), .Y(n4592) );
  INVX1 U4573 ( .A(n7260), .Y(n4593) );
  INVX1 U4574 ( .A(n7481), .Y(n4594) );
  INVX1 U4575 ( .A(n7501), .Y(n4595) );
  INVX1 U4576 ( .A(n7547), .Y(n4596) );
  INVX1 U4577 ( .A(n7564), .Y(n4597) );
  INVX1 U4578 ( .A(n7827), .Y(n4598) );
  INVX1 U4579 ( .A(n8006), .Y(n4599) );
  INVX1 U4580 ( .A(n8063), .Y(n4600) );
  INVX1 U4581 ( .A(n8489), .Y(n4601) );
  INVX1 U4582 ( .A(n8506), .Y(n4602) );
  INVX1 U4583 ( .A(n8551), .Y(n4603) );
  INVX1 U4584 ( .A(n8568), .Y(n4604) );
  INVX1 U4585 ( .A(n8661), .Y(n4605) );
  INVX1 U4586 ( .A(n8674), .Y(n4606) );
  INVX1 U4587 ( .A(n8834), .Y(n4607) );
  INVX1 U4588 ( .A(n8919), .Y(n4608) );
  INVX1 U4589 ( .A(n8932), .Y(n4609) );
  INVX1 U4590 ( .A(n9017), .Y(n4610) );
  INVX1 U4591 ( .A(n9074), .Y(n4611) );
  INVX1 U4592 ( .A(n9433), .Y(n4612) );
  INVX1 U4593 ( .A(n9450), .Y(n4613) );
  INVX1 U4594 ( .A(n9574), .Y(n4614) );
  INVX1 U4595 ( .A(n9591), .Y(n4615) );
  INVX1 U4596 ( .A(n9870), .Y(n4616) );
  INVX1 U4597 ( .A(n10052), .Y(n4617) );
  INVX1 U4598 ( .A(n10114), .Y(n4618) );
  AND2X1 U4599 ( .A(n6517), .B(n5931), .Y(n7013) );
  AND2X1 U4600 ( .A(n5932), .B(n9688), .Y(n7009) );
  AND2X1 U4601 ( .A(n6277), .B(n9632), .Y(n6910) );
  AND2X1 U4602 ( .A(n6279), .B(n6081), .Y(n7011) );
  AND2X1 U4603 ( .A(n6579), .B(n6273), .Y(n6720) );
  AND2X1 U4604 ( .A(n10291), .B(n6160), .Y(n6854) );
  AND2X1 U4605 ( .A(n6517), .B(n5933), .Y(n7092) );
  AND2X1 U4606 ( .A(n6517), .B(n5918), .Y(n6630) );
  AND2X1 U4607 ( .A(n6579), .B(n6275), .Y(n6781) );
  AND2X1 U4608 ( .A(n5820), .B(n5932), .Y(n7161) );
  AND2X1 U4609 ( .A(n6282), .B(n6083), .Y(n6962) );
  AND2X1 U4610 ( .A(n5820), .B(n5934), .Y(n7213) );
  AND2X1 U4611 ( .A(n6517), .B(n6282), .Y(n6708) );
  AND2X1 U4612 ( .A(n6579), .B(n5932), .Y(n7093) );
  AND2X1 U4613 ( .A(n6517), .B(n6275), .Y(n6724) );
  AND2X1 U4614 ( .A(n7070), .B(n5937), .Y(n7230) );
  AND2X1 U4615 ( .A(n7550), .B(n5974), .Y(n8026) );
  AND2X1 U4616 ( .A(n5973), .B(n9688), .Y(n8022) );
  AND2X1 U4617 ( .A(n5966), .B(n9632), .Y(n7940) );
  AND2X1 U4618 ( .A(n6296), .B(n6081), .Y(n8024) );
  AND2X1 U4619 ( .A(n7611), .B(n5958), .Y(n7747) );
  AND2X1 U4620 ( .A(n10291), .B(n6190), .Y(n7872) );
  AND2X1 U4621 ( .A(n7550), .B(n5975), .Y(n8125) );
  AND2X1 U4622 ( .A(n7550), .B(n5958), .Y(n7659) );
  AND2X1 U4623 ( .A(n7611), .B(n5961), .Y(n7803) );
  AND2X1 U4624 ( .A(n7662), .B(n6188), .Y(n7691) );
  AND2X1 U4625 ( .A(n5767), .B(n5974), .Y(n8182) );
  AND2X1 U4626 ( .A(n6297), .B(n9688), .Y(n7978) );
  AND2X1 U4627 ( .A(n5767), .B(n5975), .Y(n8230) );
  AND2X1 U4628 ( .A(n7550), .B(n6297), .Y(n7735) );
  AND2X1 U4629 ( .A(n7611), .B(n5973), .Y(n8126) );
  AND2X1 U4630 ( .A(n7550), .B(n5961), .Y(n7749) );
  AND2X1 U4631 ( .A(n8102), .B(n6301), .Y(n8244) );
  AND2X1 U4632 ( .A(n8554), .B(n6328), .Y(n9037) );
  AND2X1 U4633 ( .A(n6328), .B(n9688), .Y(n9033) );
  AND2X1 U4634 ( .A(n6322), .B(n9626), .Y(n9035) );
  AND2X1 U4635 ( .A(n10291), .B(n6219), .Y(n8879) );
  AND2X1 U4636 ( .A(n8554), .B(n6330), .Y(n9137) );
  AND2X1 U4637 ( .A(n8610), .B(n5276), .Y(n8810) );
  AND2X1 U4638 ( .A(n5768), .B(n6328), .Y(n9193) );
  AND2X1 U4639 ( .A(n6325), .B(n9688), .Y(n8990) );
  AND2X1 U4640 ( .A(n5768), .B(n6330), .Y(n9242) );
  AND2X1 U4641 ( .A(n8554), .B(n6325), .Y(n8742) );
  AND2X1 U4642 ( .A(n8610), .B(n6328), .Y(n9138) );
  AND2X1 U4643 ( .A(n8554), .B(n5276), .Y(n8756) );
  AND2X1 U4644 ( .A(n9114), .B(n6008), .Y(n9255) );
  AND2X1 U4645 ( .A(n6043), .B(n9688), .Y(n10068) );
  AND2X1 U4646 ( .A(n6034), .B(n9632), .Y(n9986) );
  AND2X1 U4647 ( .A(n9626), .B(n6037), .Y(n10070) );
  AND2X1 U4648 ( .A(n6342), .B(n9639), .Y(n9783) );
  AND2X1 U4649 ( .A(n10291), .B(n6246), .Y(n9918) );
  AND2X1 U4650 ( .A(n6347), .B(n9577), .Y(n10177) );
  AND2X1 U4651 ( .A(n9577), .B(n6342), .Y(n9692) );
  AND2X1 U4652 ( .A(n6032), .B(n9639), .Y(n9844) );
  AND2X1 U4653 ( .A(n9695), .B(n6244), .Y(n9725) );
  AND2X1 U4654 ( .A(n6043), .B(n5769), .Y(n10232) );
  AND2X1 U4655 ( .A(n9688), .B(n6345), .Y(n10024) );
  AND2X1 U4656 ( .A(n6347), .B(n5769), .Y(n10282) );
  AND2X1 U4657 ( .A(n6345), .B(n9577), .Y(n9770) );
  AND2X1 U4658 ( .A(n6043), .B(n9639), .Y(n10178) );
  AND2X1 U4659 ( .A(n6032), .B(n9577), .Y(n9785) );
  AND2X1 U4660 ( .A(n21), .B(n10154), .Y(n10297) );
  BUFX2 U4661 ( .A(n6584), .Y(n4619) );
  BUFX2 U4662 ( .A(n6581), .Y(n4620) );
  BUFX2 U4663 ( .A(n7616), .Y(n4621) );
  BUFX2 U4664 ( .A(n7613), .Y(n4622) );
  BUFX2 U4665 ( .A(n8618), .Y(n4623) );
  BUFX2 U4666 ( .A(n8615), .Y(n4624) );
  BUFX2 U4667 ( .A(n9648), .Y(n4625) );
  BUFX2 U4668 ( .A(n9644), .Y(n4626) );
  AND2X1 U4669 ( .A(n6517), .B(n66), .Y(n6780) );
  INVX1 U4670 ( .A(n6780), .Y(n4627) );
  AND2X1 U4671 ( .A(n6579), .B(n5934), .Y(n7160) );
  INVX1 U4672 ( .A(n7160), .Y(n4628) );
  AND2X1 U4673 ( .A(n5821), .B(n6161), .Y(n6782) );
  INVX1 U4674 ( .A(n6782), .Y(n4629) );
  AND2X1 U4675 ( .A(n6579), .B(n5937), .Y(n7212) );
  INVX1 U4676 ( .A(n7212), .Y(n4630) );
  AND2X1 U4677 ( .A(n5931), .B(n6077), .Y(n7087) );
  INVX1 U4678 ( .A(n7087), .Y(n4631) );
  AND2X1 U4679 ( .A(n10290), .B(n6174), .Y(n7138) );
  INVX1 U4680 ( .A(n7138), .Y(n4632) );
  AND2X1 U4681 ( .A(n7550), .B(n5964), .Y(n7802) );
  INVX1 U4682 ( .A(n7802), .Y(n4633) );
  AND2X1 U4683 ( .A(n7611), .B(n5975), .Y(n8181) );
  INVX1 U4684 ( .A(n8181), .Y(n4634) );
  AND2X1 U4685 ( .A(n7611), .B(n6301), .Y(n8229) );
  INVX1 U4686 ( .A(n8229), .Y(n4635) );
  AND2X1 U4687 ( .A(n5973), .B(n9632), .Y(n8131) );
  INVX1 U4688 ( .A(n8131), .Y(n4636) );
  AND2X1 U4689 ( .A(n10290), .B(n6206), .Y(n8156) );
  INVX1 U4690 ( .A(n8156), .Y(n4637) );
  AND2X1 U4691 ( .A(n8554), .B(n43), .Y(n8809) );
  INVX1 U4692 ( .A(n8809), .Y(n4638) );
  AND2X1 U4693 ( .A(n8610), .B(n6330), .Y(n9192) );
  INVX1 U4694 ( .A(n9192), .Y(n4639) );
  INVX1 U4695 ( .A(n8811), .Y(n4640) );
  AND2X1 U4696 ( .A(n8610), .B(n6332), .Y(n9241) );
  INVX1 U4697 ( .A(n9241), .Y(n4641) );
  AND2X1 U4698 ( .A(n6328), .B(n9632), .Y(n9143) );
  INVX1 U4699 ( .A(n9143), .Y(n4642) );
  INVX1 U4700 ( .A(n9168), .Y(n4643) );
  AND2X1 U4701 ( .A(n5885), .B(n9577), .Y(n9843) );
  INVX1 U4702 ( .A(n9843), .Y(n4644) );
  AND2X1 U4703 ( .A(n6347), .B(n9639), .Y(n10231) );
  INVX1 U4704 ( .A(n10231), .Y(n4645) );
  INVX1 U4705 ( .A(n9845), .Y(n4646) );
  AND2X1 U4706 ( .A(n6049), .B(n9639), .Y(n10281) );
  INVX1 U4707 ( .A(n10281), .Y(n4647) );
  AND2X1 U4708 ( .A(n6043), .B(n6077), .Y(n10183) );
  INVX1 U4709 ( .A(n10183), .Y(n4648) );
  INVX1 U4710 ( .A(n10436), .Y(n4649) );
  INVX1 U4711 ( .A(n7156), .Y(n4651) );
  INVX1 U4712 ( .A(n8187), .Y(n4654) );
  INVX1 U4713 ( .A(n9198), .Y(n4657) );
  BUFX2 U4714 ( .A(n10239), .Y(n4659) );
  INVX1 U4715 ( .A(n153), .Y(n10239) );
  INVX1 U4716 ( .A(n10237), .Y(n4661) );
  AND2X1 U4717 ( .A(n6579), .B(n6277), .Y(n6922) );
  INVX1 U4718 ( .A(n6922), .Y(n4663) );
  AND2X1 U4719 ( .A(n66), .B(n6083), .Y(n6776) );
  INVX1 U4720 ( .A(n6776), .Y(n4664) );
  AND2X1 U4721 ( .A(n4708), .B(n6155), .Y(n6790) );
  INVX1 U4722 ( .A(n6790), .Y(n4665) );
  AND2X1 U4723 ( .A(n5933), .B(n6083), .Y(n7086) );
  INVX1 U4724 ( .A(n7086), .Y(n4666) );
  AND2X1 U4725 ( .A(n6551), .B(n5932), .Y(n7215) );
  INVX1 U4726 ( .A(n7215), .Y(n4667) );
  AND2X1 U4727 ( .A(n6517), .B(n5937), .Y(n7159) );
  INVX1 U4728 ( .A(n7159), .Y(n4668) );
  AND2X1 U4729 ( .A(n6286), .B(n9688), .Y(n7235) );
  INVX1 U4730 ( .A(n7235), .Y(n4669) );
  AND2X1 U4731 ( .A(n6517), .B(n6286), .Y(n7211) );
  INVX1 U4732 ( .A(n7211), .Y(n4670) );
  AND2X1 U4733 ( .A(n10291), .B(n6174), .Y(n7358) );
  INVX1 U4734 ( .A(n7358), .Y(n4671) );
  AND2X1 U4735 ( .A(n7611), .B(n45), .Y(n7942) );
  INVX1 U4736 ( .A(n7942), .Y(n4672) );
  AND2X1 U4737 ( .A(n5965), .B(n9688), .Y(n7798) );
  INVX1 U4738 ( .A(n7798), .Y(n4673) );
  INVX1 U4739 ( .A(n8130), .Y(n4674) );
  AND2X1 U4740 ( .A(n5975), .B(n9688), .Y(n8130) );
  AND2X1 U4741 ( .A(n7586), .B(n5973), .Y(n8232) );
  INVX1 U4742 ( .A(n8232), .Y(n4675) );
  AND2X1 U4743 ( .A(n7550), .B(n6301), .Y(n8180) );
  INVX1 U4744 ( .A(n8180), .Y(n4676) );
  AND2X1 U4745 ( .A(n6303), .B(n9688), .Y(n8249) );
  INVX1 U4746 ( .A(n8249), .Y(n4677) );
  AND2X1 U4747 ( .A(n7550), .B(n6303), .Y(n8228) );
  INVX1 U4748 ( .A(n8228), .Y(n4678) );
  AND2X1 U4749 ( .A(n10291), .B(n6206), .Y(n8374) );
  INVX1 U4750 ( .A(n8374), .Y(n4679) );
  AND2X1 U4751 ( .A(n8610), .B(n6319), .Y(n8948) );
  INVX1 U4752 ( .A(n8948), .Y(n4680) );
  INVX1 U4753 ( .A(n8805), .Y(n4681) );
  AND2X1 U4754 ( .A(n6330), .B(n9688), .Y(n9142) );
  INVX1 U4755 ( .A(n9142), .Y(n4682) );
  AND2X1 U4756 ( .A(n8588), .B(n6004), .Y(n9244) );
  INVX1 U4757 ( .A(n9244), .Y(n4683) );
  AND2X1 U4758 ( .A(n8554), .B(n6008), .Y(n9191) );
  INVX1 U4759 ( .A(n9191), .Y(n4684) );
  INVX1 U4760 ( .A(n9260), .Y(n4685) );
  INVX1 U4761 ( .A(n9240), .Y(n4686) );
  AND2X1 U4762 ( .A(n10291), .B(n6233), .Y(n9384) );
  INVX1 U4763 ( .A(n9384), .Y(n4687) );
  INVX1 U4764 ( .A(n9988), .Y(n4688) );
  AND2X1 U4765 ( .A(n6034), .B(n9639), .Y(n9988) );
  AND2X1 U4766 ( .A(n9688), .B(n5885), .Y(n9839) );
  INVX1 U4767 ( .A(n9839), .Y(n4689) );
  AND2X1 U4768 ( .A(n6042), .B(n9614), .Y(n10284) );
  INVX1 U4769 ( .A(n10284), .Y(n4690) );
  AND2X1 U4770 ( .A(n6049), .B(n9577), .Y(n10230) );
  INVX1 U4771 ( .A(n10230), .Y(n4691) );
  INVX1 U4772 ( .A(n10302), .Y(n4692) );
  INVX1 U4773 ( .A(n10280), .Y(n4693) );
  INVX1 U4774 ( .A(n10208), .Y(n4694) );
  AND2X1 U4775 ( .A(n7490), .B(n6731), .Y(n6730) );
  INVX1 U4776 ( .A(n6730), .Y(n4695) );
  AND2X1 U4777 ( .A(n7233), .B(oprB[61]), .Y(n6787) );
  INVX1 U4778 ( .A(n6787), .Y(n4696) );
  AND2X1 U4779 ( .A(n6570), .B(n6155), .Y(n7147) );
  INVX1 U4780 ( .A(n7147), .Y(n4697) );
  AND2X1 U4781 ( .A(n9258), .B(n5907), .Y(n8816) );
  INVX1 U4782 ( .A(n8816), .Y(n4698) );
  INVX1 U4783 ( .A(n7089), .Y(n4699) );
  AND2X1 U4784 ( .A(n5748), .B(n8299), .Y(n8355) );
  INVX1 U4785 ( .A(n8355), .Y(n4700) );
  AND2X1 U4786 ( .A(n9498), .B(n9310), .Y(n9365) );
  INVX1 U4787 ( .A(n9365), .Y(n4701) );
  AND2X1 U4788 ( .A(n10290), .B(n6245), .Y(n9784) );
  INVX1 U4789 ( .A(n9784), .Y(n4702) );
  AND2X1 U4790 ( .A(n10498), .B(n10355), .Y(n10417) );
  INVX1 U4791 ( .A(n10417), .Y(n4703) );
  AND2X1 U4792 ( .A(n6282), .B(n6080), .Y(n7158) );
  INVX1 U4793 ( .A(n7158), .Y(n4704) );
  AND2X1 U4794 ( .A(n6297), .B(n6080), .Y(n8189) );
  INVX1 U4795 ( .A(n8189), .Y(n4705) );
  AND2X1 U4796 ( .A(n6325), .B(n6080), .Y(n9200) );
  INVX1 U4797 ( .A(n9200), .Y(n4706) );
  AND2X1 U4798 ( .A(n5800), .B(n6345), .Y(n10240) );
  INVX1 U4799 ( .A(n10240), .Y(n4707) );
  INVX1 U4800 ( .A(n6506), .Y(n4708) );
  AND2X1 U4801 ( .A(n5449), .B(n5362), .Y(n6506) );
  AND2X1 U4802 ( .A(n5931), .B(n6080), .Y(n7236) );
  INVX1 U4803 ( .A(n7236), .Y(n4709) );
  AND2X1 U4804 ( .A(n5974), .B(n6080), .Y(n8250) );
  INVX1 U4805 ( .A(n8250), .Y(n4710) );
  AND2X1 U4806 ( .A(n6004), .B(n6080), .Y(n9261) );
  INVX1 U4807 ( .A(n9261), .Y(n4711) );
  INVX1 U4808 ( .A(n10303), .Y(n4712) );
  AND2X1 U4809 ( .A(n6191), .B(n5821), .Y(n8362) );
  INVX1 U4810 ( .A(n8362), .Y(n4713) );
  INVX1 U4811 ( .A(n10424), .Y(n4714) );
  AND2X1 U4812 ( .A(n5705), .B(n6190), .Y(n8097) );
  INVX1 U4813 ( .A(n8097), .Y(n4715) );
  AND2X1 U4814 ( .A(n5706), .B(n6246), .Y(n10149) );
  INVX1 U4815 ( .A(n10149), .Y(n4716) );
  BUFX2 U4816 ( .A(n7345), .Y(n4717) );
  BUFX2 U4817 ( .A(n7860), .Y(n4718) );
  INVX1 U4818 ( .A(n4720), .Y(n4719) );
  BUFX2 U4819 ( .A(n8361), .Y(n4720) );
  BUFX2 U4820 ( .A(n9904), .Y(n4721) );
  AND2X1 U4821 ( .A(n5738), .B(n10376), .Y(n10423) );
  INVX1 U4822 ( .A(n10423), .Y(n4722) );
  BUFX2 U4823 ( .A(n9627), .Y(n4723) );
  AND2X1 U4824 ( .A(n6551), .B(n6275), .Y(n6924) );
  INVX1 U4825 ( .A(n6924), .Y(n4724) );
  AND2X1 U4826 ( .A(n6517), .B(n6627), .Y(n7488) );
  INVX1 U4827 ( .A(n7488), .Y(n4725) );
  AND2X1 U4828 ( .A(n5937), .B(n6077), .Y(n7239) );
  INVX1 U4829 ( .A(n7239), .Y(n4726) );
  AND2X1 U4830 ( .A(n6551), .B(n6277), .Y(n7016) );
  INVX1 U4831 ( .A(n7016), .Y(n4727) );
  AND2X1 U4832 ( .A(n6551), .B(n6279), .Y(n7090) );
  INVX1 U4833 ( .A(n7090), .Y(n4728) );
  AND2X1 U4834 ( .A(n7586), .B(n5961), .Y(n7944) );
  INVX1 U4835 ( .A(n7944), .Y(n4729) );
  AND2X1 U4836 ( .A(n7586), .B(n6297), .Y(n8184) );
  INVX1 U4837 ( .A(n8184), .Y(n4730) );
  AND2X1 U4838 ( .A(n7550), .B(n7656), .Y(n8496) );
  INVX1 U4839 ( .A(n8496), .Y(n4731) );
  AND2X1 U4840 ( .A(n5767), .B(n5961), .Y(n7867) );
  INVX1 U4841 ( .A(n7867), .Y(n4732) );
  AND2X1 U4842 ( .A(n6301), .B(n9632), .Y(n8253) );
  INVX1 U4843 ( .A(n8253), .Y(n4733) );
  AND2X1 U4844 ( .A(n7586), .B(n45), .Y(n8029) );
  INVX1 U4845 ( .A(n8029), .Y(n4734) );
  AND2X1 U4846 ( .A(n7586), .B(n6296), .Y(n8123) );
  INVX1 U4847 ( .A(n8123), .Y(n4735) );
  AND2X1 U4848 ( .A(n8588), .B(n5276), .Y(n8950) );
  INVX1 U4849 ( .A(n8950), .Y(n4736) );
  AND2X1 U4850 ( .A(n8679), .B(n8554), .Y(n9508) );
  INVX1 U4851 ( .A(n9508), .Y(n4737) );
  AND2X1 U4852 ( .A(n5768), .B(n5276), .Y(n8874) );
  INVX1 U4853 ( .A(n8874), .Y(n4738) );
  AND2X1 U4854 ( .A(n6332), .B(n9632), .Y(n9264) );
  INVX1 U4855 ( .A(n9264), .Y(n4739) );
  AND2X1 U4856 ( .A(n8588), .B(n6319), .Y(n9040) );
  INVX1 U4857 ( .A(n9040), .Y(n4740) );
  INVX1 U4858 ( .A(n9135), .Y(n4741) );
  AND2X1 U4859 ( .A(n8588), .B(n6322), .Y(n9135) );
  AND2X1 U4860 ( .A(n6032), .B(n9614), .Y(n9990) );
  INVX1 U4861 ( .A(n9990), .Y(n4742) );
  AND2X1 U4862 ( .A(n6345), .B(n9614), .Y(n10234) );
  INVX1 U4863 ( .A(n10234), .Y(n4743) );
  AND2X1 U4864 ( .A(n9577), .B(n9689), .Y(n10554) );
  INVX1 U4865 ( .A(n10554), .Y(n4744) );
  AND2X1 U4866 ( .A(n6032), .B(n5769), .Y(n9911) );
  INVX1 U4867 ( .A(n9911), .Y(n4745) );
  AND2X1 U4868 ( .A(n6049), .B(n9632), .Y(n10306) );
  INVX1 U4869 ( .A(n10306), .Y(n4746) );
  AND2X1 U4870 ( .A(n6034), .B(n9614), .Y(n10076) );
  INVX1 U4871 ( .A(n10076), .Y(n4747) );
  INVX1 U4872 ( .A(n10175), .Y(n4748) );
  AND2X1 U4873 ( .A(n6037), .B(n9614), .Y(n10175) );
  INVX1 U4874 ( .A(n6517), .Y(n4749) );
  AND2X1 U4875 ( .A(n5902), .B(n5899), .Y(n6733) );
  INVX1 U4876 ( .A(n6733), .Y(n4750) );
  AND2X1 U4877 ( .A(n5902), .B(n6160), .Y(n6974) );
  INVX1 U4878 ( .A(n6974), .Y(n4751) );
  AND2X1 U4879 ( .A(n6156), .B(n5890), .Y(n6731) );
  INVX1 U4880 ( .A(n6731), .Y(n4752) );
  AND2X1 U4881 ( .A(n6186), .B(n6188), .Y(n7550) );
  INVX1 U4882 ( .A(n7550), .Y(n4753) );
  AND2X1 U4883 ( .A(n6191), .B(n6189), .Y(n7755) );
  INVX1 U4884 ( .A(n7755), .Y(n4754) );
  AND2X1 U4885 ( .A(n6191), .B(n6190), .Y(n7988) );
  INVX1 U4886 ( .A(n7988), .Y(n4755) );
  AND2X1 U4887 ( .A(n6220), .B(n5907), .Y(n8762) );
  INVX1 U4888 ( .A(n8762), .Y(n4756) );
  AND2X1 U4889 ( .A(n5883), .B(n6219), .Y(n8999) );
  INVX1 U4890 ( .A(n8999), .Y(n4757) );
  INVX1 U4891 ( .A(n9577), .Y(n4758) );
  INVX1 U4892 ( .A(n9792), .Y(n4759) );
  INVX1 U4893 ( .A(n10034), .Y(n4760) );
  INVX1 U4894 ( .A(n10498), .Y(n4761) );
  AND2X1 U4895 ( .A(n5719), .B(n5363), .Y(n8171) );
  INVX1 U4896 ( .A(n8171), .Y(n4762) );
  INVX1 U4897 ( .A(n8127), .Y(n4763) );
  INVX1 U4898 ( .A(n9139), .Y(n4764) );
  INVX1 U4899 ( .A(n9475), .Y(n4765) );
  INVX1 U4900 ( .A(n10179), .Y(n4766) );
  INVX1 U4901 ( .A(n10499), .Y(n4767) );
  INVX1 U4902 ( .A(n6551), .Y(n4768) );
  INVX1 U4903 ( .A(n6778), .Y(n4769) );
  AND2X1 U4904 ( .A(n5820), .B(n5918), .Y(n6778) );
  INVX1 U4905 ( .A(n6966), .Y(n4770) );
  INVX1 U4906 ( .A(n6925), .Y(n4771) );
  INVX1 U4907 ( .A(n6967), .Y(n4772) );
  AND2X1 U4908 ( .A(n5820), .B(n6277), .Y(n6967) );
  AND2X1 U4909 ( .A(n7284), .B(n6286), .Y(n7241) );
  INVX1 U4910 ( .A(n7241), .Y(n4773) );
  INVX1 U4911 ( .A(n7586), .Y(n4774) );
  INVX1 U4912 ( .A(n7800), .Y(n4775) );
  AND2X1 U4913 ( .A(n5767), .B(n5957), .Y(n7800) );
  INVX1 U4914 ( .A(n7982), .Y(n4776) );
  AND2X1 U4915 ( .A(n7586), .B(n5964), .Y(n7982) );
  INVX1 U4916 ( .A(n7945), .Y(n4777) );
  AND2X1 U4917 ( .A(n5767), .B(n5964), .Y(n7945) );
  AND2X1 U4918 ( .A(n5767), .B(n5966), .Y(n7983) );
  INVX1 U4919 ( .A(n7983), .Y(n4778) );
  AND2X1 U4920 ( .A(n8299), .B(n6303), .Y(n8255) );
  INVX1 U4921 ( .A(n8255), .Y(n4779) );
  INVX1 U4922 ( .A(n8588), .Y(n4780) );
  INVX1 U4923 ( .A(n8807), .Y(n4781) );
  AND2X1 U4924 ( .A(n5768), .B(n6315), .Y(n8807) );
  INVX1 U4925 ( .A(n8994), .Y(n4782) );
  AND2X1 U4926 ( .A(n8588), .B(n43), .Y(n8994) );
  AND2X1 U4927 ( .A(n5768), .B(n43), .Y(n8951) );
  INVX1 U4928 ( .A(n8951), .Y(n4783) );
  AND2X1 U4929 ( .A(n5768), .B(n6319), .Y(n8995) );
  INVX1 U4930 ( .A(n8995), .Y(n4784) );
  INVX1 U4931 ( .A(n9614), .Y(n4785) );
  INVX1 U4932 ( .A(n9841), .Y(n4786) );
  AND2X1 U4933 ( .A(n6029), .B(n5769), .Y(n9841) );
  AND2X1 U4934 ( .A(n5885), .B(n9614), .Y(n10028) );
  INVX1 U4935 ( .A(n10028), .Y(n4787) );
  AND2X1 U4936 ( .A(n5885), .B(n5769), .Y(n9991) );
  INVX1 U4937 ( .A(n9991), .Y(n4788) );
  AND2X1 U4938 ( .A(n6034), .B(n5769), .Y(n10029) );
  INVX1 U4939 ( .A(n10029), .Y(n4789) );
  AND2X1 U4940 ( .A(n7491), .B(n6245), .Y(n10370) );
  INVX1 U4941 ( .A(n10370), .Y(n4790) );
  BUFX2 U4942 ( .A(n10497), .Y(n4791) );
  INVX1 U4943 ( .A(n154), .Y(n10497) );
  INVX1 U4944 ( .A(n10215), .Y(n4793) );
  AND2X1 U4945 ( .A(n7146), .B(n5889), .Y(n6721) );
  INVX1 U4946 ( .A(n6721), .Y(n4795) );
  AND2X1 U4947 ( .A(n9629), .B(n6083), .Y(n6971) );
  INVX1 U4948 ( .A(n6971), .Y(n4796) );
  AND2X1 U4949 ( .A(n5447), .B(n6155), .Y(n7407) );
  INVX1 U4950 ( .A(n7407), .Y(n4797) );
  AND2X1 U4951 ( .A(n6169), .B(n6172), .Y(n7070) );
  INVX1 U4952 ( .A(n7070), .Y(n4798) );
  INVX1 U4953 ( .A(n7611), .Y(n4799) );
  AND2X1 U4954 ( .A(n6201), .B(n6204), .Y(n8102) );
  INVX1 U4955 ( .A(n8102), .Y(n4800) );
  AND2X1 U4956 ( .A(n8299), .B(n5975), .Y(n8112) );
  INVX1 U4957 ( .A(n8112), .Y(n4801) );
  INVX1 U4958 ( .A(n8610), .Y(n4802) );
  INVX1 U4959 ( .A(n9114), .Y(n4803) );
  INVX1 U4960 ( .A(n9124), .Y(n4804) );
  AND2X1 U4961 ( .A(n9310), .B(n6330), .Y(n9124) );
  INVX1 U4962 ( .A(n9639), .Y(n4805) );
  INVX1 U4963 ( .A(n10154), .Y(n4806) );
  INVX1 U4964 ( .A(n10164), .Y(n4807) );
  AND2X1 U4965 ( .A(n10355), .B(n6347), .Y(n10164) );
  INVX1 U4966 ( .A(n6703), .Y(n4809) );
  BUFX2 U4967 ( .A(n7971), .Y(n4811) );
  INVX1 U4968 ( .A(n155), .Y(n7971) );
  INVX1 U4969 ( .A(n7731), .Y(n4813) );
  INVX1 U4970 ( .A(n8737), .Y(n4816) );
  BUFX2 U4971 ( .A(n9496), .Y(n4818) );
  INVX1 U4972 ( .A(n156), .Y(n9496) );
  INVX1 U4973 ( .A(n9254), .Y(n4820) );
  BUFX2 U4974 ( .A(n10017), .Y(n4822) );
  INVX1 U4975 ( .A(n157), .Y(n10017) );
  INVX1 U4976 ( .A(n9766), .Y(n4824) );
  INVX1 U4977 ( .A(n7308), .Y(n4826) );
  INVX1 U4978 ( .A(n8324), .Y(n4827) );
  INVX1 U4979 ( .A(n9334), .Y(n4828) );
  INVX1 U4980 ( .A(n10386), .Y(n4829) );
  INVX1 U4981 ( .A(n6628), .Y(n4830) );
  AND2X1 U4982 ( .A(n7611), .B(n5955), .Y(n7657) );
  INVX1 U4983 ( .A(n7657), .Y(n4831) );
  INVX1 U4984 ( .A(n8677), .Y(n4832) );
  AND2X1 U4985 ( .A(n6026), .B(n9639), .Y(n9690) );
  INVX1 U4986 ( .A(n9690), .Y(n4833) );
  BUFX2 U4987 ( .A(n6578), .Y(n4834) );
  BUFX2 U4988 ( .A(n6572), .Y(n4835) );
  BUFX2 U4989 ( .A(n7069), .Y(n4836) );
  BUFX2 U4990 ( .A(n7610), .Y(n4837) );
  BUFX2 U4991 ( .A(n7604), .Y(n4838) );
  BUFX2 U4992 ( .A(n8105), .Y(n4839) );
  BUFX2 U4993 ( .A(n8609), .Y(n4840) );
  BUFX2 U4994 ( .A(n8606), .Y(n4841) );
  BUFX2 U4995 ( .A(n9117), .Y(n4842) );
  BUFX2 U4996 ( .A(n9638), .Y(n4843) );
  BUFX2 U4997 ( .A(n9635), .Y(n4844) );
  BUFX2 U4998 ( .A(n10157), .Y(n4845) );
  BUFX2 U4999 ( .A(n7415), .Y(n4846) );
  BUFX2 U5000 ( .A(n10520), .Y(n4847) );
  INVX1 U5001 ( .A(n10556), .Y(n4848) );
  INVX1 U5002 ( .A(n6848), .Y(n4850) );
  INVX1 U5003 ( .A(n9194), .Y(n4853) );
  INVX1 U5004 ( .A(n7492), .Y(n4855) );
  INVX1 U5005 ( .A(n8497), .Y(n4856) );
  INVX1 U5006 ( .A(n9509), .Y(n4857) );
  AND2X1 U5007 ( .A(n8247), .B(n6189), .Y(n7809) );
  INVX1 U5008 ( .A(n7809), .Y(n4858) );
  AND2X1 U5009 ( .A(n10300), .B(n6245), .Y(n9851) );
  INVX1 U5010 ( .A(n9851), .Y(n4859) );
  INVX1 U5011 ( .A(n7162), .Y(n4861) );
  INVX1 U5012 ( .A(n10296), .Y(n4864) );
  INVX1 U5013 ( .A(n6867), .Y(n4866) );
  INVX1 U5014 ( .A(n7886), .Y(n4867) );
  INVX1 U5015 ( .A(n8892), .Y(n4868) );
  INVX1 U5016 ( .A(n9931), .Y(n4869) );
  AND2X1 U5017 ( .A(n6551), .B(n6282), .Y(n7163) );
  INVX1 U5018 ( .A(n7163), .Y(n4870) );
  AND2X1 U5019 ( .A(n8588), .B(n6325), .Y(n9195) );
  INVX1 U5020 ( .A(n9195), .Y(n4871) );
  AND2X1 U5021 ( .A(n5820), .B(n6275), .Y(n6849) );
  INVX1 U5022 ( .A(n6849), .Y(n4872) );
  INVX1 U5023 ( .A(n9266), .Y(n4873) );
  INVX1 U5024 ( .A(n10308), .Y(n4874) );
  INVX1 U5025 ( .A(n7421), .Y(n4875) );
  BUFX2 U5026 ( .A(n10575), .Y(n4876) );
  INVX1 U5027 ( .A(n8873), .Y(n4878) );
  INVX1 U5028 ( .A(n6702), .Y(n4881) );
  INVX1 U5029 ( .A(n7229), .Y(n4884) );
  INVX1 U5030 ( .A(n7730), .Y(n4887) );
  INVX1 U5031 ( .A(n8231), .Y(n4890) );
  INVX1 U5032 ( .A(n8736), .Y(n4893) );
  INVX1 U5033 ( .A(n9765), .Y(n4896) );
  BUFX2 U5034 ( .A(n7422), .Y(n4898) );
  BUFX2 U5035 ( .A(n7476), .Y(n4899) );
  BUFX2 U5036 ( .A(n8419), .Y(n4900) );
  BUFX2 U5037 ( .A(n8483), .Y(n4901) );
  BUFX2 U5038 ( .A(n9492), .Y(n4902) );
  INVX1 U5039 ( .A(n7866), .Y(n4904) );
  INVX1 U5040 ( .A(n9910), .Y(n4907) );
  INVX1 U5041 ( .A(n7014), .Y(n4910) );
  INVX1 U5042 ( .A(n7091), .Y(n4913) );
  INVX1 U5043 ( .A(n8027), .Y(n4916) );
  INVX1 U5044 ( .A(n8183), .Y(n4919) );
  INVX1 U5045 ( .A(n8243), .Y(n4922) );
  INVX1 U5046 ( .A(n9038), .Y(n4925) );
  INVX1 U5047 ( .A(n9243), .Y(n4928) );
  INVX1 U5048 ( .A(n10074), .Y(n4931) );
  INVX1 U5049 ( .A(n10233), .Y(n4934) );
  INVX1 U5050 ( .A(n10283), .Y(n4937) );
  INVX1 U5051 ( .A(n6853), .Y(n4939) );
  INVX1 U5052 ( .A(n6868), .Y(n4940) );
  AND2X1 U5053 ( .A(n5564), .B(n9846), .Y(n7871) );
  INVX1 U5054 ( .A(n7871), .Y(n4941) );
  INVX1 U5055 ( .A(n7887), .Y(n4942) );
  INVX1 U5056 ( .A(n8447), .Y(n4943) );
  INVX1 U5057 ( .A(n8878), .Y(n4944) );
  INVX1 U5058 ( .A(n8893), .Y(n4945) );
  INVX1 U5059 ( .A(n9915), .Y(n4946) );
  INVX1 U5060 ( .A(n9932), .Y(n4947) );
  INVX1 U5061 ( .A(n8239), .Y(n4948) );
  INVX1 U5062 ( .A(n6496), .Y(n4950) );
  INVX1 U5063 ( .A(n7537), .Y(n4953) );
  INVX1 U5064 ( .A(n8541), .Y(n4956) );
  BUFX2 U5065 ( .A(n9457), .Y(n4958) );
  INVX1 U5066 ( .A(n9564), .Y(n4960) );
  BUFX2 U5067 ( .A(n6783), .Y(n4962) );
  BUFX2 U5068 ( .A(n7805), .Y(n4963) );
  BUFX2 U5069 ( .A(n8812), .Y(n4964) );
  BUFX2 U5070 ( .A(n9847), .Y(n4965) );
  AND2X1 U5071 ( .A(n5820), .B(n6279), .Y(n7015) );
  INVX1 U5072 ( .A(n7015), .Y(n4966) );
  AND2X1 U5073 ( .A(n5933), .B(n6081), .Y(n7237) );
  INVX1 U5074 ( .A(n7237), .Y(n4967) );
  AND2X1 U5075 ( .A(n5767), .B(n6296), .Y(n8028) );
  INVX1 U5076 ( .A(n8028), .Y(n4968) );
  AND2X1 U5077 ( .A(n5975), .B(n9626), .Y(n8251) );
  INVX1 U5078 ( .A(n8251), .Y(n4969) );
  AND2X1 U5079 ( .A(n5768), .B(n6322), .Y(n9039) );
  INVX1 U5080 ( .A(n9039), .Y(n4970) );
  AND2X1 U5081 ( .A(n6330), .B(n6081), .Y(n9262) );
  INVX1 U5082 ( .A(n9262), .Y(n4971) );
  AND2X1 U5083 ( .A(n6037), .B(n5769), .Y(n10075) );
  INVX1 U5084 ( .A(n10075), .Y(n4972) );
  AND2X1 U5085 ( .A(n6347), .B(n6081), .Y(n10304) );
  INVX1 U5086 ( .A(n10304), .Y(n4973) );
  INVX1 U5087 ( .A(n7010), .Y(n4977) );
  INVX1 U5088 ( .A(n7214), .Y(n4980) );
  INVX1 U5089 ( .A(n8023), .Y(n4985) );
  INVX1 U5090 ( .A(n8124), .Y(n4988) );
  INVX1 U5091 ( .A(n9034), .Y(n4993) );
  INVX1 U5092 ( .A(n9136), .Y(n4996) );
  INVX1 U5093 ( .A(n10069), .Y(n5001) );
  INVX1 U5094 ( .A(n10176), .Y(n5004) );
  AND2X1 U5095 ( .A(n10290), .B(n6190), .Y(n7873) );
  INVX1 U5096 ( .A(n7873), .Y(n5006) );
  AND2X1 U5097 ( .A(n10290), .B(n6246), .Y(n9917) );
  INVX1 U5098 ( .A(n9917), .Y(n5007) );
  AND2X1 U5099 ( .A(n5841), .B(n9647), .Y(n6866) );
  INVX1 U5100 ( .A(n6866), .Y(n5008) );
  AND2X1 U5101 ( .A(n5799), .B(n9647), .Y(n7885) );
  INVX1 U5102 ( .A(n7885), .Y(n5009) );
  INVX1 U5103 ( .A(n8891), .Y(n5010) );
  AND2X1 U5104 ( .A(n5798), .B(n9647), .Y(n8891) );
  AND2X1 U5105 ( .A(n5794), .B(n9647), .Y(n9930) );
  INVX1 U5106 ( .A(n9930), .Y(n5011) );
  AND2X1 U5107 ( .A(n5890), .B(n6556), .Y(n7351) );
  INVX1 U5108 ( .A(n7351), .Y(n5012) );
  INVX1 U5109 ( .A(n6706), .Y(n5014) );
  INVX1 U5110 ( .A(n7733), .Y(n5017) );
  INVX1 U5111 ( .A(n8740), .Y(n5020) );
  INVX1 U5112 ( .A(n9768), .Y(n5023) );
  INVX1 U5113 ( .A(n6582), .Y(n5026) );
  INVX1 U5114 ( .A(mult32_A[27]), .Y(n5028) );
  AND2X1 U5115 ( .A(n6517), .B(n10487), .Y(n7221) );
  INVX1 U5116 ( .A(n7221), .Y(n5029) );
  AND2X1 U5117 ( .A(n7550), .B(n10487), .Y(n8238) );
  INVX1 U5118 ( .A(n8238), .Y(n5030) );
  AND2X1 U5119 ( .A(n8554), .B(n10487), .Y(n9250) );
  INVX1 U5120 ( .A(n9250), .Y(n5031) );
  AND2X1 U5121 ( .A(n10487), .B(n9577), .Y(n10292) );
  INVX1 U5122 ( .A(n10292), .Y(n5032) );
  INVX1 U5123 ( .A(n8949), .Y(n5034) );
  INVX1 U5124 ( .A(n6786), .Y(n5037) );
  INVX1 U5125 ( .A(n8815), .Y(n5040) );
  BUFX2 U5126 ( .A(n9454), .Y(n5042) );
  INVX1 U5127 ( .A(n6909), .Y(n5044) );
  INVX1 U5128 ( .A(n8935), .Y(n5047) );
  INVX1 U5129 ( .A(mult32_A[28]), .Y(n5049) );
  INVX1 U5130 ( .A(n9989), .Y(n5051) );
  INVX1 U5131 ( .A(n8993), .Y(n5054) );
  INVX1 U5132 ( .A(n7943), .Y(n5057) );
  INVX1 U5133 ( .A(n6923), .Y(n5060) );
  AND2X1 U5134 ( .A(n9626), .B(n6625), .Y(n10378) );
  AND2X1 U5135 ( .A(n5800), .B(n6625), .Y(n10381) );
  INVX1 U5136 ( .A(n9838), .Y(n5063) );
  INVX1 U5137 ( .A(n7797), .Y(n5066) );
  INVX1 U5138 ( .A(n6961), .Y(n5069) );
  INVX1 U5139 ( .A(n7614), .Y(n5072) );
  INVX1 U5140 ( .A(n8616), .Y(n5075) );
  INVX1 U5141 ( .A(n9645), .Y(n5078) );
  INVX1 U5142 ( .A(n6483), .Y(n5081) );
  INVX1 U5143 ( .A(n7981), .Y(n5084) );
  INVX1 U5144 ( .A(n8531), .Y(n5087) );
  INVX1 U5145 ( .A(n8743), .Y(n5090) );
  INVX1 U5146 ( .A(n10027), .Y(n5093) );
  INVX1 U5147 ( .A(n6775), .Y(n5096) );
  INVX1 U5148 ( .A(n8804), .Y(n5099) );
  INVX1 U5149 ( .A(n7939), .Y(n5102) );
  INVX1 U5150 ( .A(n8325), .Y(n5104) );
  INVX1 U5151 ( .A(n9335), .Y(n5105) );
  INVX1 U5152 ( .A(n10387), .Y(n5106) );
  INVX1 U5153 ( .A(n6709), .Y(n5108) );
  INVX1 U5154 ( .A(n6965), .Y(n5111) );
  INVX1 U5155 ( .A(n7527), .Y(n5114) );
  INVX1 U5156 ( .A(n7587), .Y(n5117) );
  INVX1 U5157 ( .A(n7736), .Y(n5120) );
  INVX1 U5158 ( .A(n7801), .Y(n5123) );
  INVX1 U5159 ( .A(n9554), .Y(n5126) );
  INVX1 U5160 ( .A(n9615), .Y(n5129) );
  INVX1 U5161 ( .A(n9771), .Y(n5132) );
  INVX1 U5162 ( .A(n9842), .Y(n5135) );
  INVX1 U5163 ( .A(n9985), .Y(n5138) );
  INVX1 U5164 ( .A(n6485), .Y(n5141) );
  INVX1 U5165 ( .A(n7529), .Y(n5144) );
  INVX1 U5166 ( .A(n8533), .Y(n5147) );
  INVX1 U5167 ( .A(n9556), .Y(n5150) );
  INVX1 U5168 ( .A(n7977), .Y(n5153) );
  INVX1 U5169 ( .A(n8989), .Y(n5156) );
  INVX1 U5170 ( .A(n7309), .Y(n5158) );
  INVX1 U5171 ( .A(n6552), .Y(n5160) );
  INVX1 U5172 ( .A(n6779), .Y(n5163) );
  INVX1 U5173 ( .A(n8589), .Y(n5166) );
  INVX1 U5174 ( .A(n8808), .Y(n5169) );
  INVX1 U5175 ( .A(n10023), .Y(n5172) );
  AND2X1 U5176 ( .A(n10290), .B(n6219), .Y(n8946) );
  INVX1 U5177 ( .A(n8946), .Y(n5174) );
  INVX1 U5178 ( .A(n10377), .Y(n5176) );
  INVX1 U5179 ( .A(n10367), .Y(n5181) );
  INVX1 U5180 ( .A(n7475), .Y(n5183) );
  INVX1 U5181 ( .A(n8482), .Y(n5184) );
  INVX1 U5182 ( .A(n9322), .Y(n5186) );
  INVX1 U5183 ( .A(n6640), .Y(n5189) );
  INVX1 U5184 ( .A(n7668), .Y(n5192) );
  INVX1 U5185 ( .A(n8684), .Y(n5195) );
  INVX1 U5186 ( .A(n9700), .Y(n5198) );
  INVX1 U5187 ( .A(n8753), .Y(n5201) );
  INVX1 U5188 ( .A(n10388), .Y(n5207) );
  INVX1 U5189 ( .A(n7310), .Y(n5214) );
  INVX1 U5190 ( .A(n8326), .Y(n5215) );
  INVX1 U5191 ( .A(n9336), .Y(n5216) );
  INVX1 U5192 ( .A(n9330), .Y(n5218) );
  INVX1 U5193 ( .A(n10380), .Y(n5221) );
  INVX1 U5194 ( .A(n9328), .Y(n5224) );
  INVX1 U5195 ( .A(n7296), .Y(n5227) );
  INVX1 U5196 ( .A(n8312), .Y(n5230) );
  INVX1 U5197 ( .A(n9782), .Y(n5233) );
  INVX1 U5198 ( .A(n7318), .Y(n5235) );
  INVX1 U5199 ( .A(n9344), .Y(n5236) );
  INVX1 U5200 ( .A(n10569), .Y(n5237) );
  INVX1 U5201 ( .A(n9502), .Y(n5238) );
  AND2X1 U5202 ( .A(n9632), .B(n6625), .Y(n10368) );
  INVX1 U5203 ( .A(n7302), .Y(n5240) );
  INVX1 U5204 ( .A(n7304), .Y(n5243) );
  INVX1 U5205 ( .A(n7746), .Y(n5246) );
  INVX1 U5206 ( .A(n8318), .Y(n5249) );
  INVX1 U5207 ( .A(n8320), .Y(n5252) );
  INVX1 U5208 ( .A(n8334), .Y(n5254) );
  INVX1 U5209 ( .A(n10396), .Y(n5255) );
  INVX1 U5210 ( .A(n6719), .Y(n5261) );
  BUFX2 U5211 ( .A(n10555), .Y(n5263) );
  INVX1 U5212 ( .A(n5265), .Y(n5264) );
  BUFX2 U5213 ( .A(n10557), .Y(n5265) );
  INVX2 U5214 ( .A(n5898), .Y(n5899) );
  AND2X2 U5215 ( .A(n6061), .B(n6261), .Y(n5765) );
  INVX2 U5216 ( .A(oprB[29]), .Y(n6219) );
  AND2X1 U5217 ( .A(n5639), .B(n6219), .Y(n9109) );
  BUFX2 U5218 ( .A(n6024), .Y(n5272) );
  INVX1 U5219 ( .A(n6010), .Y(n6011) );
  AND2X2 U5220 ( .A(n46), .B(n19), .Y(n9175) );
  INVX8 U5221 ( .A(n6248), .Y(n6247) );
  INVX8 U5222 ( .A(n6313), .Y(n5992) );
  INVX8 U5223 ( .A(n6218), .Y(n6217) );
  BUFX4 U5224 ( .A(oprA[28]), .Y(n5276) );
  BUFX4 U5225 ( .A(oprA[19]), .Y(n5278) );
  INVX1 U5226 ( .A(n6318), .Y(n5998) );
  INVX1 U5227 ( .A(n6236), .Y(n5279) );
  BUFX2 U5228 ( .A(oprA[17]), .Y(n5281) );
  BUFX2 U5229 ( .A(n6337), .Y(n5282) );
  BUFX4 U5230 ( .A(oprA[25]), .Y(n5283) );
  INVX8 U5231 ( .A(n6225), .Y(n6224) );
  BUFX4 U5232 ( .A(n6015), .Y(n5286) );
  INVX1 U5233 ( .A(n6454), .Y(n5287) );
  AND2X1 U5234 ( .A(n6085), .B(n7253), .Y(n7254) );
  INVX1 U5235 ( .A(n7254), .Y(n5288) );
  AND2X1 U5236 ( .A(n3145), .B(n5776), .Y(n9547) );
  INVX1 U5237 ( .A(n9547), .Y(n5289) );
  AND2X1 U5238 ( .A(n6076), .B(n6054), .Y(n6466) );
  INVX1 U5239 ( .A(n6466), .Y(n5290) );
  AND2X1 U5240 ( .A(n6085), .B(n7820), .Y(n7821) );
  INVX1 U5241 ( .A(n7821), .Y(n5291) );
  AND2X1 U5242 ( .A(n3146), .B(n5776), .Y(n9607) );
  INVX1 U5243 ( .A(n9607), .Y(n5292) );
  AND2X1 U5244 ( .A(n6076), .B(n6332), .Y(n6445) );
  INVX1 U5245 ( .A(n6445), .Y(n5293) );
  AND2X1 U5246 ( .A(n6076), .B(n6347), .Y(n6463) );
  INVX1 U5247 ( .A(n6463), .Y(n5294) );
  AND2X1 U5248 ( .A(n6085), .B(n8827), .Y(n8828) );
  INVX1 U5249 ( .A(n8828), .Y(n5295) );
  AND2X1 U5250 ( .A(n3147), .B(n5776), .Y(n9685) );
  INVX1 U5251 ( .A(n9685), .Y(n5296) );
  AND2X1 U5252 ( .A(n6076), .B(n6322), .Y(n6441) );
  INVX1 U5253 ( .A(n6441), .Y(n5297) );
  INVX1 U5254 ( .A(n6465), .Y(n5298) );
  AND2X1 U5255 ( .A(n6085), .B(n9863), .Y(n9864) );
  INVX1 U5256 ( .A(n9864), .Y(n5299) );
  AND2X1 U5257 ( .A(n3148), .B(n5776), .Y(n9763) );
  INVX1 U5258 ( .A(n9763), .Y(n5300) );
  AND2X1 U5259 ( .A(n6076), .B(n5993), .Y(n6434) );
  INVX1 U5260 ( .A(n6434), .Y(n5301) );
  AND2X1 U5261 ( .A(n6076), .B(n5277), .Y(n6460) );
  INVX1 U5262 ( .A(n6460), .Y(n5302) );
  AND2X1 U5263 ( .A(n6085), .B(n7850), .Y(n7851) );
  INVX1 U5264 ( .A(n7851), .Y(n5303) );
  AND2X1 U5265 ( .A(n3161), .B(n5776), .Y(n6476) );
  INVX1 U5266 ( .A(n6476), .Y(n5304) );
  AND2X1 U5267 ( .A(n3129), .B(n5776), .Y(n8524) );
  INVX1 U5268 ( .A(n8524), .Y(n5305) );
  INVX1 U5269 ( .A(mult32_B[1]), .Y(n5306) );
  AND2X1 U5270 ( .A(n6076), .B(n6319), .Y(n6440) );
  INVX1 U5271 ( .A(n6440), .Y(n5307) );
  AND2X1 U5272 ( .A(n6076), .B(n6042), .Y(n6462) );
  INVX1 U5273 ( .A(n6462), .Y(n5308) );
  BUFX2 U5274 ( .A(n6545), .Y(n5309) );
  AND2X1 U5275 ( .A(n6085), .B(n8087), .Y(n8088) );
  INVX1 U5276 ( .A(n8088), .Y(n5310) );
  AND2X1 U5277 ( .A(n3163), .B(n5776), .Y(n6622) );
  INVX1 U5278 ( .A(n6622), .Y(n5311) );
  AND2X1 U5279 ( .A(n3132), .B(n5776), .Y(n8734) );
  INVX1 U5280 ( .A(n8734), .Y(n5312) );
  AND2X1 U5281 ( .A(n6076), .B(n6018), .Y(n6448) );
  INVX1 U5282 ( .A(n6448), .Y(n5313) );
  AND2X1 U5283 ( .A(n6076), .B(n6034), .Y(n6459) );
  INVX1 U5284 ( .A(n6459), .Y(n5314) );
  INVX1 U5285 ( .A(n10479), .Y(n5315) );
  BUFX2 U5286 ( .A(n6825), .Y(n5316) );
  BUFX2 U5287 ( .A(n6901), .Y(n5317) );
  AND2X1 U5288 ( .A(n6085), .B(n8858), .Y(n8859) );
  INVX1 U5289 ( .A(n8859), .Y(n5318) );
  AND2X1 U5290 ( .A(n3164), .B(n5776), .Y(n6700) );
  INVX1 U5291 ( .A(n6700), .Y(n5319) );
  AND2X1 U5292 ( .A(n3133), .B(n5776), .Y(n8797) );
  INVX1 U5293 ( .A(n8797), .Y(n5320) );
  AND2X1 U5294 ( .A(n530), .B(n5773), .Y(n7131) );
  INVX1 U5295 ( .A(n7131), .Y(n5321) );
  BUFX2 U5296 ( .A(n7132), .Y(n5322) );
  AND2X1 U5297 ( .A(n6076), .B(n5286), .Y(n6447) );
  INVX1 U5298 ( .A(n6447), .Y(n5323) );
  AND2X1 U5299 ( .A(n6076), .B(n6356), .Y(n6468) );
  INVX1 U5300 ( .A(n6468), .Y(n5324) );
  BUFX2 U5301 ( .A(n8927), .Y(n5325) );
  AND2X1 U5302 ( .A(n6085), .B(n9099), .Y(n9100) );
  INVX1 U5303 ( .A(n9100), .Y(n5326) );
  AND2X1 U5304 ( .A(n3166), .B(n5776), .Y(n6824) );
  INVX1 U5305 ( .A(n6824), .Y(n5327) );
  AND2X1 U5306 ( .A(n3134), .B(n5776), .Y(n8849) );
  INVX1 U5307 ( .A(n8849), .Y(n5328) );
  AND2X1 U5308 ( .A(n527), .B(n5773), .Y(n6951) );
  INVX1 U5309 ( .A(n6951), .Y(n5329) );
  BUFX2 U5310 ( .A(n6952), .Y(n5330) );
  AND2X1 U5311 ( .A(n415), .B(n5778), .Y(n7483) );
  INVX1 U5312 ( .A(n7483), .Y(n5331) );
  AND2X1 U5313 ( .A(n6076), .B(n6061), .Y(n6469) );
  INVX1 U5314 ( .A(n6469), .Y(n5332) );
  AND2X1 U5315 ( .A(n6076), .B(n6026), .Y(n6453) );
  INVX1 U5316 ( .A(n6453), .Y(n5333) );
  BUFX2 U5317 ( .A(n7135), .Y(n5334) );
  BUFX2 U5318 ( .A(n9032), .Y(n5335) );
  AND2X1 U5319 ( .A(n6085), .B(n6801), .Y(n6802) );
  INVX1 U5320 ( .A(n6802), .Y(n5336) );
  BUFX2 U5321 ( .A(n7698), .Y(n5337) );
  AND2X1 U5322 ( .A(n6085), .B(n9894), .Y(n9895) );
  INVX1 U5323 ( .A(n9895), .Y(n5338) );
  AND2X1 U5324 ( .A(n1310), .B(n6125), .Y(n6751) );
  INVX1 U5325 ( .A(n6751), .Y(n5339) );
  AND2X1 U5326 ( .A(n3169), .B(n5776), .Y(n7007) );
  INVX1 U5327 ( .A(n7007), .Y(n5340) );
  AND2X1 U5328 ( .A(n3136), .B(n5776), .Y(n8982) );
  INVX1 U5329 ( .A(n8982), .Y(n5341) );
  BUFX2 U5330 ( .A(n7115), .Y(n5342) );
  BUFX2 U5331 ( .A(n9293), .Y(n5343) );
  AND2X1 U5332 ( .A(n531), .B(n5773), .Y(n7206) );
  INVX1 U5333 ( .A(n7206), .Y(n5344) );
  BUFX2 U5334 ( .A(n7207), .Y(n5345) );
  INVX1 U5335 ( .A(n8592), .Y(n5346) );
  INVX1 U5336 ( .A(n6435), .Y(n5347) );
  AND2X1 U5337 ( .A(n6076), .B(n6354), .Y(n6467) );
  INVX1 U5338 ( .A(n6467), .Y(n5348) );
  BUFX2 U5339 ( .A(n7338), .Y(n5349) );
  BUFX2 U5340 ( .A(n8776), .Y(n5350) );
  BUFX2 U5341 ( .A(n9090), .Y(n5351) );
  BUFX2 U5342 ( .A(n9655), .Y(n5352) );
  AND2X1 U5343 ( .A(n6085), .B(n7178), .Y(n7179) );
  INVX1 U5344 ( .A(n7179), .Y(n5353) );
  AND2X1 U5345 ( .A(n3177), .B(n5776), .Y(n7520) );
  INVX1 U5346 ( .A(n7520), .Y(n5354) );
  AND2X1 U5347 ( .A(n3170), .B(n5776), .Y(n7064) );
  INVX1 U5348 ( .A(n7064), .Y(n5355) );
  AND2X1 U5349 ( .A(n3137), .B(n5776), .Y(n9031) );
  INVX1 U5350 ( .A(n9031), .Y(n5356) );
  BUFX2 U5351 ( .A(n9896), .Y(n5357) );
  BUFX2 U5352 ( .A(n6817), .Y(n5358) );
  BUFX2 U5353 ( .A(n9600), .Y(n5359) );
  BUFX2 U5354 ( .A(n6750), .Y(n5360) );
  AND2X1 U5355 ( .A(n5841), .B(n5821), .Y(n6627) );
  INVX1 U5356 ( .A(n6627), .Y(n5361) );
  AND2X1 U5357 ( .A(n5840), .B(n6497), .Y(n6570) );
  INVX1 U5358 ( .A(n6570), .Y(n5362) );
  AND2X1 U5359 ( .A(n7490), .B(n5834), .Y(n7298) );
  INVX1 U5360 ( .A(n7298), .Y(n5363) );
  AND2X1 U5361 ( .A(n5875), .B(n5874), .Y(n7491) );
  INVX1 U5362 ( .A(n7491), .Y(n5364) );
  AND2X1 U5363 ( .A(n1570), .B(n6123), .Y(n6932) );
  INVX1 U5364 ( .A(n6932), .Y(n5365) );
  BUFX2 U5365 ( .A(n6933), .Y(n5366) );
  AND2X1 U5366 ( .A(n9183), .B(n10491), .Y(n9184) );
  INVX1 U5367 ( .A(n9184), .Y(n5367) );
  AND2X1 U5368 ( .A(n775), .B(n5825), .Y(n9424) );
  INVX1 U5369 ( .A(n9424), .Y(n5368) );
  INVX1 U5370 ( .A(n6446), .Y(n5369) );
  AND2X1 U5371 ( .A(n6076), .B(n21), .Y(n6464) );
  INVX1 U5372 ( .A(n6464), .Y(n5370) );
  BUFX2 U5373 ( .A(n9165), .Y(n5371) );
  BUFX2 U5374 ( .A(n9810), .Y(n5372) );
  BUFX2 U5375 ( .A(n9306), .Y(n5373) );
  BUFX2 U5376 ( .A(n7210), .Y(n5374) );
  BUFX2 U5377 ( .A(n9733), .Y(n5375) );
  AND2X1 U5378 ( .A(n6085), .B(n8195), .Y(n8196) );
  INVX1 U5379 ( .A(n8196), .Y(n5376) );
  BUFX2 U5380 ( .A(n8832), .Y(n5377) );
  AND2X1 U5381 ( .A(n3178), .B(n5776), .Y(n7579) );
  INVX1 U5382 ( .A(n7579), .Y(n5378) );
  AND2X1 U5383 ( .A(n1285), .B(n6125), .Y(n9219) );
  INVX1 U5384 ( .A(n9219), .Y(n5379) );
  AND2X1 U5385 ( .A(n3171), .B(n5776), .Y(n7134) );
  INVX1 U5386 ( .A(n7134), .Y(n5380) );
  AND2X1 U5387 ( .A(n3138), .B(n5776), .Y(n9089) );
  INVX1 U5388 ( .A(n9089), .Y(n5381) );
  BUFX2 U5389 ( .A(n10112), .Y(n5382) );
  BUFX2 U5390 ( .A(n8082), .Y(n5383) );
  AND2X1 U5391 ( .A(n1102), .B(n6127), .Y(n6804) );
  INVX1 U5392 ( .A(n6804), .Y(n5384) );
  BUFX2 U5393 ( .A(n6543), .Y(n5385) );
  BUFX2 U5394 ( .A(n6880), .Y(n5386) );
  BUFX2 U5395 ( .A(n7572), .Y(n5387) );
  BUFX2 U5396 ( .A(n10008), .Y(n5388) );
  BUFX2 U5397 ( .A(n6748), .Y(n5389) );
  BUFX2 U5398 ( .A(n6828), .Y(n5390) );
  AND2X1 U5399 ( .A(n1087), .B(n6127), .Y(n9897) );
  INVX1 U5400 ( .A(n9897), .Y(n5391) );
  AND2X1 U5401 ( .A(n5813), .B(n6490), .Y(n6431) );
  INVX1 U5402 ( .A(n6431), .Y(n5392) );
  AND2X1 U5403 ( .A(n6557), .B(n7222), .Y(n6625) );
  INVX1 U5404 ( .A(n6625), .Y(n5393) );
  AND2X1 U5405 ( .A(n5798), .B(n5821), .Y(n8679) );
  INVX1 U5406 ( .A(n8679), .Y(n5394) );
  BUFX2 U5407 ( .A(n8600), .Y(n5395) );
  INVX1 U5408 ( .A(n8599), .Y(n5396) );
  INVX1 U5409 ( .A(n10356), .Y(n5397) );
  INVX1 U5410 ( .A(n9324), .Y(n5398) );
  BUFX2 U5411 ( .A(n10372), .Y(n5399) );
  AND2X1 U5412 ( .A(n6497), .B(n5874), .Y(n7490) );
  INVX1 U5413 ( .A(n7490), .Y(n5400) );
  INVX1 U5414 ( .A(mult32_B[7]), .Y(n5401) );
  INVX1 U5415 ( .A(mult32_B[19]), .Y(n5402) );
  INVX1 U5416 ( .A(mult32_B[18]), .Y(n5403) );
  INVX1 U5417 ( .A(mult32_B[20]), .Y(n5404) );
  INVX1 U5418 ( .A(mult32_B[23]), .Y(n5405) );
  AND2X1 U5419 ( .A(n3834), .B(n5775), .Y(n8471) );
  INVX1 U5420 ( .A(n8471), .Y(n5406) );
  AND2X1 U5421 ( .A(n399), .B(n5778), .Y(n8491) );
  INVX1 U5422 ( .A(n8491), .Y(n5407) );
  BUFX2 U5423 ( .A(n7923), .Y(n5408) );
  AND2X1 U5424 ( .A(n6076), .B(n6337), .Y(n6449) );
  INVX1 U5425 ( .A(n6449), .Y(n5409) );
  AND2X1 U5426 ( .A(n6076), .B(n6345), .Y(n6461) );
  INVX1 U5427 ( .A(n6461), .Y(n5410) );
  AND2X1 U5428 ( .A(n776), .B(n5825), .Y(n9534) );
  INVX1 U5429 ( .A(n9534), .Y(n5411) );
  BUFX2 U5430 ( .A(n7403), .Y(n5412) );
  BUFX2 U5431 ( .A(n6936), .Y(n5413) );
  BUFX2 U5432 ( .A(n8669), .Y(n5414) );
  BUFX2 U5433 ( .A(n10323), .Y(n5415) );
  BUFX2 U5434 ( .A(n7281), .Y(n5416) );
  BUFX2 U5435 ( .A(n6955), .Y(n5417) );
  BUFX2 U5436 ( .A(n9239), .Y(n5418) );
  BUFX2 U5437 ( .A(n6669), .Y(n5419) );
  AND2X1 U5438 ( .A(n6085), .B(n9206), .Y(n9207) );
  INVX1 U5439 ( .A(n9207), .Y(n5420) );
  BUFX2 U5440 ( .A(n6898), .Y(n5421) );
  AND2X1 U5441 ( .A(n6085), .B(n6895), .Y(n6896) );
  INVX1 U5442 ( .A(n6896), .Y(n5422) );
  BUFX2 U5443 ( .A(n6991), .Y(n5423) );
  BUFX2 U5444 ( .A(n10077), .Y(n5424) );
  AND2X1 U5445 ( .A(n3179), .B(n5776), .Y(n7653) );
  INVX1 U5446 ( .A(n7653), .Y(n5425) );
  AND2X1 U5447 ( .A(n1312), .B(n6125), .Y(n6829) );
  INVX1 U5448 ( .A(n6829), .Y(n5426) );
  AND2X1 U5449 ( .A(n3172), .B(n5776), .Y(n7209) );
  INVX1 U5450 ( .A(n7209), .Y(n5427) );
  AND2X1 U5451 ( .A(n3139), .B(n5776), .Y(n9164) );
  INVX1 U5452 ( .A(n9164), .Y(n5428) );
  OR2X1 U5453 ( .A(n5574), .B(n5505), .Y(n10488) );
  INVX1 U5454 ( .A(n10488), .Y(n5429) );
  BUFX2 U5455 ( .A(n9428), .Y(n5430) );
  AND2X1 U5456 ( .A(n1325), .B(n5848), .Y(n8652) );
  INVX1 U5457 ( .A(n8652), .Y(n5431) );
  BUFX2 U5458 ( .A(n9218), .Y(n5432) );
  BUFX2 U5459 ( .A(n8636), .Y(n5433) );
  BUFX2 U5460 ( .A(n10122), .Y(n5434) );
  AND2X1 U5461 ( .A(n811), .B(n5857), .Y(n8655) );
  BUFX2 U5462 ( .A(n9093), .Y(n5435) );
  BUFX2 U5463 ( .A(n7513), .Y(n5436) );
  BUFX2 U5464 ( .A(n9540), .Y(n5437) );
  BUFX2 U5465 ( .A(n8777), .Y(n5438) );
  AND2X1 U5466 ( .A(n1119), .B(n5826), .Y(n7853) );
  INVX1 U5467 ( .A(n7853), .Y(n5439) );
  AND2X1 U5468 ( .A(n6153), .B(n6152), .Y(n9688) );
  AND2X1 U5469 ( .A(n5813), .B(n5812), .Y(n6430) );
  INVX1 U5470 ( .A(n6430), .Y(n5440) );
  INVX1 U5471 ( .A(n9046), .Y(n5441) );
  AND2X1 U5472 ( .A(n5821), .B(n5794), .Y(n9689) );
  INVX1 U5473 ( .A(n9689), .Y(n5442) );
  BUFX4 U5474 ( .A(oprB[28]), .Y(n5882) );
  AND2X1 U5475 ( .A(n5819), .B(n6206), .Y(n8300) );
  INVX1 U5476 ( .A(n8300), .Y(n5443) );
  AND2X1 U5477 ( .A(n6189), .B(n7491), .Y(n8314) );
  INVX1 U5478 ( .A(n8314), .Y(n5444) );
  AND2X1 U5479 ( .A(n10167), .B(n9647), .Y(n9767) );
  INVX1 U5480 ( .A(n9767), .Y(n5445) );
  AND2X1 U5481 ( .A(n5833), .B(n6557), .Y(n7172) );
  INVX1 U5482 ( .A(n7172), .Y(n5446) );
  OR2X1 U5483 ( .A(shift_amount[3]), .B(n6635), .Y(n6918) );
  INVX1 U5484 ( .A(n6918), .Y(n5447) );
  OR2X1 U5485 ( .A(shift_amount[3]), .B(n9718), .Y(n9976) );
  INVX1 U5486 ( .A(n9976), .Y(n5448) );
  AND2X1 U5487 ( .A(n5840), .B(n5850), .Y(n7146) );
  INVX1 U5488 ( .A(n7146), .Y(n5449) );
  INVX1 U5489 ( .A(n9310), .Y(n5450) );
  INVX1 U5490 ( .A(n6505), .Y(n5451) );
  BUFX2 U5491 ( .A(n9326), .Y(n5452) );
  INVX1 U5492 ( .A(mult32_B[2]), .Y(n5453) );
  INVX1 U5493 ( .A(mult32_B[5]), .Y(n5454) );
  INVX1 U5494 ( .A(mult32_B[27]), .Y(n5455) );
  INVX1 U5495 ( .A(mult32_B[15]), .Y(n5456) );
  AND2X2 U5496 ( .A(n191), .B(n1178), .Y(mult32_B[16]) );
  INVX1 U5497 ( .A(mult32_B[16]), .Y(n5457) );
  INVX1 U5498 ( .A(mult32_B[26]), .Y(n5458) );
  INVX1 U5499 ( .A(mult32_B[24]), .Y(n5459) );
  BUFX2 U5500 ( .A(n10413), .Y(n5461) );
  AND2X1 U5501 ( .A(n517), .B(n5773), .Y(n10412) );
  INVX1 U5502 ( .A(n10412), .Y(n5462) );
  BUFX2 U5503 ( .A(n8351), .Y(n5463) );
  AND2X1 U5504 ( .A(n549), .B(n6143), .Y(n8350) );
  INVX1 U5505 ( .A(n8350), .Y(n5464) );
  AND2X1 U5506 ( .A(n5788), .B(n6332), .Y(n9050) );
  INVX1 U5507 ( .A(n9050), .Y(n5465) );
  AND2X1 U5508 ( .A(n5952), .B(n9632), .Y(n7590) );
  INVX1 U5509 ( .A(n7590), .Y(n5466) );
  AND2X1 U5510 ( .A(n6076), .B(n6325), .Y(n6442) );
  INVX1 U5511 ( .A(n6442), .Y(n5467) );
  INVX1 U5512 ( .A(n10353), .Y(n5468) );
  BUFX2 U5513 ( .A(n10348), .Y(n5469) );
  BUFX2 U5514 ( .A(n10347), .Y(n5470) );
  BUFX2 U5515 ( .A(n7252), .Y(n5471) );
  BUFX2 U5516 ( .A(n9862), .Y(n5472) );
  BUFX2 U5517 ( .A(n7276), .Y(n5473) );
  BUFX2 U5518 ( .A(n9301), .Y(n5474) );
  OR2X1 U5519 ( .A(n7102), .B(n10315), .Y(n7103) );
  INVX1 U5520 ( .A(n7103), .Y(n5475) );
  BUFX2 U5521 ( .A(n7623), .Y(n5476) );
  AND2X1 U5522 ( .A(n6085), .B(n10139), .Y(n10140) );
  INVX1 U5523 ( .A(n10140), .Y(n5477) );
  BUFX2 U5524 ( .A(n8924), .Y(n5478) );
  AND2X1 U5525 ( .A(n6085), .B(n8921), .Y(n8922) );
  INVX1 U5526 ( .A(n8922), .Y(n5479) );
  OR2X1 U5527 ( .A(n9846), .B(n6284), .Y(n7073) );
  INVX1 U5528 ( .A(n7073), .Y(n5480) );
  AND2X1 U5529 ( .A(n3180), .B(n5776), .Y(n7728) );
  INVX1 U5530 ( .A(n7728), .Y(n5481) );
  AND2X1 U5531 ( .A(n799), .B(n5825), .Y(n6900) );
  INVX1 U5532 ( .A(n6900), .Y(n5482) );
  BUFX2 U5533 ( .A(n7768), .Y(n5483) );
  AND2X1 U5534 ( .A(n1264), .B(n5785), .Y(n9890) );
  INVX1 U5535 ( .A(n9890), .Y(n5484) );
  AND2X1 U5536 ( .A(n3174), .B(n5776), .Y(n7337) );
  INVX1 U5537 ( .A(n7337), .Y(n5485) );
  AND2X1 U5538 ( .A(n3140), .B(n5776), .Y(n9238) );
  INVX1 U5539 ( .A(n9238), .Y(n5486) );
  AND2X1 U5540 ( .A(n2284), .B(n5838), .Y(n9962) );
  BUFX2 U5541 ( .A(n6992), .Y(n5487) );
  BUFX2 U5542 ( .A(n9778), .Y(n5488) );
  BUFX2 U5543 ( .A(n9586), .Y(n5489) );
  BUFX2 U5544 ( .A(n8671), .Y(n5490) );
  BUFX2 U5545 ( .A(n7288), .Y(n5491) );
  BUFX2 U5546 ( .A(n10134), .Y(n5492) );
  BUFX2 U5547 ( .A(n9314), .Y(n5493) );
  AND2X1 U5548 ( .A(n1103), .B(n5826), .Y(n6836) );
  INVX1 U5549 ( .A(n6836), .Y(n5494) );
  AND2X1 U5550 ( .A(n907), .B(n6133), .Y(n8710) );
  INVX1 U5551 ( .A(n8710), .Y(n5495) );
  BUFX2 U5552 ( .A(n6799), .Y(n5496) );
  BUFX2 U5553 ( .A(n9756), .Y(n5497) );
  BUFX2 U5554 ( .A(n10271), .Y(n5498) );
  BUFX2 U5555 ( .A(n8825), .Y(n5499) );
  BUFX2 U5556 ( .A(n9063), .Y(n5500) );
  AND2X1 U5557 ( .A(n7804), .B(n6189), .Y(n8035) );
  INVX1 U5558 ( .A(n8035), .Y(n5501) );
  AND2X1 U5559 ( .A(n6782), .B(n5900), .Y(n7022) );
  INVX1 U5560 ( .A(n7022), .Y(n5502) );
  AND2X1 U5561 ( .A(n5799), .B(n5821), .Y(n7656) );
  INVX1 U5562 ( .A(n7656), .Y(n5503) );
  AND2X1 U5563 ( .A(n6791), .B(n6083), .Y(n6590) );
  INVX1 U5564 ( .A(n6590), .Y(n5504) );
  INVX1 U5565 ( .A(n10486), .Y(n5505) );
  AND2X1 U5566 ( .A(n9127), .B(n9647), .Y(n8738) );
  INVX1 U5567 ( .A(n8738), .Y(n5506) );
  AND2X1 U5568 ( .A(n7491), .B(n6657), .Y(n6926) );
  INVX1 U5569 ( .A(n6926), .Y(n5507) );
  AND2X1 U5570 ( .A(n5852), .B(n5874), .Y(n6557) );
  INVX1 U5571 ( .A(n6557), .Y(n5508) );
  OR2X1 U5572 ( .A(shift_amount[3]), .B(n8697), .Y(n8944) );
  INVX1 U5573 ( .A(n8944), .Y(n5509) );
  INVX1 U5574 ( .A(mult32_A[31]), .Y(n5510) );
  AND2X1 U5575 ( .A(n5911), .B(n5730), .Y(n6432) );
  INVX1 U5576 ( .A(n6432), .Y(n5511) );
  AND2X1 U5577 ( .A(n6076), .B(n5880), .Y(n6433) );
  INVX1 U5578 ( .A(n6433), .Y(n5512) );
  INVX1 U5579 ( .A(n10355), .Y(n5513) );
  AND2X1 U5580 ( .A(n6202), .B(n6204), .Y(n8299) );
  INVX1 U5581 ( .A(n8299), .Y(n5514) );
  INVX1 U5582 ( .A(n7148), .Y(n5515) );
  BUFX2 U5583 ( .A(n6634), .Y(n5516) );
  BUFX2 U5584 ( .A(n6633), .Y(n5517) );
  BUFX2 U5585 ( .A(n8316), .Y(n5518) );
  AND2X1 U5586 ( .A(n5840), .B(n5851), .Y(n9500) );
  INVX1 U5587 ( .A(n9500), .Y(n5519) );
  INVX1 U5588 ( .A(n8968), .Y(n5520) );
  INVX1 U5589 ( .A(mult32_B[8]), .Y(n5521) );
  INVX1 U5590 ( .A(mult32_B[22]), .Y(n5522) );
  INVX1 U5591 ( .A(mult32_B[25]), .Y(n5523) );
  AND2X1 U5592 ( .A(n1538), .B(n5779), .Y(n8959) );
  INVX1 U5593 ( .A(n8959), .Y(n5524) );
  BUFX2 U5594 ( .A(n8960), .Y(n5525) );
  AND2X1 U5595 ( .A(n5765), .B(n10290), .Y(n10374) );
  INVX1 U5596 ( .A(n10374), .Y(n5526) );
  BUFX2 U5597 ( .A(n9968), .Y(n5527) );
  AND2X1 U5598 ( .A(n59), .B(n6077), .Y(n9618) );
  INVX1 U5599 ( .A(n9618), .Y(n5528) );
  AND2X1 U5600 ( .A(n6076), .B(n6330), .Y(n6444) );
  INVX1 U5601 ( .A(n6444), .Y(n5529) );
  BUFX2 U5602 ( .A(n9364), .Y(n5530) );
  BUFX2 U5603 ( .A(n7913), .Y(n5531) );
  BUFX2 U5604 ( .A(n9096), .Y(n5532) );
  BUFX2 U5605 ( .A(n10103), .Y(n5533) );
  BUFX2 U5606 ( .A(n6769), .Y(n5534) );
  BUFX2 U5607 ( .A(n7469), .Y(n5535) );
  BUFX2 U5608 ( .A(n10067), .Y(n5536) );
  OR2X1 U5609 ( .A(n9273), .B(n10315), .Y(n9274) );
  INVX1 U5610 ( .A(n9274), .Y(n5537) );
  BUFX2 U5611 ( .A(n6592), .Y(n5538) );
  AND2X1 U5612 ( .A(n6085), .B(n7919), .Y(n7920) );
  INVX1 U5613 ( .A(n7920), .Y(n5539) );
  BUFX2 U5614 ( .A(n7048), .Y(n5540) );
  BUFX2 U5615 ( .A(n7769), .Y(n5541) );
  AND2X1 U5616 ( .A(n1356), .B(n5772), .Y(n6544) );
  INVX1 U5617 ( .A(n6544), .Y(n5542) );
  AND2X1 U5618 ( .A(n3185), .B(n5776), .Y(n8020) );
  INVX1 U5619 ( .A(n8020), .Y(n5543) );
  AND2X1 U5620 ( .A(n763), .B(n5825), .Y(n8668) );
  INVX1 U5621 ( .A(n8668), .Y(n5544) );
  AND2X1 U5622 ( .A(n1011), .B(n6129), .Y(n10135) );
  INVX1 U5623 ( .A(n10135), .Y(n5545) );
  AND2X1 U5624 ( .A(n1269), .B(n6125), .Y(n10259) );
  INVX1 U5625 ( .A(n10259), .Y(n5546) );
  BUFX2 U5626 ( .A(n8775), .Y(n5547) );
  AND2X1 U5627 ( .A(n3173), .B(n5776), .Y(n7275) );
  INVX1 U5628 ( .A(n7275), .Y(n5548) );
  AND2X1 U5629 ( .A(n3141), .B(n5776), .Y(n9300) );
  INVX1 U5630 ( .A(n9300), .Y(n5549) );
  BUFX2 U5631 ( .A(n10322), .Y(n5550) );
  BUFX2 U5632 ( .A(n9015), .Y(n5551) );
  BUFX2 U5633 ( .A(n7279), .Y(n5552) );
  BUFX2 U5634 ( .A(n10141), .Y(n5553) );
  BUFX2 U5635 ( .A(n8659), .Y(n5554) );
  BUFX2 U5636 ( .A(n9861), .Y(n5555) );
  BUFX2 U5637 ( .A(n7000), .Y(n5556) );
  BUFX2 U5638 ( .A(n6680), .Y(n5557) );
  BUFX2 U5639 ( .A(n9231), .Y(n5558) );
  BUFX2 U5640 ( .A(n7251), .Y(n5559) );
  AND2X1 U5641 ( .A(n1110), .B(n6127), .Y(n7289) );
  INVX1 U5642 ( .A(n7289), .Y(n5560) );
  AND2X1 U5643 ( .A(n1078), .B(n6127), .Y(n9315) );
  INVX1 U5644 ( .A(n9315), .Y(n5561) );
  AND2X1 U5645 ( .A(n6556), .B(n6155), .Y(n6626) );
  INVX1 U5646 ( .A(n6626), .Y(n5562) );
  AND2X1 U5647 ( .A(n5747), .B(n7284), .Y(n7339) );
  INVX1 U5648 ( .A(n7339), .Y(n5563) );
  AND2X1 U5649 ( .A(n5821), .B(n6192), .Y(n7804) );
  INVX1 U5650 ( .A(n7804), .Y(n5564) );
  INVX1 U5651 ( .A(oprB[44]), .Y(n6192) );
  INVX1 U5652 ( .A(n9109), .Y(n5565) );
  BUFX2 U5653 ( .A(n6565), .Y(n5566) );
  OR2X1 U5654 ( .A(n6064), .B(n5943), .Y(n6564) );
  INVX1 U5655 ( .A(n6564), .Y(n5567) );
  INVX1 U5656 ( .A(n7285), .Y(n5568) );
  AND2X1 U5657 ( .A(n8115), .B(n9647), .Y(n7732) );
  INVX1 U5658 ( .A(n7732), .Y(n5569) );
  AND2X1 U5659 ( .A(n7491), .B(n8691), .Y(n8952) );
  INVX1 U5660 ( .A(n8952), .Y(n5570) );
  INVX1 U5661 ( .A(n9127), .Y(n5571) );
  INVX1 U5662 ( .A(n6579), .Y(n5572) );
  OR2X1 U5663 ( .A(shift_amount[3]), .B(n7683), .Y(n7930) );
  INVX1 U5664 ( .A(n7930), .Y(n5573) );
  AND2X2 U5665 ( .A(n5573), .B(n6155), .Y(n5861) );
  AND2X1 U5666 ( .A(n5853), .B(n5874), .Y(n10487) );
  INVX1 U5667 ( .A(n10487), .Y(n5574) );
  INVX8 U5668 ( .A(n6219), .Y(n5907) );
  INVX1 U5669 ( .A(mult32_A[12]), .Y(n5575) );
  AND2X1 U5670 ( .A(n5961), .B(n5730), .Y(n6455) );
  INVX1 U5671 ( .A(n6455), .Y(n5576) );
  AND2X1 U5672 ( .A(n6076), .B(n6032), .Y(n6456) );
  INVX1 U5673 ( .A(n6456), .Y(n5577) );
  AND2X1 U5674 ( .A(n7490), .B(n5833), .Y(n8954) );
  INVX1 U5675 ( .A(n8954), .Y(n5578) );
  INVX1 U5676 ( .A(n9187), .Y(n5579) );
  BUFX2 U5677 ( .A(n8695), .Y(n5580) );
  BUFX2 U5678 ( .A(n8696), .Y(n5581) );
  BUFX2 U5679 ( .A(n7300), .Y(n5582) );
  AND2X1 U5680 ( .A(n5851), .B(n5869), .Y(n8910) );
  INVX1 U5681 ( .A(n8910), .Y(n5583) );
  INVX1 U5682 ( .A(n10226), .Y(n5584) );
  BUFX2 U5683 ( .A(n9717), .Y(n5585) );
  BUFX2 U5684 ( .A(n9716), .Y(n5586) );
  INVX1 U5685 ( .A(n6791), .Y(n5587) );
  AND2X1 U5686 ( .A(n5840), .B(n5875), .Y(n10290) );
  INVX1 U5687 ( .A(n10290), .Y(n5588) );
  AND2X1 U5688 ( .A(n5656), .B(n9846), .Y(n10104) );
  INVX1 U5689 ( .A(n10104), .Y(n5589) );
  AND2X2 U5690 ( .A(n194), .B(n1182), .Y(mult32_B[11]) );
  AND2X1 U5691 ( .A(n5720), .B(n5871), .Y(n10564) );
  INVX1 U5692 ( .A(mult32_B[4]), .Y(n5591) );
  INVX1 U5693 ( .A(mult32_B[12]), .Y(n5592) );
  AND2X1 U5694 ( .A(n5813), .B(n5814), .Y(n6363) );
  AND2X1 U5695 ( .A(n3208), .B(n5827), .Y(n7470) );
  INVX1 U5696 ( .A(n7470), .Y(n5594) );
  AND2X1 U5697 ( .A(n5792), .B(n5937), .Y(n7026) );
  INVX1 U5698 ( .A(n7026), .Y(n5595) );
  AND2X1 U5699 ( .A(n5787), .B(n6301), .Y(n8039) );
  INVX1 U5700 ( .A(n8039), .Y(n5596) );
  AND2X1 U5701 ( .A(n5793), .B(n6049), .Y(n10088) );
  INVX1 U5702 ( .A(n10088), .Y(n5597) );
  AND2X1 U5703 ( .A(n5912), .B(n6077), .Y(n6555) );
  INVX1 U5704 ( .A(n6555), .Y(n5598) );
  AND2X1 U5705 ( .A(n6076), .B(n6004), .Y(n6443) );
  INVX1 U5706 ( .A(n6443), .Y(n5599) );
  AND2X1 U5707 ( .A(n2276), .B(n5838), .Y(n9429) );
  INVX1 U5708 ( .A(n9429), .Y(n5600) );
  BUFX2 U5709 ( .A(n8963), .Y(n5601) );
  BUFX2 U5710 ( .A(n9491), .Y(n5602) );
  BUFX2 U5711 ( .A(n8625), .Y(n5603) );
  AND2X1 U5712 ( .A(n6085), .B(n6833), .Y(n6834) );
  INVX1 U5713 ( .A(n6834), .Y(n5604) );
  AND2X1 U5714 ( .A(n6085), .B(n10246), .Y(n10247) );
  INVX1 U5715 ( .A(n10247), .Y(n5605) );
  AND2X1 U5716 ( .A(n1795), .B(n5777), .Y(n6935) );
  INVX1 U5717 ( .A(n6935), .Y(n5606) );
  AND2X1 U5718 ( .A(n767), .B(n5825), .Y(n8926) );
  INVX1 U5719 ( .A(n8926), .Y(n5607) );
  AND2X1 U5720 ( .A(n1043), .B(n6129), .Y(n8083) );
  INVX1 U5721 ( .A(n8083), .Y(n5608) );
  AND2X1 U5722 ( .A(n1747), .B(n5777), .Y(n9957) );
  INVX1 U5723 ( .A(n9957), .Y(n5609) );
  AND2X1 U5724 ( .A(n1062), .B(n5786), .Y(n7280) );
  INVX1 U5725 ( .A(n7280), .Y(n5610) );
  BUFX2 U5726 ( .A(n9809), .Y(n5611) );
  AND2X1 U5727 ( .A(n1296), .B(n5785), .Y(n7846) );
  INVX1 U5728 ( .A(n7846), .Y(n5612) );
  AND2X1 U5729 ( .A(n3804), .B(n6108), .Y(n6615) );
  INVX1 U5730 ( .A(n6615), .Y(n5613) );
  AND2X1 U5731 ( .A(n3168), .B(n5776), .Y(n6954) );
  INVX1 U5732 ( .A(n6954), .Y(n5614) );
  AND2X1 U5733 ( .A(n3175), .B(n5776), .Y(n7402) );
  INVX1 U5734 ( .A(n7402), .Y(n5615) );
  AND2X1 U5735 ( .A(n3142), .B(n5776), .Y(n9363) );
  INVX1 U5736 ( .A(n9363), .Y(n5616) );
  BUFX2 U5737 ( .A(n8005), .Y(n5617) );
  BUFX2 U5738 ( .A(n9072), .Y(n5618) );
  BUFX2 U5739 ( .A(n9928), .Y(n5619) );
  BUFX2 U5740 ( .A(n6903), .Y(n5620) );
  BUFX2 U5741 ( .A(n7911), .Y(n5621) );
  BUFX2 U5742 ( .A(n9094), .Y(n5622) );
  BUFX2 U5743 ( .A(n9304), .Y(n5623) );
  BUFX2 U5744 ( .A(n8448), .Y(n5624) );
  BUFX2 U5745 ( .A(n10102), .Y(n5625) );
  BUFX2 U5746 ( .A(n10256), .Y(n5626) );
  BUFX2 U5747 ( .A(n6678), .Y(n5627) );
  INVX1 U5748 ( .A(n6071), .Y(n5628) );
  AND2X1 U5749 ( .A(n6347), .B(n6083), .Y(n10182) );
  INVX1 U5750 ( .A(n10182), .Y(n5629) );
  AND2X1 U5751 ( .A(n6189), .B(n10290), .Y(n7748) );
  INVX1 U5752 ( .A(n7748), .Y(n5630) );
  AND2X1 U5753 ( .A(n5900), .B(n10290), .Y(n6723) );
  INVX1 U5754 ( .A(n6723), .Y(n5631) );
  AND2X1 U5755 ( .A(n5883), .B(n5821), .Y(n9371) );
  INVX1 U5756 ( .A(n9371), .Y(n5632) );
  BUFX2 U5757 ( .A(n7598), .Y(n5633) );
  OR2X1 U5758 ( .A(n6064), .B(n6307), .Y(n7597) );
  INVX1 U5759 ( .A(n7597), .Y(n5634) );
  INVX1 U5760 ( .A(n9996), .Y(n5635) );
  AND2X1 U5761 ( .A(n7491), .B(n7686), .Y(n7946) );
  INVX1 U5762 ( .A(n7946), .Y(n5636) );
  INVX1 U5763 ( .A(n9309), .Y(n5637) );
  AND2X1 U5764 ( .A(n6170), .B(n6172), .Y(n7284) );
  INVX1 U5765 ( .A(n7284), .Y(n5638) );
  INVX1 U5766 ( .A(n8876), .Y(n5639) );
  OR2X1 U5767 ( .A(n5896), .B(n6546), .Y(n6851) );
  INVX1 U5768 ( .A(n6851), .Y(n5640) );
  INVX1 U5769 ( .A(n6913), .Y(n5641) );
  INVX1 U5770 ( .A(n8939), .Y(n5642) );
  BUFX2 U5771 ( .A(n6515), .Y(n5643) );
  INVX1 U5772 ( .A(n5643), .Y(n6499) );
  AND2X1 U5773 ( .A(n6731), .B(n6557), .Y(n8485) );
  INVX1 U5774 ( .A(n8485), .Y(n5644) );
  INVX1 U5775 ( .A(mult32_A[15]), .Y(n5645) );
  AND2X1 U5776 ( .A(n5952), .B(n5730), .Y(n6451) );
  INVX1 U5777 ( .A(n6451), .Y(n5646) );
  AND2X1 U5778 ( .A(n6076), .B(n59), .Y(n6452) );
  INVX1 U5779 ( .A(n6452), .Y(n5647) );
  OR2X1 U5780 ( .A(shift_amount[3]), .B(n7678), .Y(n7933) );
  INVX1 U5781 ( .A(n7933), .Y(n5648) );
  OR2X1 U5782 ( .A(shift_amount[3]), .B(n9711), .Y(n9979) );
  INVX1 U5783 ( .A(n9979), .Y(n5649) );
  AND2X1 U5784 ( .A(n10290), .B(n6160), .Y(n6920) );
  INVX1 U5785 ( .A(n6920), .Y(n5650) );
  INVX1 U5786 ( .A(n8176), .Y(n5651) );
  BUFX2 U5787 ( .A(n7663), .Y(n5652) );
  BUFX2 U5788 ( .A(n7664), .Y(n5653) );
  INVX1 U5789 ( .A(n10371), .Y(n5654) );
  INVX1 U5790 ( .A(n9774), .Y(n5655) );
  AND2X1 U5791 ( .A(n5851), .B(n5874), .Y(n9969) );
  AND2X1 U5792 ( .A(n5840), .B(n5853), .Y(n10291) );
  INVX1 U5793 ( .A(n10291), .Y(n5656) );
  AND2X2 U5794 ( .A(n196), .B(n1184), .Y(mult32_B[9]) );
  INVX1 U5795 ( .A(mult32_B[3]), .Y(n5658) );
  AND2X2 U5796 ( .A(n80), .B(n1187), .Y(mult32_B[6]) );
  INVX1 U5797 ( .A(mult32_B[6]), .Y(n5659) );
  INVX1 U5798 ( .A(mult32_B[10]), .Y(n5660) );
  INVX1 U5799 ( .A(mult32_B[13]), .Y(n5661) );
  AND2X1 U5800 ( .A(n5813), .B(n5815), .Y(n6361) );
  INVX1 U5801 ( .A(mult32_B[28]), .Y(n5662) );
  INVX1 U5802 ( .A(mult32_B[17]), .Y(n5663) );
  INVX1 U5803 ( .A(mult32_B[21]), .Y(n5664) );
  INVX1 U5804 ( .A(mult32_B[29]), .Y(n5665) );
  AND2X1 U5805 ( .A(n3224), .B(n5827), .Y(n8477) );
  INVX1 U5806 ( .A(n8477), .Y(n5666) );
  AND2X1 U5807 ( .A(n2585), .B(n5831), .Y(n8657) );
  INVX1 U5808 ( .A(n8657), .Y(n5667) );
  AND2X1 U5809 ( .A(n3452), .B(n5847), .Y(n8672) );
  INVX1 U5810 ( .A(n8672), .Y(n5668) );
  INVX1 U5811 ( .A(n10567), .Y(n5669) );
  AND2X1 U5812 ( .A(n3898), .B(n5828), .Y(n10565) );
  INVX1 U5813 ( .A(n10565), .Y(n5670) );
  BUFX2 U5814 ( .A(n10566), .Y(n5671) );
  OR2X1 U5815 ( .A(n10316), .B(n10315), .Y(n10317) );
  INVX1 U5816 ( .A(n10317), .Y(n5672) );
  AND2X1 U5817 ( .A(n6085), .B(n9964), .Y(n9965) );
  INVX1 U5818 ( .A(n9965), .Y(n5673) );
  AND2X1 U5819 ( .A(n3153), .B(n5776), .Y(n10066) );
  INVX1 U5820 ( .A(n10066), .Y(n5674) );
  AND2X1 U5821 ( .A(n1763), .B(n5777), .Y(n8962) );
  INVX1 U5822 ( .A(n8962), .Y(n5675) );
  AND2X1 U5823 ( .A(n1779), .B(n5777), .Y(n7912) );
  INVX1 U5824 ( .A(n7912), .Y(n5676) );
  AND2X1 U5825 ( .A(n1027), .B(n5786), .Y(n9095) );
  INVX1 U5826 ( .A(n9095), .Y(n5677) );
  AND2X1 U5827 ( .A(n1280), .B(n6125), .Y(n8854) );
  INVX1 U5828 ( .A(n8854), .Y(n5678) );
  AND2X1 U5829 ( .A(n3165), .B(n5776), .Y(n6768) );
  INVX1 U5830 ( .A(n6768), .Y(n5679) );
  AND2X1 U5831 ( .A(n3176), .B(n5776), .Y(n7468) );
  INVX1 U5832 ( .A(n7468), .Y(n5680) );
  AND2X1 U5833 ( .A(n3772), .B(n6108), .Y(n8648) );
  INVX1 U5834 ( .A(n8648), .Y(n5681) );
  AND2X1 U5835 ( .A(n3144), .B(n5776), .Y(n9490) );
  INVX1 U5836 ( .A(n9490), .Y(n5682) );
  AND2X1 U5837 ( .A(n3544), .B(n5830), .Y(n8449) );
  INVX1 U5838 ( .A(n8449), .Y(n5683) );
  AND2X1 U5839 ( .A(n1030), .B(n6129), .Y(n9305) );
  INVX1 U5840 ( .A(n9305), .Y(n5684) );
  AND2X1 U5841 ( .A(n1290), .B(n5785), .Y(n9531) );
  INVX1 U5842 ( .A(n9531), .Y(n5685) );
  AND2X1 U5843 ( .A(n808), .B(n5825), .Y(n7507) );
  INVX1 U5844 ( .A(n7507), .Y(n5686) );
  BUFX2 U5845 ( .A(n8929), .Y(n5687) );
  BUFX2 U5846 ( .A(n8863), .Y(n5688) );
  AND2X1 U5847 ( .A(n1578), .B(n6123), .Y(n7450) );
  INVX1 U5848 ( .A(n7450), .Y(n5689) );
  BUFX2 U5849 ( .A(n8454), .Y(n5690) );
  BUFX2 U5850 ( .A(n9430), .Y(n5691) );
  BUFX2 U5851 ( .A(n9216), .Y(n5692) );
  BUFX2 U5852 ( .A(n10258), .Y(n5693) );
  AND2X1 U5853 ( .A(n1091), .B(n6127), .Y(n10142) );
  INVX1 U5854 ( .A(n10142), .Y(n5694) );
  AND2X1 U5855 ( .A(n6790), .B(n6083), .Y(n9731) );
  INVX1 U5856 ( .A(n9731), .Y(n5695) );
  AND2X1 U5857 ( .A(n9845), .B(n6245), .Y(n10082) );
  INVX1 U5858 ( .A(n10082), .Y(n5696) );
  AND2X1 U5859 ( .A(n5840), .B(n5852), .Y(n6556) );
  INVX1 U5860 ( .A(n6556), .Y(n5697) );
  INVX1 U5861 ( .A(n9498), .Y(n5698) );
  AND2X1 U5862 ( .A(n6189), .B(n6192), .Y(n8115) );
  INVX1 U5863 ( .A(n8115), .Y(n5699) );
  AND2X1 U5864 ( .A(n5858), .B(n9647), .Y(n6704) );
  INVX1 U5865 ( .A(n6704), .Y(n5700) );
  AND2X1 U5866 ( .A(n8999), .B(n5821), .Y(n9460) );
  INVX1 U5867 ( .A(n9460), .Y(n5701) );
  AND2X1 U5868 ( .A(n7491), .B(n9720), .Y(n9992) );
  INVX1 U5869 ( .A(n9992), .Y(n5702) );
  INVX1 U5870 ( .A(n10167), .Y(n5703) );
  INVX1 U5871 ( .A(n7405), .Y(n5704) );
  INVX1 U5872 ( .A(n7869), .Y(n5705) );
  INVX1 U5873 ( .A(n9913), .Y(n5706) );
  AND2X1 U5874 ( .A(n7687), .B(n6188), .Y(n7950) );
  INVX1 U5875 ( .A(n7950), .Y(n5707) );
  INVX1 U5876 ( .A(n9474), .Y(n5708) );
  OR2X1 U5877 ( .A(n6203), .B(n8158), .Y(n8414) );
  INVX1 U5878 ( .A(n8414), .Y(n5709) );
  INVX1 U5879 ( .A(n10507), .Y(n5710) );
  AND2X1 U5880 ( .A(n5908), .B(n10290), .Y(n8755) );
  INVX1 U5881 ( .A(n8755), .Y(n5711) );
  INVX1 U5882 ( .A(n8368), .Y(n5712) );
  INVX1 U5883 ( .A(n10430), .Y(n5713) );
  INVX1 U5884 ( .A(n9378), .Y(n5714) );
  AND2X1 U5885 ( .A(n6155), .B(n6157), .Y(n7222) );
  INVX1 U5886 ( .A(n7222), .Y(n5715) );
  OR2X1 U5887 ( .A(shift_amount[3]), .B(n6650), .Y(n6938) );
  INVX1 U5888 ( .A(n6938), .Y(n5716) );
  OR2X1 U5889 ( .A(shift_amount[3]), .B(n8715), .Y(n8965) );
  INVX1 U5890 ( .A(n8965), .Y(n5717) );
  INVX1 U5891 ( .A(n7352), .Y(n5718) );
  AND2X1 U5892 ( .A(n6570), .B(n5889), .Y(n10375) );
  INVX1 U5893 ( .A(n10375), .Y(n5719) );
  OR2X1 U5894 ( .A(op[3]), .B(op[2]), .Y(n7984) );
  INVX1 U5895 ( .A(n7984), .Y(n5720) );
  AND2X1 U5896 ( .A(n5834), .B(n6557), .Y(n10500) );
  INVX1 U5897 ( .A(n10500), .Y(n5721) );
  AND2X1 U5898 ( .A(n8910), .B(n6142), .Y(n10480) );
  INVX1 U5899 ( .A(n10480), .Y(n5722) );
  AND2X1 U5900 ( .A(n5851), .B(n5872), .Y(n10502) );
  INVX1 U5901 ( .A(n10216), .Y(n5723) );
  AND2X1 U5902 ( .A(n9688), .B(n6625), .Y(n9576) );
  INVX1 U5903 ( .A(n9576), .Y(n5724) );
  INVX1 U5904 ( .A(n7167), .Y(n5725) );
  AND2X1 U5905 ( .A(n6203), .B(n6201), .Y(n8163) );
  INVX1 U5906 ( .A(n8163), .Y(n5726) );
  INVX1 U5907 ( .A(n9175), .Y(n5727) );
  INVX1 U5908 ( .A(n9803), .Y(n5728) );
  AND2X1 U5909 ( .A(shift_amount[3]), .B(n6152), .Y(n9626) );
  AND2X1 U5910 ( .A(n5886), .B(n6153), .Y(n9632) );
  AND2X1 U5911 ( .A(n7490), .B(n6156), .Y(n10085) );
  INVX1 U5912 ( .A(n10085), .Y(n5729) );
  INVX1 U5913 ( .A(n6457), .Y(n5730) );
  AND2X1 U5914 ( .A(n5850), .B(n5874), .Y(n9629) );
  INVX1 U5915 ( .A(n9629), .Y(n5731) );
  AND2X1 U5916 ( .A(n9688), .B(n6626), .Y(n10354) );
  INVX1 U5917 ( .A(n10354), .Y(n5732) );
  INVX1 U5918 ( .A(n10093), .Y(n5733) );
  INVX2 U5919 ( .A(n6291), .Y(n5947) );
  INVX2 U5920 ( .A(n5971), .Y(n5974) );
  INVX2 U5921 ( .A(n6302), .Y(n5977) );
  INVX8 U5922 ( .A(n6258), .Y(n6257) );
  INVX8 U5923 ( .A(n6238), .Y(n6237) );
  INVX8 U5924 ( .A(n6270), .Y(n6269) );
  INVX2 U5925 ( .A(n6176), .Y(n6175) );
  INVX8 U5926 ( .A(n5884), .Y(n5885) );
  INVX2 U5927 ( .A(oprA[0]), .Y(n6359) );
  INVX2 U5928 ( .A(n6293), .Y(n5955) );
  INVX1 U5929 ( .A(oprB[13]), .Y(n6246) );
  INVX1 U5930 ( .A(n6335), .Y(n6015) );
  INVX1 U5931 ( .A(n6307), .Y(n5985) );
  INVX8 U5932 ( .A(n6040), .Y(n6041) );
  INVX2 U5933 ( .A(n5971), .Y(n5972) );
  INVX2 U5934 ( .A(oprB[12]), .Y(n6248) );
  INVX1 U5935 ( .A(n6062), .Y(n6080) );
  INVX1 U5936 ( .A(n6062), .Y(n6079) );
  AND2X1 U5937 ( .A(n8485), .B(n9688), .Y(n5735) );
  INVX1 U5938 ( .A(n6084), .Y(n6083) );
  INVX1 U5939 ( .A(n4717), .Y(n7418) );
  INVX1 U5940 ( .A(n5722), .Y(n6112) );
  INVX1 U5941 ( .A(n5440), .Y(n6074) );
  INVX1 U5942 ( .A(n5392), .Y(n6075) );
  INVX1 U5943 ( .A(n9793), .Y(n9703) );
  INVX1 U5944 ( .A(n5452), .Y(n9258) );
  INVX1 U5945 ( .A(n5582), .Y(n7233) );
  INVX1 U5946 ( .A(n5518), .Y(n8247) );
  INVX1 U5947 ( .A(n9185), .Y(n9461) );
  INVX1 U5948 ( .A(n5399), .Y(n10300) );
  BUFX2 U5949 ( .A(n5695), .Y(n6069) );
  INVX1 U5950 ( .A(n8174), .Y(n8426) );
  BUFX2 U5951 ( .A(n5695), .Y(n6070) );
  INVX1 U5952 ( .A(n10224), .Y(n10506) );
  INVX1 U5953 ( .A(n4847), .Y(n10447) );
  INVX1 U5954 ( .A(n4846), .Y(n7369) );
  INVX1 U5955 ( .A(n7413), .Y(n7371) );
  INVX1 U5956 ( .A(n10518), .Y(n10449) );
  INVX1 U5957 ( .A(n5042), .Y(n9375) );
  INVX1 U5958 ( .A(n9688), .Y(n6084) );
  INVX1 U5959 ( .A(n6095), .Y(n6094) );
  INVX1 U5960 ( .A(n6099), .Y(n6098) );
  INVX1 U5961 ( .A(n6078), .Y(n6077) );
  INVX1 U5962 ( .A(n6144), .Y(n6143) );
  INVX1 U5963 ( .A(n4808), .Y(n6705) );
  INVX1 U5964 ( .A(n6109), .Y(n6108) );
  INVX1 U5965 ( .A(n6118), .Y(n6117) );
  INVX1 U5966 ( .A(n6120), .Y(n6119) );
  INVX1 U5967 ( .A(n6111), .Y(n6110) );
  INVX1 U5968 ( .A(n6126), .Y(n6125) );
  INVX1 U5969 ( .A(n6146), .Y(n6145) );
  INVX1 U5970 ( .A(n6107), .Y(n6106) );
  AND2X1 U5971 ( .A(n5907), .B(n10291), .Y(n5737) );
  INVX1 U5972 ( .A(n6148), .Y(n6147) );
  INVX1 U5973 ( .A(n6140), .Y(n6139) );
  INVX1 U5974 ( .A(n6122), .Y(n6121) );
  INVX1 U5975 ( .A(n6124), .Y(n6123) );
  INVX1 U5976 ( .A(n6116), .Y(n6115) );
  INVX1 U5977 ( .A(n6150), .Y(n6149) );
  INVX1 U5978 ( .A(n6130), .Y(n6129) );
  INVX1 U5979 ( .A(n10522), .Y(n6088) );
  INVX1 U5980 ( .A(n6082), .Y(n6081) );
  INVX1 U5981 ( .A(n6036), .Y(n6038) );
  BUFX2 U5982 ( .A(oprB[28]), .Y(n5883) );
  BUFX2 U5983 ( .A(oprA[31]), .Y(n5879) );
  BUFX2 U5984 ( .A(n5990), .Y(n5880) );
  INVX1 U5985 ( .A(n6358), .Y(n6058) );
  INVX1 U5986 ( .A(n6338), .Y(n6022) );
  INVX1 U5987 ( .A(n6429), .Y(n6076) );
  INVX1 U5988 ( .A(n6846), .Y(n6847) );
  INVX1 U5989 ( .A(n7150), .Y(n6636) );
  INVX1 U5990 ( .A(n10489), .Y(n10376) );
  INVX1 U5991 ( .A(n6921), .Y(n6656) );
  INVX1 U5992 ( .A(n5739), .Y(n10574) );
  INVX1 U5993 ( .A(n6480), .Y(n6498) );
  INVX1 U5994 ( .A(n8877), .Y(n9372) );
  INVX1 U5995 ( .A(n8698), .Y(n9183) );
  INVX1 U5996 ( .A(n7870), .Y(n8363) );
  INVX1 U5997 ( .A(n6732), .Y(n9791) );
  INVX1 U5998 ( .A(n10505), .Y(n7428) );
  INVX1 U5999 ( .A(n10491), .Y(n7408) );
  INVX1 U6000 ( .A(n8966), .Y(n8721) );
  INVX1 U6001 ( .A(n8996), .Y(n8683) );
  INVX1 U6002 ( .A(n4815), .Y(n8739) );
  INVX1 U6003 ( .A(n9969), .Y(n6095) );
  INVX1 U6004 ( .A(n10502), .Y(n6099) );
  INVX1 U6005 ( .A(n7427), .Y(n7140) );
  INVX1 U6006 ( .A(n9632), .Y(n6078) );
  INVX1 U6007 ( .A(n9626), .Y(n6082) );
  INVX1 U6008 ( .A(n6789), .Y(n10383) );
  INVX1 U6009 ( .A(n8553), .Y(n9441) );
  INVX1 U6010 ( .A(n7549), .Y(n8433) );
  INVX1 U6011 ( .A(n5772), .Y(n6140) );
  INVX1 U6012 ( .A(n5774), .Y(n6107) );
  INVX1 U6013 ( .A(n5775), .Y(n6109) );
  INVX1 U6014 ( .A(n5771), .Y(n6146) );
  INVX1 U6015 ( .A(n5777), .Y(n6122) );
  INVX1 U6016 ( .A(n5778), .Y(n6118) );
  INVX1 U6017 ( .A(n5790), .Y(n6120) );
  INVX1 U6018 ( .A(n5779), .Y(n6124) );
  INVX1 U6019 ( .A(n5780), .Y(n6111) );
  INVX1 U6020 ( .A(n5781), .Y(n6116) );
  INVX1 U6021 ( .A(n5784), .Y(n6148) );
  INVX1 U6022 ( .A(n5783), .Y(n6150) );
  INVX1 U6023 ( .A(n5786), .Y(n6130) );
  INVX1 U6024 ( .A(n5785), .Y(n6126) );
  AND2X1 U6025 ( .A(n6517), .B(n5911), .Y(n5743) );
  AND2X1 U6026 ( .A(n7550), .B(n5952), .Y(n5744) );
  AND2X1 U6027 ( .A(n6173), .B(n10290), .Y(n5745) );
  AND2X1 U6028 ( .A(n9577), .B(n59), .Y(n5746) );
  AND2X1 U6029 ( .A(n6205), .B(n5819), .Y(n5748) );
  INVX1 U6030 ( .A(n4650), .Y(n7404) );
  INVX1 U6031 ( .A(n4623), .Y(n8881) );
  INVX1 U6032 ( .A(n4621), .Y(n7875) );
  INVX1 U6033 ( .A(n4619), .Y(n6856) );
  INVX1 U6034 ( .A(n8301), .Y(n8435) );
  INVX1 U6035 ( .A(n4624), .Y(n8883) );
  INVX1 U6036 ( .A(n4620), .Y(n6858) );
  INVX1 U6037 ( .A(n4626), .Y(n9922) );
  INVX1 U6038 ( .A(n4622), .Y(n7877) );
  AND2X1 U6039 ( .A(n6626), .B(n9632), .Y(n5749) );
  INVX1 U6040 ( .A(n9311), .Y(n9443) );
  AND2X1 U6041 ( .A(n5800), .B(n6626), .Y(n5750) );
  AND2X1 U6042 ( .A(n9626), .B(n6626), .Y(n5751) );
  INVX1 U6043 ( .A(n6105), .Y(n6104) );
  INVX1 U6044 ( .A(n6101), .Y(n6100) );
  INVX1 U6045 ( .A(n6136), .Y(n6135) );
  INVX1 U6046 ( .A(n6128), .Y(n6127) );
  AND2X1 U6047 ( .A(n8999), .B(n9647), .Y(n5752) );
  AND2X1 U6048 ( .A(n6974), .B(n9647), .Y(n5753) );
  AND2X1 U6049 ( .A(n10034), .B(n9647), .Y(n5754) );
  AND2X1 U6050 ( .A(n7988), .B(n9647), .Y(n5755) );
  INVX1 U6051 ( .A(n7612), .Y(n7874) );
  INVX1 U6052 ( .A(n9696), .Y(n9977) );
  INVX1 U6053 ( .A(n6138), .Y(n6137) );
  INVX1 U6054 ( .A(n7677), .Y(n7932) );
  INVX1 U6055 ( .A(n6649), .Y(n6937) );
  INVX1 U6056 ( .A(n8718), .Y(n8964) );
  INVX1 U6057 ( .A(n9710), .Y(n9978) );
  INVX1 U6058 ( .A(n6087), .Y(n6086) );
  INVX1 U6059 ( .A(n9914), .Y(n10425) );
  INVX1 U6060 ( .A(n6852), .Y(n7346) );
  INVX1 U6061 ( .A(n7524), .Y(n7538) );
  INVX1 U6062 ( .A(n8528), .Y(n8542) );
  INVX1 U6063 ( .A(n9551), .Y(n9565) );
  AND2X1 U6064 ( .A(n10291), .B(n6245), .Y(n5757) );
  INVX1 U6065 ( .A(n6134), .Y(n6133) );
  INVX1 U6066 ( .A(n6132), .Y(n6131) );
  INVX1 U6067 ( .A(n6097), .Y(n6096) );
  INVX1 U6068 ( .A(n6093), .Y(n6092) );
  AND2X1 U6069 ( .A(n5899), .B(n10291), .Y(n5758) );
  INVX1 U6070 ( .A(n9719), .Y(n10222) );
  INVX1 U6071 ( .A(n7684), .Y(n8172) );
  INVX1 U6072 ( .A(n9169), .Y(n9473) );
  INVX1 U6073 ( .A(n8157), .Y(n8413) );
  INVX1 U6074 ( .A(n7685), .Y(n7931) );
  INVX1 U6075 ( .A(n10209), .Y(n10495) );
  AND2X1 U6076 ( .A(n6189), .B(n10291), .Y(n5759) );
  INVX1 U6077 ( .A(n6103), .Y(n6102) );
  INVX1 U6078 ( .A(n6722), .Y(n7224) );
  INVX1 U6079 ( .A(n5801), .Y(n6073) );
  INVX1 U6080 ( .A(n5773), .Y(n6144) );
  AND2X1 U6081 ( .A(n7284), .B(n5934), .Y(n5760) );
  INVX1 U6082 ( .A(n5800), .Y(n6062) );
  INVX1 U6083 ( .A(n6114), .Y(n6113) );
  INVX1 U6084 ( .A(n5782), .Y(n6114) );
  AND2X1 U6085 ( .A(n5899), .B(n7491), .Y(n5763) );
  AND2X1 U6086 ( .A(n6173), .B(n10291), .Y(n5764) );
  INVX1 U6087 ( .A(n6091), .Y(n6090) );
  INVX1 U6088 ( .A(n10564), .Y(n6089) );
  INVX1 U6089 ( .A(n6190), .Y(n6189) );
  INVX1 U6090 ( .A(n5996), .Y(n5997) );
  INVX1 U6091 ( .A(n6044), .Y(n6046) );
  INVX1 U6092 ( .A(n6306), .Y(n5981) );
  INVX1 U6093 ( .A(n6353), .Y(n6055) );
  INVX1 U6094 ( .A(n6346), .Y(n6039) );
  INVX1 U6095 ( .A(n6283), .Y(n5928) );
  INVX1 U6096 ( .A(n6300), .Y(n5975) );
  INVX1 U6097 ( .A(n6), .Y(n6047) );
  INVX1 U6098 ( .A(n6010), .Y(n6012) );
  INVX1 U6099 ( .A(n6161), .Y(n5901) );
  INVX1 U6100 ( .A(n6040), .Y(n6042) );
  INVX1 U6101 ( .A(n6358), .Y(n6356) );
  INVX1 U6102 ( .A(n5894), .Y(n5895) );
  INVX1 U6103 ( .A(n5891), .Y(n5892) );
  INVX1 U6104 ( .A(n5894), .Y(n5896) );
  INVX1 U6105 ( .A(n6331), .Y(n6330) );
  INVX1 U6106 ( .A(n6162), .Y(n5905) );
  INVX1 U6107 ( .A(n6162), .Y(n5906) );
  INVX1 U6108 ( .A(n6162), .Y(n5904) );
  INVX1 U6109 ( .A(op[0]), .Y(n6142) );
  INVX1 U6110 ( .A(n6324), .Y(n6322) );
  INVX1 U6111 ( .A(n6323), .Y(n6321) );
  INVX1 U6112 ( .A(oprA[17]), .Y(n6020) );
  INVX1 U6113 ( .A(n6291), .Y(n5946) );
  INVX1 U6114 ( .A(n10441), .Y(n9630) );
  INVX1 U6115 ( .A(n9389), .Y(n8602) );
  INVX1 U6116 ( .A(n8379), .Y(n7600) );
  INVX1 U6117 ( .A(n7363), .Y(n6567) );
  INVX1 U6118 ( .A(n8871), .Y(n8872) );
  INVX1 U6119 ( .A(n7864), .Y(n7865) );
  BUFX2 U6120 ( .A(n9795), .Y(n6065) );
  BUFX2 U6121 ( .A(n9797), .Y(n6066) );
  INVX1 U6122 ( .A(n5766), .Y(n9647) );
  INVX1 U6123 ( .A(n7080), .Y(n7075) );
  AND2X1 U6124 ( .A(n9629), .B(n6156), .Y(n5770) );
  INVX1 U6125 ( .A(n10155), .Y(n10439) );
  AND2X1 U6126 ( .A(n5857), .B(n6141), .Y(n5771) );
  AND2X1 U6127 ( .A(n5848), .B(n6141), .Y(n5772) );
  AND2X1 U6128 ( .A(n5849), .B(n6141), .Y(n5773) );
  AND2X1 U6129 ( .A(n5847), .B(n6141), .Y(n5774) );
  AND2X1 U6130 ( .A(n5845), .B(n6141), .Y(n5775) );
  AND2X1 U6131 ( .A(n5844), .B(n6141), .Y(n5776) );
  AND2X1 U6132 ( .A(n5840), .B(n5812), .Y(n5777) );
  AND2X1 U6133 ( .A(n5840), .B(n5855), .Y(n5778) );
  AND2X1 U6134 ( .A(n5840), .B(n5815), .Y(n5779) );
  AND2X1 U6135 ( .A(n5835), .B(n6142), .Y(n5780) );
  AND2X1 U6136 ( .A(n5856), .B(n6142), .Y(n5781) );
  AND2X1 U6137 ( .A(n5843), .B(n6142), .Y(n5782) );
  AND2X1 U6138 ( .A(n5842), .B(n6142), .Y(n5783) );
  AND2X1 U6139 ( .A(n5846), .B(n6142), .Y(n5784) );
  AND2X1 U6140 ( .A(n6490), .B(n5840), .Y(n5785) );
  AND2X1 U6141 ( .A(n5814), .B(n5840), .Y(n5786) );
  INVX1 U6142 ( .A(n9179), .Y(n8700) );
  INVX1 U6143 ( .A(n8376), .Y(n8116) );
  AND2X1 U6144 ( .A(n6203), .B(n6202), .Y(n5787) );
  INVX1 U6145 ( .A(n6152), .Y(n5886) );
  INVX1 U6146 ( .A(n6973), .Y(n10033) );
  AND2X1 U6147 ( .A(n8939), .B(n6219), .Y(n5789) );
  AND2X1 U6148 ( .A(n5840), .B(n5854), .Y(n5790) );
  INVX1 U6149 ( .A(n6152), .Y(n5887) );
  AND2X1 U6150 ( .A(n6156), .B(n6557), .Y(n5791) );
  INVX1 U6151 ( .A(n6155), .Y(n5890) );
  AND2X1 U6152 ( .A(n6974), .B(n5821), .Y(n5795) );
  BUFX2 U6153 ( .A(n6084), .Y(n6064) );
  BUFX2 U6154 ( .A(n6084), .Y(n6063) );
  AND2X1 U6155 ( .A(n7988), .B(n5821), .Y(n5796) );
  AND2X1 U6156 ( .A(n10034), .B(n5821), .Y(n5797) );
  AND2X1 U6157 ( .A(n6190), .B(n6192), .Y(n5799) );
  AND2X1 U6158 ( .A(shift_amount[3]), .B(n5888), .Y(n5800) );
  INVX1 U6159 ( .A(n5967), .Y(n6296) );
  INVX1 U6160 ( .A(n9386), .Y(n9128) );
  INVX1 U6161 ( .A(n6152), .Y(n5888) );
  INVX1 U6162 ( .A(n10438), .Y(n10168) );
  INVX1 U6163 ( .A(n6287), .Y(n6286) );
  INVX1 U6164 ( .A(n5823), .Y(n6136) );
  INVX1 U6165 ( .A(n5824), .Y(n6134) );
  INVX1 U6166 ( .A(n5825), .Y(n6138) );
  INVX1 U6167 ( .A(n5839), .Y(n6132) );
  INVX1 U6168 ( .A(n5828), .Y(n6097) );
  INVX1 U6169 ( .A(n5829), .Y(n6087) );
  INVX1 U6170 ( .A(n5830), .Y(n6093) );
  INVX1 U6171 ( .A(n5827), .Y(n6101) );
  INVX1 U6172 ( .A(n5831), .Y(n6103) );
  INVX1 U6173 ( .A(n5838), .Y(n6105) );
  INVX1 U6174 ( .A(n4625), .Y(n9919) );
  INVX1 U6175 ( .A(n5818), .Y(n6091) );
  INVX1 U6176 ( .A(n4653), .Y(n8415) );
  INVX1 U6177 ( .A(n6309), .Y(n6308) );
  INVX1 U6178 ( .A(n6580), .Y(n6855) );
  INVX1 U6179 ( .A(n8604), .Y(n8882) );
  INVX1 U6180 ( .A(n8611), .Y(n8880) );
  INVX1 U6181 ( .A(n9633), .Y(n9921) );
  INVX1 U6182 ( .A(n6569), .Y(n6857) );
  INVX1 U6183 ( .A(n9640), .Y(n9920) );
  AND2X1 U6184 ( .A(n7755), .B(n5821), .Y(n5802) );
  INVX1 U6185 ( .A(n7602), .Y(n7876) );
  AND2X1 U6186 ( .A(n6733), .B(n5821), .Y(n5803) );
  AND2X1 U6187 ( .A(n9792), .B(n5821), .Y(n5804) );
  INVX1 U6188 ( .A(n7142), .Y(n7430) );
  INVX1 U6189 ( .A(n9115), .Y(n9387) );
  INVX1 U6190 ( .A(n7071), .Y(n7361) );
  INVX1 U6191 ( .A(n8103), .Y(n8377) );
  INVX1 U6192 ( .A(n6067), .Y(n6068) );
  AND2X1 U6193 ( .A(n8762), .B(n5821), .Y(n5805) );
  INVX1 U6194 ( .A(n9908), .Y(n9909) );
  INVX1 U6195 ( .A(n5826), .Y(n6128) );
  INVX1 U6196 ( .A(n8106), .Y(n8375) );
  INVX1 U6197 ( .A(n9118), .Y(n9385) );
  AND2X1 U6198 ( .A(n7950), .B(n6190), .Y(n5806) );
  AND2X1 U6199 ( .A(n6579), .B(n67), .Y(n5807) );
  AND2X1 U6200 ( .A(n5903), .B(n5821), .Y(n5808) );
  AND2X1 U6201 ( .A(n8610), .B(n43), .Y(n5809) );
  AND2X1 U6202 ( .A(n7611), .B(n5964), .Y(n5810) );
  AND2X1 U6203 ( .A(n5885), .B(n9639), .Y(n5811) );
  INVX1 U6204 ( .A(n10315), .Y(n6085) );
  INVX1 U6205 ( .A(n6280), .Y(n6279) );
  INVX1 U6206 ( .A(op[0]), .Y(n6141) );
  INVX1 U6207 ( .A(oprB[35]), .Y(n6210) );
  INVX1 U6208 ( .A(n6355), .Y(n6354) );
  INVX1 U6209 ( .A(oprB[51]), .Y(n6178) );
  INVX1 U6210 ( .A(oprB[50]), .Y(n6180) );
  INVX1 U6211 ( .A(oprB[52]), .Y(n6176) );
  INVX1 U6212 ( .A(oprB[49]), .Y(n6182) );
  INVX1 U6213 ( .A(oprB[18]), .Y(n6238) );
  INVX2 U6214 ( .A(n6168), .Y(n6167) );
  INVX1 U6215 ( .A(oprB[56]), .Y(n6168) );
  INVX1 U6216 ( .A(oprB[41]), .Y(n6198) );
  INVX1 U6217 ( .A(oprB[40]), .Y(n6200) );
  INVX1 U6218 ( .A(oprB[42]), .Y(n6196) );
  INVX1 U6219 ( .A(oprB[8]), .Y(n6256) );
  INVX1 U6220 ( .A(oprB[9]), .Y(n6254) );
  INVX1 U6221 ( .A(oprB[48]), .Y(n6184) );
  INVX1 U6222 ( .A(n6458), .Y(mult32_A[11]) );
  INVX1 U6223 ( .A(oprB[43]), .Y(n6194) );
  AND2X1 U6224 ( .A(n5870), .B(n5868), .Y(n5812) );
  INVX1 U6225 ( .A(oprB[46]), .Y(n6188) );
  INVX1 U6226 ( .A(oprB[47]), .Y(n6186) );
  INVX1 U6227 ( .A(oprB[57]), .Y(n6166) );
  INVX1 U6228 ( .A(oprB[54]), .Y(n6172) );
  AND2X1 U6229 ( .A(n5869), .B(n6142), .Y(n5813) );
  AND2X1 U6230 ( .A(n5816), .B(n5868), .Y(n5814) );
  AND2X1 U6231 ( .A(n5871), .B(n5868), .Y(n5815) );
  INVX1 U6232 ( .A(n6364), .Y(n6490) );
  INVX1 U6233 ( .A(oprA[39]), .Y(n5971) );
  AND2X1 U6234 ( .A(n5817), .B(n6516), .Y(n5816) );
  INVX1 U6235 ( .A(n6346), .Y(n6345) );
  INVX1 U6236 ( .A(n6326), .Y(n6325) );
  AND2X1 U6237 ( .A(n6362), .B(n6471), .Y(n5817) );
  INVX1 U6238 ( .A(oprB[61]), .Y(n5898) );
  INVX1 U6239 ( .A(oprA[16]), .Y(n6023) );
  INVX1 U6240 ( .A(oprB[59]), .Y(n6162) );
  INVX1 U6241 ( .A(oprB[62]), .Y(n5894) );
  INVX1 U6242 ( .A(n6318), .Y(n6317) );
  INVX1 U6243 ( .A(oprA[6]), .Y(n6044) );
  INVX1 U6244 ( .A(n6157), .Y(n6156) );
  AND2X1 U6245 ( .A(n5840), .B(n5876), .Y(n5819) );
  INVX1 U6246 ( .A(n5819), .Y(n9846) );
  AND2X1 U6247 ( .A(n5896), .B(n6158), .Y(n5820) );
  AND2X1 U6248 ( .A(n5876), .B(n5874), .Y(n5821) );
  AND2X1 U6249 ( .A(n7146), .B(n6155), .Y(n5822) );
  AND2X1 U6250 ( .A(n5872), .B(n5855), .Y(n5823) );
  AND2X1 U6251 ( .A(n5872), .B(n5854), .Y(n5824) );
  AND2X1 U6252 ( .A(n5854), .B(n5874), .Y(n5825) );
  AND2X1 U6253 ( .A(n5814), .B(n5874), .Y(n5826) );
  INVX1 U6254 ( .A(n6298), .Y(n6297) );
  AND2X1 U6255 ( .A(n5850), .B(n5872), .Y(n5827) );
  AND2X1 U6256 ( .A(n6497), .B(n5872), .Y(n5828) );
  AND2X1 U6257 ( .A(n5853), .B(n5872), .Y(n5829) );
  AND2X1 U6258 ( .A(n5875), .B(n5872), .Y(n5830) );
  AND2X1 U6259 ( .A(n5852), .B(n5872), .Y(n5831) );
  AND2X1 U6260 ( .A(n5816), .B(n5877), .Y(n5832) );
  INVX1 U6261 ( .A(n5832), .Y(n10522) );
  AND2X1 U6262 ( .A(n6156), .B(n6155), .Y(n5833) );
  AND2X1 U6263 ( .A(n5889), .B(n6157), .Y(n5834) );
  AND2X1 U6264 ( .A(n5853), .B(n5869), .Y(n5835) );
  AND2X1 U6265 ( .A(n9908), .B(n6155), .Y(n5836) );
  AND2X1 U6266 ( .A(n8871), .B(n6155), .Y(n5837) );
  AND2X1 U6267 ( .A(n5876), .B(n5872), .Y(n5838) );
  AND2X1 U6268 ( .A(n5855), .B(n5874), .Y(n5839) );
  AND2X1 U6269 ( .A(n6489), .B(n6488), .Y(n5840) );
  INVX1 U6270 ( .A(n10517), .Y(n6067) );
  AND2X1 U6271 ( .A(n5874), .B(n5812), .Y(n5842) );
  AND2X1 U6272 ( .A(n5876), .B(n5869), .Y(n5843) );
  AND2X1 U6273 ( .A(n5850), .B(n5869), .Y(n5844) );
  AND2X1 U6274 ( .A(n6497), .B(n5869), .Y(n5845) );
  AND2X1 U6275 ( .A(n5815), .B(n5874), .Y(n5846) );
  AND2X1 U6276 ( .A(n5875), .B(n5869), .Y(n5847) );
  AND2X1 U6277 ( .A(n6490), .B(n5874), .Y(n5848) );
  AND2X1 U6278 ( .A(n5869), .B(n5855), .Y(n5849) );
  AND2X1 U6279 ( .A(n5866), .B(n6471), .Y(n5850) );
  AND2X1 U6280 ( .A(n5873), .B(n5816), .Y(n5851) );
  AND2X1 U6281 ( .A(n5873), .B(n5871), .Y(n5852) );
  AND2X1 U6282 ( .A(n5873), .B(n5870), .Y(n5853) );
  AND2X1 U6283 ( .A(n5877), .B(n5870), .Y(n5854) );
  AND2X1 U6284 ( .A(n5877), .B(n5871), .Y(n5855) );
  AND2X1 U6285 ( .A(n5852), .B(n5869), .Y(n5856) );
  AND2X1 U6286 ( .A(n5854), .B(n5869), .Y(n5857) );
  INVX1 U6287 ( .A(n6306), .Y(n6305) );
  AND2X1 U6288 ( .A(n5900), .B(n6161), .Y(n5858) );
  INVX1 U6289 ( .A(n10158), .Y(n10437) );
  AND2X1 U6290 ( .A(n6846), .B(n6155), .Y(n5859) );
  INVX1 U6291 ( .A(n7068), .Y(n7360) );
  AND2X1 U6292 ( .A(n7864), .B(n6155), .Y(n5862) );
  AND2X1 U6293 ( .A(n6913), .B(n6160), .Y(n5864) );
  AND2X1 U6294 ( .A(n5878), .B(n6516), .Y(n5866) );
  INVX1 U6295 ( .A(n6283), .Y(n6282) );
  INVX1 U6296 ( .A(n6304), .Y(n6303) );
  INVX1 U6297 ( .A(n6155), .Y(n6154) );
  INVX1 U6298 ( .A(n6302), .Y(n6301) );
  INVX1 U6299 ( .A(oprB[58]), .Y(n6164) );
  AND2X1 U6300 ( .A(op[5]), .B(n6362), .Y(n5867) );
  AND2X1 U6301 ( .A(op[2]), .B(n6360), .Y(n5868) );
  INVX1 U6302 ( .A(oprA[49]), .Y(n6291) );
  INVX1 U6303 ( .A(oprA[24]), .Y(n6326) );
  INVX1 U6304 ( .A(oprA[27]), .Y(n6318) );
  INVX1 U6305 ( .A(op[4]), .Y(n6516) );
  INVX1 U6306 ( .A(oprB[31]), .Y(n6151) );
  INVX1 U6307 ( .A(oprB[63]), .Y(n6158) );
  AND2X1 U6308 ( .A(ww[0]), .B(n6489), .Y(n5869) );
  AND2X1 U6309 ( .A(op[4]), .B(n5867), .Y(n5870) );
  AND2X1 U6310 ( .A(n5817), .B(op[4]), .Y(n5871) );
  INVX1 U6311 ( .A(oprA[51]), .Y(n6289) );
  INVX1 U6312 ( .A(oprA[35]), .Y(n6306) );
  INVX1 U6313 ( .A(oprA[36]), .Y(n6304) );
  INVX1 U6314 ( .A(op[5]), .Y(n6471) );
  INVX1 U6315 ( .A(oprA[19]), .Y(n6335) );
  INVX1 U6316 ( .A(ww[1]), .Y(n6489) );
  INVX1 U6317 ( .A(op[1]), .Y(n6362) );
  AND2X1 U6318 ( .A(ww[0]), .B(ww[1]), .Y(n5872) );
  AND2X1 U6319 ( .A(op[3]), .B(op[2]), .Y(n5873) );
  AND2X1 U6320 ( .A(ww[1]), .B(n6488), .Y(n5874) );
  INVX1 U6321 ( .A(shift_amount[2]), .Y(n6155) );
  INVX1 U6322 ( .A(shift_amount[3]), .Y(n6153) );
  INVX1 U6323 ( .A(n6470), .Y(n6497) );
  AND2X1 U6324 ( .A(n5866), .B(op[5]), .Y(n5875) );
  AND2X1 U6325 ( .A(n6499), .B(op[2]), .Y(n5876) );
  AND2X1 U6326 ( .A(op[3]), .B(n6472), .Y(n5877) );
  INVX1 U6327 ( .A(shift_amount[1]), .Y(n6157) );
  INVX1 U6328 ( .A(ww[0]), .Y(n6488) );
  INVX1 U6329 ( .A(oprA[57]), .Y(n6281) );
  INVX1 U6330 ( .A(n6021), .Y(n6339) );
  INVX1 U6331 ( .A(n6001), .Y(n6324) );
  INVX1 U6332 ( .A(n6350), .Y(n6050) );
  INVX1 U6333 ( .A(oprA[55]), .Y(n6284) );
  INVX1 U6334 ( .A(oprA[39]), .Y(n6299) );
  INVX1 U6335 ( .A(oprA[33]), .Y(n6310) );
  INVX1 U6336 ( .A(n6278), .Y(n6277) );
  INVX1 U6337 ( .A(n6274), .Y(n6273) );
  INVX1 U6338 ( .A(oprA[52]), .Y(n6287) );
  INVX1 U6339 ( .A(n37), .Y(n5884) );
  INVX1 U6340 ( .A(n6071), .Y(n6072) );
  INVX8 U6341 ( .A(n6164), .Y(n6163) );
  AOI22X1 U6342 ( .A(n6361), .B(n5991), .C(n6074), .D(n5911), .Y(n6366) );
  NAND3X1 U6343 ( .A(n5868), .B(n5867), .C(n6516), .Y(n6364) );
  AOI22X1 U6344 ( .A(n6363), .B(n5267), .C(n6075), .D(n9), .Y(n6365) );
  AOI22X1 U6345 ( .A(n6361), .B(n5992), .C(n6074), .D(n5915), .Y(n6368) );
  AOI22X1 U6346 ( .A(n6363), .B(n6217), .C(n6075), .D(n5897), .Y(n6367) );
  AOI22X1 U6347 ( .A(n6361), .B(n6314), .C(n6074), .D(n5918), .Y(n6370) );
  AOI22X1 U6348 ( .A(n6363), .B(n5908), .C(n6075), .D(n5899), .Y(n6369) );
  AOI22X1 U6349 ( .A(n6361), .B(n5276), .C(n6074), .D(n6275), .Y(n6372) );
  AOI22X1 U6350 ( .A(n6363), .B(n5882), .C(n6075), .D(n5902), .Y(n6371) );
  AOI22X1 U6351 ( .A(n6361), .B(n44), .C(n6074), .D(n67), .Y(n6374) );
  AOI22X1 U6352 ( .A(n6363), .B(n6222), .C(n6075), .D(n5906), .Y(n6373) );
  AOI22X1 U6353 ( .A(n6361), .B(n6319), .C(n6074), .D(n5925), .Y(n6376) );
  AOI22X1 U6354 ( .A(n6363), .B(n6224), .C(n6075), .D(n6163), .Y(n6375) );
  AOI22X1 U6355 ( .A(n6361), .B(n5283), .C(n6074), .D(n5927), .Y(n6378) );
  AOI22X1 U6356 ( .A(n6363), .B(n56), .C(n6075), .D(n6165), .Y(n6377) );
  AOI22X1 U6357 ( .A(n6361), .B(n5274), .C(n6074), .D(n6282), .Y(n6380) );
  AOI22X1 U6358 ( .A(n6363), .B(n6228), .C(n6075), .D(n6167), .Y(n6379) );
  AOI22X1 U6359 ( .A(n6361), .B(n6328), .C(n6074), .D(n5932), .Y(n6382) );
  AOI22X1 U6360 ( .A(n6363), .B(n46), .C(n6075), .D(n6169), .Y(n6381) );
  AOI22X1 U6361 ( .A(n6361), .B(n6330), .C(n6074), .D(n5933), .Y(n6384) );
  AOI22X1 U6362 ( .A(n6363), .B(n20), .C(n6431), .D(n6171), .Y(n6383) );
  AOI22X1 U6363 ( .A(n6361), .B(n6332), .C(n6074), .D(n5938), .Y(n6386) );
  AOI22X1 U6364 ( .A(n6363), .B(n6232), .C(n6075), .D(n6173), .Y(n6385) );
  AOI22X1 U6365 ( .A(n6361), .B(n6334), .C(n6074), .D(n5940), .Y(n6388) );
  AOI22X1 U6366 ( .A(n6363), .B(n6234), .C(n6431), .D(n6175), .Y(n6387) );
  AOI22X1 U6367 ( .A(n6361), .B(n5286), .C(n6074), .D(n6288), .Y(n6390) );
  AOI22X1 U6368 ( .A(n6363), .B(n5279), .C(n6075), .D(n6177), .Y(n6389) );
  AOI22X1 U6369 ( .A(n6361), .B(n6018), .C(n6074), .D(n5944), .Y(n6392) );
  AOI22X1 U6370 ( .A(n6363), .B(n6237), .C(n6075), .D(n6179), .Y(n6391) );
  AOI22X1 U6371 ( .A(n6361), .B(n6337), .C(n6074), .D(n5947), .Y(n6394) );
  AOI22X1 U6372 ( .A(n6363), .B(n6239), .C(n6431), .D(n6181), .Y(n6393) );
  AOI22X1 U6373 ( .A(n6361), .B(n5271), .C(n6074), .D(n5948), .Y(n6396) );
  AOI22X1 U6374 ( .A(n6363), .B(n6241), .C(n6075), .D(n6183), .Y(n6395) );
  AOI22X1 U6375 ( .A(n6361), .B(oprA[15]), .C(n6074), .D(n5952), .Y(n6398) );
  AOI22X1 U6376 ( .A(n6363), .B(n70), .C(n6075), .D(n6185), .Y(n6397) );
  AOI22X1 U6377 ( .A(n6361), .B(n6026), .C(n6074), .D(n5955), .Y(n6400) );
  AOI22X1 U6378 ( .A(n6363), .B(n6243), .C(n6075), .D(n6187), .Y(n6399) );
  AOI22X1 U6379 ( .A(n6361), .B(n6342), .C(n6074), .D(n5958), .Y(n6402) );
  AOI22X1 U6380 ( .A(n6363), .B(n6245), .C(n6431), .D(n6189), .Y(n6401) );
  AOI22X1 U6381 ( .A(n6361), .B(n6032), .C(n6074), .D(n5960), .Y(n6404) );
  AOI22X1 U6382 ( .A(n6363), .B(n6247), .C(n6075), .D(n6191), .Y(n6403) );
  AOI22X1 U6383 ( .A(n6361), .B(n37), .C(n6074), .D(n5964), .Y(n6406) );
  AOI22X1 U6384 ( .A(n6363), .B(n6249), .C(n6075), .D(n6193), .Y(n6405) );
  AOI22X1 U6385 ( .A(n6361), .B(n6034), .C(n6430), .D(n45), .Y(n6408) );
  AOI22X1 U6386 ( .A(n6363), .B(n6251), .C(n6431), .D(n6195), .Y(n6407) );
  AOI22X1 U6387 ( .A(n6361), .B(n6037), .C(n6430), .D(n5968), .Y(n6410) );
  AOI22X1 U6388 ( .A(n6363), .B(n6253), .C(n6075), .D(n6197), .Y(n6409) );
  AOI22X1 U6389 ( .A(n6361), .B(n6345), .C(n6430), .D(n6297), .Y(n6412) );
  AOI22X1 U6390 ( .A(n6363), .B(n6255), .C(n6431), .D(n6199), .Y(n6411) );
  AOI22X1 U6391 ( .A(n6361), .B(n6042), .C(n6430), .D(n5974), .Y(n6414) );
  AOI22X1 U6392 ( .A(n6363), .B(n6257), .C(n6075), .D(n6201), .Y(n6413) );
  AOI22X1 U6393 ( .A(n6361), .B(n6046), .C(n6430), .D(n5976), .Y(n6416) );
  AOI22X1 U6394 ( .A(n6363), .B(n6259), .C(n6431), .D(n6203), .Y(n6415) );
  AOI22X1 U6395 ( .A(n6361), .B(n6049), .C(n6430), .D(n5977), .Y(n6418) );
  AOI22X1 U6396 ( .A(n6363), .B(n6261), .C(n6075), .D(n6205), .Y(n6417) );
  AOI22X1 U6397 ( .A(n6361), .B(n6351), .C(n6074), .D(n6303), .Y(n6420) );
  AOI22X1 U6398 ( .A(n6363), .B(n6263), .C(n6075), .D(n6207), .Y(n6419) );
  AOI22X1 U6399 ( .A(n6361), .B(n6054), .C(n6430), .D(n5982), .Y(n6422) );
  AOI22X1 U6400 ( .A(n6363), .B(n3), .C(n6431), .D(n6209), .Y(n6421) );
  AOI22X1 U6401 ( .A(n6361), .B(n6354), .C(n6430), .D(n5984), .Y(n6424) );
  AOI22X1 U6402 ( .A(n6363), .B(n6267), .C(n6075), .D(n6211), .Y(n6423) );
  AOI22X1 U6403 ( .A(n6361), .B(n6356), .C(n6430), .D(n6308), .Y(n6426) );
  AOI22X1 U6404 ( .A(n6363), .B(n6269), .C(n6431), .D(n6213), .Y(n6425) );
  AOI22X1 U6405 ( .A(n6361), .B(n6061), .C(n6430), .D(n5988), .Y(n6428) );
  AOI22X1 U6406 ( .A(n6363), .B(n6271), .C(n6075), .D(n6215), .Y(n6427) );
  OAI21X1 U6407 ( .A(n5815), .B(n5814), .C(n5813), .Y(n6429) );
  OAI21X1 U6408 ( .A(n6457), .B(n5913), .C(n5301), .Y(mult32_A[30]) );
  OAI21X1 U6409 ( .A(n6457), .B(n6274), .C(n5347), .Y(mult32_A[29]) );
  OAI21X1 U6410 ( .A(n6457), .B(n6278), .C(n5307), .Y(mult32_A[26]) );
  OAI21X1 U6411 ( .A(n6457), .B(n6280), .C(n5297), .Y(mult32_A[25]) );
  OAI21X1 U6412 ( .A(n6457), .B(n6283), .C(n5467), .Y(mult32_A[24]) );
  OAI21X1 U6413 ( .A(n6457), .B(n6284), .C(n5599), .Y(mult32_A[23]) );
  OAI21X1 U6414 ( .A(n6457), .B(n6285), .C(n5529), .Y(mult32_A[22]) );
  OAI21X1 U6415 ( .A(n6457), .B(n5936), .C(n5293), .Y(mult32_A[21]) );
  OAI21X1 U6416 ( .A(n6457), .B(n6287), .C(n5369), .Y(mult32_A[20]) );
  OAI21X1 U6417 ( .A(n6457), .B(n6289), .C(n5323), .Y(mult32_A[19]) );
  OAI21X1 U6418 ( .A(n6457), .B(n5943), .C(n5313), .Y(mult32_A[18]) );
  OAI21X1 U6419 ( .A(n6457), .B(n6291), .C(n5409), .Y(mult32_A[17]) );
  OAI21X1 U6420 ( .A(n6457), .B(n6292), .C(n1917), .Y(mult32_A[16]) );
  OAI21X1 U6421 ( .A(n6457), .B(n6293), .C(n5333), .Y(mult32_A[14]) );
  OAI21X1 U6422 ( .A(n6457), .B(n6294), .C(n5287), .Y(mult32_A[13]) );
  AOI22X1 U6423 ( .A(n5964), .B(n5730), .C(n6076), .D(n37), .Y(n6458) );
  OAI21X1 U6424 ( .A(n6457), .B(n6295), .C(n5314), .Y(mult32_A[10]) );
  OAI21X1 U6425 ( .A(n6457), .B(n5967), .C(n5302), .Y(mult32_A[9]) );
  OAI21X1 U6426 ( .A(n6457), .B(n6298), .C(n5410), .Y(mult32_A[8]) );
  OAI21X1 U6427 ( .A(n6457), .B(n6299), .C(n5308), .Y(mult32_A[7]) );
  OAI21X1 U6428 ( .A(n6457), .B(n6300), .C(n5294), .Y(mult32_A[6]) );
  OAI21X1 U6429 ( .A(n6457), .B(n6302), .C(n5370), .Y(mult32_A[5]) );
  OAI21X1 U6430 ( .A(n6457), .B(n6304), .C(n5298), .Y(mult32_A[4]) );
  OAI21X1 U6431 ( .A(n6457), .B(n6306), .C(n5290), .Y(mult32_A[3]) );
  OAI21X1 U6432 ( .A(n6457), .B(n6307), .C(n5348), .Y(mult32_A[2]) );
  OAI21X1 U6433 ( .A(n6457), .B(n6309), .C(n5324), .Y(mult32_A[1]) );
  OAI21X1 U6434 ( .A(n6457), .B(n6311), .C(n5332), .Y(mult32_A[0]) );
  NAND3X1 U6435 ( .A(op[4]), .B(n6471), .C(n5878), .Y(n6470) );
  AOI22X1 U6436 ( .A(n3803), .B(n6108), .C(n3482), .D(n6106), .Y(n6477) );
  AOI22X1 U6437 ( .A(n1355), .B(n5772), .C(n841), .D(n6145), .Y(n6474) );
  NAND3X1 U6438 ( .A(n2378), .B(n5304), .C(n6475), .Y(n6542) );
  NAND3X1 U6439 ( .A(n4724), .B(n4769), .C(n4830), .Y(n6479) );
  NAND3X1 U6440 ( .A(n4870), .B(n6478), .C(n4966), .Y(n6783) );
  MUX2X1 U6441 ( .B(n2763), .A(n4962), .S(n5899), .Y(n6480) );
  AOI22X1 U6442 ( .A(n5820), .B(n6290), .C(n6551), .D(n5949), .Y(n6482) );
  AOI22X1 U6443 ( .A(n6579), .B(n5944), .C(n6517), .D(n5942), .Y(n6481) );
  AOI22X1 U6444 ( .A(n5820), .B(n5937), .C(n6551), .D(n5941), .Y(n6483) );
  AOI22X1 U6445 ( .A(n6733), .B(n5235), .C(n6974), .D(n5080), .Y(n6484) );
  OAI21X1 U6446 ( .A(n5902), .B(n6480), .C(n1740), .Y(n6487) );
  AOI22X1 U6447 ( .A(n5933), .B(n6077), .C(n5938), .D(n9626), .Y(n6485) );
  AOI22X1 U6448 ( .A(n6487), .B(n9647), .C(n9774), .D(n5140), .Y(n6495) );
  AOI22X1 U6449 ( .A(n3514), .B(n5830), .C(n3835), .D(n5828), .Y(n6494) );
  AOI22X1 U6450 ( .A(n3193), .B(n5827), .C(n1789), .D(n6121), .Y(n6492) );
  AOI22X1 U6451 ( .A(n1050), .B(n5786), .C(n1307), .D(n5785), .Y(n6491) );
  OAI21X1 U6452 ( .A(n6506), .B(n6155), .C(n5520), .Y(n10087) );
  AOI22X1 U6453 ( .A(n4949), .B(n10087), .C(n6498), .D(n5733), .Y(n6504) );
  NAND3X1 U6454 ( .A(op[3]), .B(n5867), .C(n6516), .Y(n6515) );
  OAI21X1 U6455 ( .A(n5900), .B(n10104), .C(n5650), .Y(n6502) );
  AOI22X1 U6456 ( .A(n5945), .B(n9632), .C(n6290), .D(n6081), .Y(n6501) );
  AOI22X1 U6457 ( .A(n5948), .B(n6080), .C(n5942), .D(n9688), .Y(n6500) );
  AOI22X1 U6458 ( .A(n5743), .B(n6502), .C(n5742), .D(n5214), .Y(n6503) );
  OAI21X1 U6459 ( .A(n6062), .B(n5587), .C(n1918), .Y(n9793) );
  OAI21X1 U6460 ( .A(n6082), .B(n5587), .C(n1919), .Y(n9795) );
  AOI22X1 U6461 ( .A(n5922), .B(n9793), .C(n5918), .D(n6065), .Y(n6512) );
  OAI21X1 U6462 ( .A(n6078), .B(n5587), .C(n1920), .Y(n9797) );
  OAI21X1 U6463 ( .A(n5911), .B(n6091), .C(n6089), .Y(n6510) );
  AOI22X1 U6464 ( .A(n5915), .B(n6066), .C(n8), .D(n6510), .Y(n6511) );
  NOR3X1 U6465 ( .A(n3689), .B(n4224), .C(n4586), .Y(n6534) );
  AOI22X1 U6466 ( .A(n2551), .B(n5831), .C(n2872), .D(n5829), .Y(n6526) );
  AOI22X1 U6467 ( .A(n472), .B(n6131), .C(n793), .D(n5825), .Y(n6525) );
  AOI22X1 U6468 ( .A(n5931), .B(n9969), .C(n1098), .D(n5826), .Y(n6523) );
  OAI21X1 U6469 ( .A(op[2]), .B(n5643), .C(n6089), .Y(n10315) );
  NAND3X1 U6470 ( .A(n4725), .B(n5724), .C(n6085), .Y(n7415) );
  NAND3X1 U6471 ( .A(n5720), .B(n5867), .C(n6516), .Y(n10517) );
  MUX2X1 U6472 ( .B(n6091), .A(n6068), .S(n8), .Y(n6519) );
  OAI21X1 U6473 ( .A(n4749), .B(n5008), .C(n6070), .Y(n6518) );
  NAND3X1 U6474 ( .A(n7369), .B(n5736), .C(n3650), .Y(n6521) );
  MUX2X1 U6475 ( .B(n6088), .A(n2786), .S(n5912), .Y(n6522) );
  AOI22X1 U6476 ( .A(n416), .B(n6117), .C(n552), .D(n5823), .Y(n6528) );
  AOI22X1 U6477 ( .A(n737), .B(n6119), .C(n2230), .D(n6104), .Y(n6527) );
  AOI22X1 U6478 ( .A(n1564), .B(n5779), .C(n873), .D(n6133), .Y(n6530) );
  AOI22X1 U6479 ( .A(n67), .B(n9500), .C(n5991), .D(n10502), .Y(n6529) );
  NOR3X1 U6480 ( .A(n3694), .B(n4225), .C(n4587), .Y(n6533) );
  AOI22X1 U6481 ( .A(n2972), .B(n6141), .C(n1837), .D(n5783), .Y(n6540) );
  AOI22X1 U6482 ( .A(n1612), .B(n6147), .C(n5951), .D(n6112), .Y(n6539) );
  AOI22X1 U6483 ( .A(n2840), .B(n6110), .C(n2519), .D(n6115), .Y(n6537) );
  NAND3X1 U6484 ( .A(n2379), .B(n2999), .C(n6538), .Y(n6541) );
  AOI22X1 U6485 ( .A(n3483), .B(n6106), .C(n3162), .D(n5776), .Y(n6545) );
  AOI22X1 U6486 ( .A(n842), .B(n5771), .C(n521), .D(n5773), .Y(n6543) );
  NAND3X1 U6487 ( .A(n5309), .B(n5542), .C(n5385), .Y(n6618) );
  AOI22X1 U6488 ( .A(n2520), .B(n6115), .C(n2199), .D(n6113), .Y(n6616) );
  MUX2X1 U6489 ( .B(n5915), .A(n5911), .S(n9), .Y(n6546) );
  AOI21X1 U6490 ( .A(n6517), .B(n5916), .C(n6720), .Y(n6547) );
  NAND3X1 U6491 ( .A(n4872), .B(n4770), .C(n3634), .Y(n6548) );
  AOI22X1 U6492 ( .A(n5863), .B(n4939), .C(n3357), .D(n5208), .Y(n6554) );
  AOI21X1 U6493 ( .A(n6517), .B(n6278), .C(n2363), .Y(n6578) );
  NAND3X1 U6494 ( .A(n4834), .B(n4768), .C(n3651), .Y(n6584) );
  AOI22X1 U6495 ( .A(n5820), .B(n5940), .C(n6551), .D(n5942), .Y(n6552) );
  AOI22X1 U6496 ( .A(n5758), .B(n6856), .C(n5753), .D(n5159), .Y(n6553) );
  AOI22X1 U6497 ( .A(n67), .B(n9793), .C(n5922), .D(n6065), .Y(n6561) );
  OAI21X1 U6498 ( .A(n5916), .B(n6091), .C(n6089), .Y(n6558) );
  OAI21X1 U6499 ( .A(n6063), .B(n5913), .C(n5598), .Y(n6846) );
  OAI21X1 U6500 ( .A(n6156), .B(n5508), .C(n5697), .Y(n9916) );
  AOI22X1 U6501 ( .A(n5897), .B(n6558), .C(n5859), .D(n9916), .Y(n6559) );
  NAND3X1 U6502 ( .A(n2381), .B(n3061), .C(n3379), .Y(n6562) );
  AOI21X1 U6503 ( .A(n6290), .B(n9632), .C(n5567), .Y(n6565) );
  OAI21X1 U6504 ( .A(n6082), .B(n6292), .C(n5566), .Y(n7363) );
  OAI21X1 U6505 ( .A(n6153), .B(n6292), .C(n5566), .Y(n7362) );
  OAI21X1 U6506 ( .A(n6567), .B(n5731), .C(n1921), .Y(n7353) );
  AOI21X1 U6507 ( .A(n6083), .B(n6278), .C(n2364), .Y(n6572) );
  OAI21X1 U6508 ( .A(n5926), .B(n6078), .C(n4835), .Y(n6569) );
  AOI22X1 U6509 ( .A(n6731), .B(n7353), .C(n6857), .D(n10375), .Y(n6574) );
  NAND3X1 U6510 ( .A(n4835), .B(n6062), .C(n3652), .Y(n6581) );
  AOI22X1 U6511 ( .A(n8968), .B(n4940), .C(n3515), .D(n6092), .Y(n6573) );
  AOI22X1 U6512 ( .A(n6579), .B(n6290), .C(n6517), .D(n5945), .Y(n6577) );
  AOI22X1 U6513 ( .A(n5820), .B(n10487), .C(n5896), .D(n7491), .Y(n6575) );
  OR2X2 U6514 ( .A(n1962), .B(n6292), .Y(n6576) );
  OAI21X1 U6515 ( .A(n5766), .B(n3352), .C(n6576), .Y(n7359) );
  OAI21X1 U6516 ( .A(n6279), .B(n5572), .C(n4834), .Y(n6580) );
  AOI22X1 U6517 ( .A(n6733), .B(n7359), .C(n6723), .D(n6855), .Y(n6587) );
  AOI21X1 U6518 ( .A(n6288), .B(n6079), .C(n7086), .Y(n6582) );
  AOI22X1 U6519 ( .A(n9774), .B(n5025), .C(n6704), .D(n4866), .Y(n6585) );
  NAND3X1 U6520 ( .A(n2382), .B(n3062), .C(n3380), .Y(n6588) );
  MUX2X1 U6521 ( .B(n6090), .A(n6067), .S(n5896), .Y(n6591) );
  NAND3X1 U6522 ( .A(n6591), .B(n6069), .C(n9803), .Y(n6592) );
  MUX2X1 U6523 ( .B(n6088), .A(n5538), .S(n5915), .Y(n6595) );
  AOI22X1 U6524 ( .A(n794), .B(n6137), .C(n5934), .D(n9969), .Y(n6593) );
  NAND3X1 U6525 ( .A(n6595), .B(n3064), .C(n3381), .Y(n6600) );
  AOI22X1 U6526 ( .A(n738), .B(n5790), .C(n2231), .D(n6104), .Y(n6598) );
  AOI22X1 U6527 ( .A(n2873), .B(n5829), .C(n473), .D(n6131), .Y(n6596) );
  NAND3X1 U6528 ( .A(n2383), .B(n3065), .C(n3382), .Y(n6599) );
  AOI22X1 U6529 ( .A(n5925), .B(n9500), .C(n5993), .D(n10502), .Y(n6602) );
  AOI22X1 U6530 ( .A(n417), .B(n5778), .C(n553), .D(n5823), .Y(n6601) );
  AOI22X1 U6531 ( .A(n3836), .B(n6096), .C(n3194), .D(n5827), .Y(n6605) );
  AOI22X1 U6532 ( .A(n1308), .B(n6125), .C(n874), .D(n5824), .Y(n6603) );
  NOR3X1 U6533 ( .A(n6607), .B(n4226), .C(n4295), .Y(n6608) );
  NAND3X1 U6534 ( .A(n2718), .B(n3063), .C(n6608), .Y(n6611) );
  OAI21X1 U6535 ( .A(n5722), .B(n6293), .C(n1922), .Y(n6613) );
  AOI21X1 U6536 ( .A(n2841), .B(n5780), .C(n6613), .Y(n6614) );
  NAND3X1 U6537 ( .A(n2380), .B(n5613), .C(n3635), .Y(n6617) );
  AOI22X1 U6538 ( .A(n3805), .B(n6108), .C(n3484), .D(n5774), .Y(n6623) );
  AOI22X1 U6539 ( .A(n1357), .B(n5772), .C(n843), .D(n5771), .Y(n6620) );
  NAND3X1 U6540 ( .A(n2384), .B(n5311), .C(n6621), .Y(n6696) );
  AOI22X1 U6541 ( .A(n5915), .B(n9632), .C(n5911), .D(n6081), .Y(n6624) );
  OAI21X1 U6542 ( .A(n6063), .B(n6274), .C(n1742), .Y(n7417) );
  OAI21X1 U6543 ( .A(oprB[61]), .B(n9846), .C(n5361), .Y(n6968) );
  AOI22X1 U6544 ( .A(n7417), .B(n6072), .C(n6968), .D(n5258), .Y(n6639) );
  NAND3X1 U6545 ( .A(n4727), .B(n4771), .C(n3653), .Y(n6632) );
  AOI22X1 U6546 ( .A(n5940), .B(n9632), .C(n6288), .D(n9626), .Y(n6634) );
  AOI22X1 U6547 ( .A(n5944), .B(n6079), .C(n5937), .D(n9688), .Y(n6633) );
  MUX2X1 U6548 ( .B(n6290), .A(n5949), .S(n5886), .Y(n6635) );
  MUX2X1 U6549 ( .B(n5515), .A(n5447), .S(n5889), .Y(n7150) );
  AOI22X1 U6550 ( .A(n8954), .B(n5515), .C(n6636), .D(n5770), .Y(n6637) );
  NAND3X1 U6551 ( .A(n2385), .B(n3066), .C(n3383), .Y(n6648) );
  AOI22X1 U6552 ( .A(n5820), .B(n6288), .C(n6551), .D(n5945), .Y(n6640) );
  NAND3X1 U6553 ( .A(n6974), .B(n7491), .C(n5188), .Y(n6642) );
  OAI21X1 U6554 ( .A(n9703), .B(n6278), .C(n1894), .Y(n6643) );
  AOI21X1 U6555 ( .A(n66), .B(n6065), .C(n6643), .Y(n6646) );
  OAI21X1 U6556 ( .A(n5918), .B(n6091), .C(n6089), .Y(n6644) );
  AOI22X1 U6557 ( .A(n17), .B(n6066), .C(n5900), .D(n6644), .Y(n6645) );
  MUX2X1 U6558 ( .B(n5948), .A(n6290), .S(n9688), .Y(n7427) );
  MUX2X1 U6559 ( .B(n5929), .A(n5926), .S(n9688), .Y(n6649) );
  AOI22X1 U6560 ( .A(n6730), .B(n7140), .C(n10375), .D(n6937), .Y(n6654) );
  MUX2X1 U6561 ( .B(n5927), .A(n5929), .S(n5887), .Y(n6650) );
  AOI21X1 U6562 ( .A(n5932), .B(n9626), .C(n5716), .Y(n6651) );
  OAI21X1 U6563 ( .A(n6062), .B(n6285), .C(n1895), .Y(n6939) );
  AOI22X1 U6564 ( .A(n3516), .B(n6092), .C(n3837), .D(n6096), .Y(n6652) );
  NAND3X1 U6565 ( .A(n2386), .B(n3067), .C(n3384), .Y(n6667) );
  MUX2X1 U6566 ( .B(n6280), .A(n6283), .S(n9), .Y(n6655) );
  MUX2X1 U6567 ( .B(n5929), .A(n5927), .S(n6517), .Y(n6921) );
  AOI22X1 U6568 ( .A(n5758), .B(n6662), .C(n6723), .D(n6656), .Y(n6665) );
  MUX2X1 U6569 ( .B(n6292), .A(n6291), .S(n6517), .Y(n6657) );
  MUX2X1 U6570 ( .B(n6291), .A(n6292), .S(n9), .Y(n6658) );
  MUX2X1 U6571 ( .B(n170), .A(n5641), .S(n5900), .Y(n6659) );
  OAI21X1 U6572 ( .A(n6160), .B(n5507), .C(n1923), .Y(n7171) );
  AOI22X1 U6573 ( .A(n5716), .B(n6721), .C(n6704), .D(n4974), .Y(n6663) );
  NAND3X1 U6574 ( .A(n2387), .B(n3068), .C(n3386), .Y(n6666) );
  MUX2X1 U6575 ( .B(n6090), .A(n6067), .S(n5900), .Y(n6668) );
  NAND3X1 U6576 ( .A(n6668), .B(n6069), .C(n9803), .Y(n6669) );
  MUX2X1 U6577 ( .B(n6088), .A(n5419), .S(n5918), .Y(n6672) );
  AOI22X1 U6578 ( .A(n795), .B(n6137), .C(n5938), .D(n9969), .Y(n6670) );
  NAND3X1 U6579 ( .A(n6672), .B(n3070), .C(n3387), .Y(n6677) );
  AOI22X1 U6580 ( .A(n739), .B(n5790), .C(n2232), .D(n6104), .Y(n6675) );
  AOI22X1 U6581 ( .A(n2874), .B(n5829), .C(n474), .D(n6131), .Y(n6673) );
  NAND3X1 U6582 ( .A(n2388), .B(n3071), .C(n3388), .Y(n6676) );
  AOI22X1 U6583 ( .A(n875), .B(n5824), .C(n5926), .D(n9500), .Y(n6680) );
  AOI22X1 U6584 ( .A(n418), .B(n5778), .C(n554), .D(n5823), .Y(n6678) );
  NAND3X1 U6585 ( .A(n5557), .B(n3072), .C(n5627), .Y(n6684) );
  AOI22X1 U6586 ( .A(n3195), .B(n6100), .C(n1791), .D(n6121), .Y(n6683) );
  AOI22X1 U6587 ( .A(n1309), .B(n6125), .C(n1566), .D(n6123), .Y(n6681) );
  NOR3X1 U6588 ( .A(n6685), .B(n4128), .C(n4299), .Y(n6686) );
  NAND3X1 U6589 ( .A(n2719), .B(n3069), .C(n6686), .Y(n6689) );
  AOI22X1 U6590 ( .A(n2942), .B(n6141), .C(n1839), .D(n6149), .Y(n6694) );
  AOI22X1 U6591 ( .A(n1614), .B(n6147), .C(n5958), .D(n6112), .Y(n6693) );
  AOI22X1 U6592 ( .A(n2842), .B(n6110), .C(n2521), .D(n6115), .Y(n6691) );
  NAND3X1 U6593 ( .A(n2389), .B(n3000), .C(n6692), .Y(n6695) );
  AOI22X1 U6594 ( .A(n3806), .B(n5775), .C(n3485), .D(n6106), .Y(n6701) );
  AOI22X1 U6595 ( .A(n1358), .B(n5772), .C(n844), .D(n5771), .Y(n6698) );
  NAND3X1 U6596 ( .A(n2390), .B(n5319), .C(n6699), .Y(n6764) );
  AOI21X1 U6597 ( .A(n5937), .B(n6079), .C(n6962), .Y(n6702) );
  AOI22X1 U6598 ( .A(n8968), .B(n4880), .C(n3517), .D(n6092), .Y(n6716) );
  AOI22X1 U6599 ( .A(n3838), .B(n6096), .C(n3196), .D(n5827), .Y(n6715) );
  AOI21X1 U6600 ( .A(n6551), .B(n5937), .C(n7093), .Y(n6703) );
  NAND3X1 U6601 ( .A(n5902), .B(n5948), .C(n7491), .Y(n7300) );
  OAI21X1 U6602 ( .A(n6705), .B(n5700), .C(n4696), .Y(n6713) );
  AOI22X1 U6603 ( .A(n6288), .B(n9632), .C(n5945), .D(n9626), .Y(n6706) );
  AOI22X1 U6604 ( .A(n5820), .B(n5944), .C(n6551), .D(n6290), .Y(n6709) );
  AOI22X1 U6605 ( .A(n5758), .B(n6708), .C(n5753), .D(n5107), .Y(n6711) );
  OAI21X1 U6606 ( .A(n158), .B(n5655), .C(n1758), .Y(n6712) );
  AOI22X1 U6607 ( .A(n5918), .B(n9632), .C(n5915), .D(n9626), .Y(n6718) );
  AOI22X1 U6608 ( .A(n5911), .B(n6080), .C(n5922), .D(n6083), .Y(n6717) );
  AOI22X1 U6609 ( .A(n5820), .B(n5915), .C(n6551), .D(n5912), .Y(n6719) );
  AOI22X1 U6610 ( .A(n5183), .B(n6072), .C(n6968), .D(n5260), .Y(n6729) );
  OAI21X1 U6611 ( .A(n6063), .B(n4795), .C(n5719), .Y(n6722) );
  NAND3X1 U6612 ( .A(n4728), .B(n4772), .C(n3654), .Y(n6726) );
  AOI22X1 U6613 ( .A(n5929), .B(n2775), .C(n3358), .D(n5208), .Y(n6728) );
  OAI21X1 U6614 ( .A(n4752), .B(n4796), .C(n4695), .Y(n6732) );
  OAI21X1 U6615 ( .A(n4750), .B(n5029), .C(n9791), .Y(n6734) );
  AOI22X1 U6616 ( .A(n5949), .B(n6734), .C(n5927), .D(n9793), .Y(n6738) );
  OAI21X1 U6617 ( .A(n5922), .B(n6091), .C(n6089), .Y(n6735) );
  AOI22X1 U6618 ( .A(n67), .B(n6066), .C(n5903), .D(n6735), .Y(n6736) );
  NOR3X1 U6619 ( .A(n3699), .B(n4227), .C(n4306), .Y(n6756) );
  AOI22X1 U6620 ( .A(n2233), .B(n5838), .C(n2554), .D(n6102), .Y(n6747) );
  AOI22X1 U6621 ( .A(n2875), .B(n5829), .C(n475), .D(n6131), .Y(n6746) );
  AOI22X1 U6622 ( .A(n796), .B(n5825), .C(n5940), .D(n9969), .Y(n6744) );
  MUX2X1 U6623 ( .B(n6091), .A(n6068), .S(n5903), .Y(n6740) );
  NOR3X1 U6624 ( .A(n5728), .B(n9731), .C(n6740), .Y(n6741) );
  MUX2X1 U6625 ( .B(n10522), .A(n6741), .S(n5922), .Y(n6742) );
  AOI21X1 U6626 ( .A(n1101), .B(n5826), .C(n6742), .Y(n6743) );
  AOI22X1 U6627 ( .A(n5276), .B(n10502), .C(n419), .D(n5778), .Y(n6749) );
  AOI22X1 U6628 ( .A(n555), .B(n5823), .C(n740), .D(n6119), .Y(n6748) );
  AOI22X1 U6629 ( .A(n1792), .B(n5777), .C(n1053), .D(n6129), .Y(n6752) );
  AOI22X1 U6630 ( .A(n1567), .B(n5779), .C(n876), .D(n5824), .Y(n6750) );
  NAND3X1 U6631 ( .A(n2391), .B(n5339), .C(n5360), .Y(n6753) );
  NOR3X1 U6632 ( .A(n3703), .B(n4228), .C(n4310), .Y(n6755) );
  AOI22X1 U6633 ( .A(n2973), .B(n6141), .C(n1840), .D(n6149), .Y(n6762) );
  AOI22X1 U6634 ( .A(n1615), .B(n6147), .C(n5960), .D(n6112), .Y(n6761) );
  AOI22X1 U6635 ( .A(n2843), .B(n5780), .C(n2522), .D(n6115), .Y(n6759) );
  NAND3X1 U6636 ( .A(n2392), .B(n3001), .C(n6760), .Y(n6763) );
  AOI22X1 U6637 ( .A(n3807), .B(n6108), .C(n3486), .D(n5774), .Y(n6769) );
  AOI22X1 U6638 ( .A(n1359), .B(n6139), .C(n845), .D(n5771), .Y(n6766) );
  NAND3X1 U6639 ( .A(n5534), .B(n5679), .C(n6767), .Y(n6820) );
  AOI22X1 U6640 ( .A(n5753), .B(n5235), .C(n9774), .D(n5214), .Y(n6774) );
  AOI22X1 U6641 ( .A(n6704), .B(n5080), .C(n8968), .D(n5140), .Y(n6773) );
  AOI22X1 U6642 ( .A(n3518), .B(n6092), .C(n3839), .D(n6096), .Y(n6771) );
  AOI22X1 U6643 ( .A(n3197), .B(n6100), .C(n1793), .D(n6121), .Y(n6770) );
  AOI22X1 U6644 ( .A(n5922), .B(n9632), .C(n5918), .D(n9626), .Y(n6775) );
  AOI21X1 U6645 ( .A(n6551), .B(n5916), .C(n6778), .Y(n6779) );
  AOI22X1 U6646 ( .A(n5095), .B(n6072), .C(n6968), .D(n5162), .Y(n6785) );
  OAI21X1 U6647 ( .A(n9846), .B(n6160), .C(n5502), .Y(n6964) );
  AOI22X1 U6648 ( .A(n5743), .B(n6964), .C(n5208), .D(n4962), .Y(n6784) );
  OAI21X1 U6649 ( .A(n10375), .B(n6723), .C(n6282), .Y(n6786) );
  OAI21X1 U6650 ( .A(n6063), .B(n5012), .C(n5519), .Y(n6789) );
  OAI21X1 U6651 ( .A(n6063), .B(n5721), .C(n10383), .Y(n9853) );
  OAI21X1 U6652 ( .A(n67), .B(n6091), .C(n6089), .Y(n6792) );
  AOI22X1 U6653 ( .A(n5905), .B(n6792), .C(n4949), .D(n6073), .Y(n6793) );
  NOR3X1 U6654 ( .A(n3708), .B(n4229), .C(n4311), .Y(n6812) );
  AOI22X1 U6655 ( .A(n1054), .B(n5786), .C(n1311), .D(n5785), .Y(n6800) );
  AOI22X1 U6656 ( .A(n1568), .B(n5779), .C(n877), .D(n5824), .Y(n6799) );
  AOI22X1 U6657 ( .A(n27), .B(n10502), .C(n420), .D(n5778), .Y(n6797) );
  AOI22X1 U6658 ( .A(n556), .B(n5823), .C(n741), .D(n5790), .Y(n6796) );
  NAND3X1 U6659 ( .A(n2393), .B(n5496), .C(n6798), .Y(n6810) );
  MUX2X1 U6660 ( .B(n6090), .A(n6067), .S(n5905), .Y(n6801) );
  MUX2X1 U6661 ( .B(n5832), .A(n5336), .S(n67), .Y(n6805) );
  AOI22X1 U6662 ( .A(n797), .B(n6137), .C(n6288), .D(n9969), .Y(n6803) );
  NAND3X1 U6663 ( .A(n6805), .B(n5384), .C(n3389), .Y(n6809) );
  AOI22X1 U6664 ( .A(n2234), .B(n5838), .C(n2555), .D(n6102), .Y(n6807) );
  AOI22X1 U6665 ( .A(n2876), .B(n5829), .C(n476), .D(n6131), .Y(n6806) );
  NOR3X1 U6666 ( .A(n3713), .B(n4129), .C(n4588), .Y(n6811) );
  AOI22X1 U6667 ( .A(n2974), .B(n6141), .C(n1841), .D(n6149), .Y(n6818) );
  AOI22X1 U6668 ( .A(n1616), .B(n5784), .C(n5964), .D(n6112), .Y(n6817) );
  AOI22X1 U6669 ( .A(n2844), .B(n6110), .C(n2523), .D(n6115), .Y(n6815) );
  NAND3X1 U6670 ( .A(n2394), .B(n5358), .C(n6816), .Y(n6819) );
  AOI22X1 U6671 ( .A(n3808), .B(n5775), .C(n3487), .D(n6106), .Y(n6825) );
  AOI22X1 U6672 ( .A(n1360), .B(n5772), .C(n846), .D(n5771), .Y(n6822) );
  NAND3X1 U6673 ( .A(n5316), .B(n5327), .C(n6823), .Y(n6883) );
  AOI22X1 U6674 ( .A(n5916), .B(n9500), .C(n6319), .D(n10502), .Y(n6827) );
  AOI22X1 U6675 ( .A(n421), .B(n5778), .C(n557), .D(n5823), .Y(n6826) );
  AOI22X1 U6676 ( .A(n1794), .B(n5777), .C(n1055), .D(n6129), .Y(n6830) );
  AOI22X1 U6677 ( .A(n1569), .B(n5779), .C(n878), .D(n5824), .Y(n6828) );
  NAND3X1 U6678 ( .A(n2395), .B(n5426), .C(n5390), .Y(n6831) );
  MUX2X1 U6679 ( .B(n6090), .A(n6067), .S(n6163), .Y(n6833) );
  MUX2X1 U6680 ( .B(n6088), .A(n5604), .S(n5924), .Y(n6837) );
  AOI22X1 U6681 ( .A(n798), .B(n6137), .C(n5944), .D(n9969), .Y(n6835) );
  NAND3X1 U6682 ( .A(n6837), .B(n5494), .C(n3390), .Y(n6842) );
  AOI22X1 U6683 ( .A(n742), .B(n5790), .C(n2235), .D(n5838), .Y(n6840) );
  AOI22X1 U6684 ( .A(n2877), .B(n5829), .C(n477), .D(n6131), .Y(n6838) );
  NAND3X1 U6685 ( .A(n2396), .B(n3073), .C(n3391), .Y(n6841) );
  OAI21X1 U6686 ( .A(n5924), .B(n6091), .C(n6089), .Y(n6843) );
  AOI21X1 U6687 ( .A(n6163), .B(n6843), .C(n5036), .Y(n6863) );
  AOI22X1 U6688 ( .A(n67), .B(n9632), .C(n5922), .D(n9626), .Y(n6845) );
  AOI22X1 U6689 ( .A(n5918), .B(n6079), .C(n5924), .D(n9688), .Y(n6844) );
  MUX2X1 U6690 ( .B(n7089), .A(n6847), .S(n5889), .Y(n7340) );
  AOI21X1 U6691 ( .A(n6517), .B(n5924), .C(n5807), .Y(n6848) );
  MUX2X1 U6692 ( .B(n4849), .A(n5640), .S(n5899), .Y(n6852) );
  AOI22X1 U6693 ( .A(n7340), .B(n9916), .C(n7346), .D(n4939), .Y(n6862) );
  AOI22X1 U6694 ( .A(n6856), .B(n6854), .C(n6855), .D(n6920), .Y(n6860) );
  AOI22X1 U6695 ( .A(n6858), .B(n5822), .C(n6857), .D(n7147), .Y(n6859) );
  AOI22X1 U6696 ( .A(n8968), .B(n5025), .C(n3519), .D(n6092), .Y(n6865) );
  AOI22X1 U6697 ( .A(n3840), .B(n5828), .C(n3198), .D(n5827), .Y(n6864) );
  AOI22X1 U6698 ( .A(n6974), .B(n7359), .C(n6704), .D(n5159), .Y(n6871) );
  AOI22X1 U6699 ( .A(n5833), .B(n7353), .C(n6791), .D(n4940), .Y(n6869) );
  NOR3X1 U6700 ( .A(n3714), .B(n4230), .C(n4314), .Y(n6873) );
  NAND3X1 U6701 ( .A(n2720), .B(n3074), .C(n6873), .Y(n6876) );
  AOI22X1 U6702 ( .A(n2943), .B(n6141), .C(n1842), .D(n6149), .Y(n6881) );
  AOI22X1 U6703 ( .A(n1617), .B(n5784), .C(n45), .D(n6112), .Y(n6880) );
  AOI22X1 U6704 ( .A(n2845), .B(n6110), .C(n2524), .D(n6115), .Y(n6878) );
  NAND3X1 U6705 ( .A(n2397), .B(n5386), .C(n6879), .Y(n6882) );
  AOI22X1 U6706 ( .A(n2557), .B(n6102), .C(n2878), .D(n5829), .Y(n6888) );
  OAI21X1 U6707 ( .A(n5583), .B(n5967), .C(n1924), .Y(n6885) );
  AOI21X1 U6708 ( .A(n1361), .B(n5848), .C(n6885), .Y(n6886) );
  AOI22X1 U6709 ( .A(n558), .B(n5823), .C(n743), .D(n5790), .Y(n6890) );
  AOI22X1 U6710 ( .A(n879), .B(n5824), .C(n5918), .D(n9500), .Y(n6892) );
  AOI22X1 U6711 ( .A(n6322), .B(n10502), .C(n422), .D(n5778), .Y(n6891) );
  NOR3X1 U6712 ( .A(n3719), .B(n4231), .C(n4589), .Y(n6949) );
  AOI22X1 U6713 ( .A(n2846), .B(n5835), .C(n478), .D(n5839), .Y(n6901) );
  AOI22X1 U6714 ( .A(n6290), .B(n6094), .C(n1104), .D(n5826), .Y(n6898) );
  MUX2X1 U6715 ( .B(n6090), .A(n6067), .S(n6165), .Y(n6895) );
  MUX2X1 U6716 ( .B(n5832), .A(n5422), .S(n5926), .Y(n6897) );
  NAND3X1 U6717 ( .A(n5317), .B(n5482), .C(n6899), .Y(n6908) );
  AOI22X1 U6718 ( .A(n3809), .B(n5845), .C(n2204), .D(n5843), .Y(n6903) );
  AOI22X1 U6719 ( .A(n1618), .B(n5846), .C(n1843), .D(n5842), .Y(n6905) );
  AOI22X1 U6720 ( .A(n3167), .B(n5844), .C(n3488), .D(n5847), .Y(n6904) );
  NOR3X1 U6721 ( .A(n3723), .B(n4232), .C(n4590), .Y(n6948) );
  AOI22X1 U6722 ( .A(n17), .B(n6080), .C(n5927), .D(n6083), .Y(n6909) );
  AOI22X1 U6723 ( .A(n7417), .B(n10574), .C(n6964), .D(n5258), .Y(n6912) );
  OAI21X1 U6724 ( .A(n6071), .B(n164), .C(n1774), .Y(n6917) );
  AOI21X1 U6725 ( .A(n6090), .B(n6280), .C(n10564), .Y(n6915) );
  NAND3X1 U6726 ( .A(n5903), .B(n10487), .C(n5864), .Y(n6914) );
  OAI21X1 U6727 ( .A(n2759), .B(n6166), .C(n1896), .Y(n6916) );
  NOR3X1 U6728 ( .A(n6917), .B(n6916), .C(n5036), .Y(n6931) );
  AOI22X1 U6729 ( .A(n7407), .B(n5770), .C(n6662), .D(n6854), .Y(n6919) );
  OAI21X1 U6730 ( .A(n6921), .B(n5650), .C(n1790), .Y(n6929) );
  AOI21X1 U6731 ( .A(n6517), .B(n6279), .C(n6922), .Y(n6923) );
  AOI22X1 U6732 ( .A(n6968), .B(n5059), .C(n6926), .D(n6974), .Y(n6927) );
  OAI21X1 U6733 ( .A(n7427), .B(n5578), .C(n1806), .Y(n6928) );
  AOI22X1 U6734 ( .A(n3841), .B(n6096), .C(n3199), .D(n5827), .Y(n6936) );
  AOI22X1 U6735 ( .A(n1056), .B(n5786), .C(n1313), .D(n5785), .Y(n6933) );
  NAND3X1 U6736 ( .A(n5413), .B(n5606), .C(n6934), .Y(n6945) );
  AOI22X1 U6737 ( .A(n5716), .B(n5822), .C(n7147), .D(n6937), .Y(n6944) );
  AOI22X1 U6738 ( .A(n6704), .B(n5188), .C(n6866), .D(n4974), .Y(n6943) );
  OAI21X1 U6739 ( .A(n7148), .B(n5520), .C(n1925), .Y(n6941) );
  AOI21X1 U6740 ( .A(n3520), .B(n6092), .C(n6941), .Y(n6942) );
  NOR3X1 U6741 ( .A(n4121), .B(n4130), .C(n4321), .Y(n6947) );
  NAND3X1 U6742 ( .A(n6949), .B(n6948), .C(n6947), .Y(n6950) );
  AOI22X1 U6743 ( .A(n3810), .B(n6108), .C(n3489), .D(n5774), .Y(n6955) );
  AOI22X1 U6744 ( .A(n1362), .B(n5772), .C(n848), .D(n5771), .Y(n6952) );
  NAND3X1 U6745 ( .A(n5417), .B(n5614), .C(n6953), .Y(n7003) );
  AOI22X1 U6746 ( .A(n6704), .B(n5107), .C(n6866), .D(n4808), .Y(n6960) );
  AOI22X1 U6747 ( .A(n6791), .B(n4880), .C(n8968), .D(n5013), .Y(n6959) );
  AOI22X1 U6748 ( .A(n3521), .B(n6092), .C(n3842), .D(n6096), .Y(n6957) );
  AOI22X1 U6749 ( .A(n3200), .B(n5827), .C(n1796), .D(n6121), .Y(n6956) );
  AOI22X1 U6750 ( .A(n5927), .B(n9632), .C(n5925), .D(n9626), .Y(n6961) );
  AOI22X1 U6751 ( .A(n6964), .B(n5260), .C(n5068), .D(n6072), .Y(n6970) );
  AOI21X1 U6752 ( .A(n6579), .B(n6279), .C(n6708), .Y(n6965) );
  AOI22X1 U6753 ( .A(n6968), .B(n5110), .C(n6708), .D(n6854), .Y(n6969) );
  NAND3X1 U6754 ( .A(n5729), .B(n6095), .C(n3655), .Y(n6973) );
  OAI21X1 U6755 ( .A(n4751), .B(n5029), .C(n10033), .Y(n6975) );
  OAI21X1 U6756 ( .A(n6282), .B(n6091), .C(n6089), .Y(n6976) );
  AOI22X1 U6757 ( .A(n6167), .B(n6976), .C(n5183), .D(n10574), .Y(n6977) );
  NOR3X1 U6758 ( .A(n3724), .B(n4233), .C(n4326), .Y(n6995) );
  AOI22X1 U6759 ( .A(n1057), .B(n5786), .C(n1314), .D(n5785), .Y(n6984) );
  AOI22X1 U6760 ( .A(n1571), .B(n5779), .C(n880), .D(n5824), .Y(n6983) );
  AOI22X1 U6761 ( .A(n5922), .B(n9500), .C(n5274), .D(n10502), .Y(n6981) );
  AOI22X1 U6762 ( .A(n423), .B(n6117), .C(n559), .D(n5823), .Y(n6980) );
  AOI21X1 U6763 ( .A(n5822), .B(n9688), .C(n6570), .Y(n6985) );
  NAND3X1 U6764 ( .A(n2698), .B(n5588), .C(n6085), .Y(n10557) );
  MUX2X1 U6765 ( .B(n6090), .A(n6067), .S(n6167), .Y(n6986) );
  MUX2X1 U6766 ( .B(n6088), .A(n2937), .S(n6282), .Y(n6990) );
  AOI22X1 U6767 ( .A(n479), .B(n5839), .C(n800), .D(n5825), .Y(n6988) );
  AOI22X1 U6768 ( .A(n744), .B(n5790), .C(n2237), .D(n6104), .Y(n6992) );
  AOI22X1 U6769 ( .A(n2558), .B(n6102), .C(n2879), .D(n6086), .Y(n6991) );
  NOR3X1 U6770 ( .A(n3729), .B(n4131), .C(n4591), .Y(n6994) );
  AOI22X1 U6771 ( .A(n2975), .B(n6141), .C(n1844), .D(n6149), .Y(n7001) );
  AOI22X1 U6772 ( .A(n1619), .B(n5784), .C(n5970), .D(n6112), .Y(n7000) );
  AOI22X1 U6773 ( .A(n2847), .B(n5780), .C(n2526), .D(n5781), .Y(n6998) );
  NAND3X1 U6774 ( .A(n2398), .B(n5556), .C(n6999), .Y(n7002) );
  AOI22X1 U6775 ( .A(n3811), .B(n5775), .C(n3490), .D(n6106), .Y(n7008) );
  AOI22X1 U6776 ( .A(n1363), .B(n5772), .C(n849), .D(n5771), .Y(n7005) );
  NAND3X1 U6777 ( .A(n2399), .B(n5340), .C(n7006), .Y(n7060) );
  OAI21X1 U6778 ( .A(n6063), .B(n5446), .C(n6095), .Y(n10072) );
  AOI21X1 U6779 ( .A(n5925), .B(n5800), .C(n7009), .Y(n7010) );
  AOI22X1 U6780 ( .A(n5912), .B(n10072), .C(n6625), .D(n4976), .Y(n7021) );
  AOI21X1 U6781 ( .A(n6579), .B(n5929), .C(n7013), .Y(n7014) );
  AOI22X1 U6782 ( .A(n10500), .B(n5095), .C(n6627), .D(n4909), .Y(n7020) );
  AOI22X1 U6783 ( .A(n3522), .B(n6092), .C(n3843), .D(n6096), .Y(n7018) );
  AOI22X1 U6784 ( .A(n3201), .B(n6100), .C(n1797), .D(n6121), .Y(n7017) );
  AOI22X1 U6785 ( .A(n5743), .B(n5795), .C(n6704), .D(n5235), .Y(n7024) );
  AOI22X1 U6786 ( .A(n6866), .B(n5080), .C(n7022), .D(n5162), .Y(n7023) );
  OAI21X1 U6787 ( .A(n5932), .B(n6091), .C(n6089), .Y(n7025) );
  OAI21X1 U6788 ( .A(n5729), .B(n6292), .C(n5582), .Y(n7151) );
  AOI21X1 U6789 ( .A(n6169), .B(n7025), .C(n7151), .Y(n7034) );
  OAI21X1 U6790 ( .A(n6287), .B(n5725), .C(n5595), .Y(n7027) );
  AOI21X1 U6791 ( .A(n7070), .B(n5934), .C(n7027), .Y(n7030) );
  AOI22X1 U6792 ( .A(n5792), .B(n6290), .C(n7167), .D(n5949), .Y(n7029) );
  AOI22X1 U6793 ( .A(n7070), .B(n5945), .C(n7284), .D(n6288), .Y(n7028) );
  MUX2X1 U6794 ( .B(n2764), .A(n7308), .S(n6173), .Y(n7031) );
  AOI22X1 U6795 ( .A(n5140), .B(n6073), .C(n7031), .D(n5733), .Y(n7032) );
  NOR3X1 U6796 ( .A(n3734), .B(n4234), .C(n4329), .Y(n7052) );
  AOI22X1 U6797 ( .A(n1058), .B(n5786), .C(n1315), .D(n5785), .Y(n7040) );
  AOI22X1 U6798 ( .A(n1572), .B(n6123), .C(n881), .D(n5824), .Y(n7039) );
  AOI22X1 U6799 ( .A(n6288), .B(n9500), .C(n6004), .D(n10502), .Y(n7037) );
  AOI22X1 U6800 ( .A(n408), .B(n5778), .C(n560), .D(n5823), .Y(n7036) );
  NAND3X1 U6801 ( .A(n7284), .B(n5589), .C(n6174), .Y(n7041) );
  MUX2X1 U6802 ( .B(n6091), .A(n6068), .S(n6169), .Y(n7042) );
  AOI21X1 U6803 ( .A(n7138), .B(n7284), .C(n7042), .Y(n7043) );
  NAND3X1 U6804 ( .A(n7492), .B(n6085), .C(n3636), .Y(n7044) );
  MUX2X1 U6805 ( .B(n6088), .A(n2787), .S(n5932), .Y(n7047) );
  AOI22X1 U6806 ( .A(n480), .B(n6131), .C(n801), .D(n5825), .Y(n7045) );
  AOI22X1 U6807 ( .A(n729), .B(n5790), .C(n2238), .D(n5838), .Y(n7049) );
  AOI22X1 U6808 ( .A(n2559), .B(n6102), .C(n2880), .D(n6086), .Y(n7048) );
  NOR3X1 U6809 ( .A(n3739), .B(n4135), .C(n4592), .Y(n7051) );
  AOI22X1 U6810 ( .A(n2976), .B(n6141), .C(n1845), .D(n6149), .Y(n7058) );
  AOI22X1 U6811 ( .A(n1620), .B(n6147), .C(n5974), .D(n6112), .Y(n7057) );
  AOI22X1 U6812 ( .A(n2848), .B(n6110), .C(n2527), .D(n6115), .Y(n7055) );
  NAND3X1 U6813 ( .A(n2400), .B(n3002), .C(n7056), .Y(n7059) );
  AOI22X1 U6814 ( .A(n3812), .B(n5775), .C(n3491), .D(n5774), .Y(n7065) );
  AOI22X1 U6815 ( .A(n1364), .B(n5772), .C(n850), .D(n5771), .Y(n7062) );
  NAND3X1 U6816 ( .A(n2401), .B(n5355), .C(n7063), .Y(n7130) );
  AOI22X1 U6817 ( .A(n5859), .B(n5791), .C(n5858), .D(n7359), .Y(n7079) );
  AOI21X1 U6818 ( .A(n7284), .B(n5943), .C(n2365), .Y(n7069) );
  NAND3X1 U6819 ( .A(n4836), .B(n5725), .C(n3656), .Y(n7068) );
  OAI21X1 U6820 ( .A(n6290), .B(n4798), .C(n4836), .Y(n7071) );
  AOI21X1 U6821 ( .A(n5792), .B(n6286), .C(n7230), .Y(n7072) );
  OAI21X1 U6822 ( .A(n6289), .B(n5725), .C(n1897), .Y(n7080) );
  AOI22X1 U6823 ( .A(n5480), .B(n7070), .C(n5760), .D(n5589), .Y(n7074) );
  OAI21X1 U6824 ( .A(n7075), .B(n5656), .C(n1838), .Y(n7076) );
  AOI22X1 U6825 ( .A(n5745), .B(n7361), .C(n7076), .D(n6174), .Y(n7077) );
  OAI21X1 U6826 ( .A(n5760), .B(n7080), .C(n7138), .Y(n7081) );
  OAI21X1 U6827 ( .A(n5801), .B(n162), .C(n7081), .Y(n7085) );
  AOI21X1 U6828 ( .A(n6090), .B(n6285), .C(n10564), .Y(n7083) );
  AOI21X1 U6829 ( .A(n5863), .B(n5808), .C(n7151), .Y(n7082) );
  OAI21X1 U6830 ( .A(n2760), .B(n6172), .C(n1898), .Y(n7084) );
  NOR3X1 U6831 ( .A(n3744), .B(n7085), .C(n7084), .Y(n7122) );
  AOI21X1 U6832 ( .A(n5929), .B(n9626), .C(n5718), .Y(n7088) );
  OAI21X1 U6833 ( .A(n6062), .B(n6280), .C(n1899), .Y(n7354) );
  AOI22X1 U6834 ( .A(n6625), .B(n7354), .C(n10375), .D(n7362), .Y(n7096) );
  AOI21X1 U6835 ( .A(n5820), .B(n5929), .C(n7090), .Y(n7091) );
  AOI22X1 U6836 ( .A(n6627), .B(n4912), .C(n3523), .D(n6092), .Y(n7094) );
  NAND3X1 U6837 ( .A(n2402), .B(n3075), .C(n3392), .Y(n7101) );
  AOI22X1 U6838 ( .A(n6721), .B(n7363), .C(n6866), .D(n5159), .Y(n7099) );
  AOI22X1 U6839 ( .A(n5834), .B(n7353), .C(n6626), .D(n5718), .Y(n7097) );
  NAND3X1 U6840 ( .A(n2403), .B(n3076), .C(n3393), .Y(n7100) );
  AOI22X1 U6841 ( .A(n481), .B(n5839), .C(n802), .D(n5825), .Y(n7107) );
  MUX2X1 U6842 ( .B(n6091), .A(n6068), .S(n6171), .Y(n7102) );
  MUX2X1 U6843 ( .B(n10522), .A(n5475), .S(n5933), .Y(n7104) );
  AOI21X1 U6844 ( .A(n1107), .B(n6127), .C(n7104), .Y(n7105) );
  NAND3X1 U6845 ( .A(n2404), .B(n3078), .C(n3637), .Y(n7112) );
  AOI22X1 U6846 ( .A(n561), .B(n5823), .C(n730), .D(n6119), .Y(n7110) );
  AOI22X1 U6847 ( .A(n2560), .B(n6102), .C(n2881), .D(n6086), .Y(n7108) );
  NAND3X1 U6848 ( .A(n2405), .B(n3079), .C(n3394), .Y(n7111) );
  AOI22X1 U6849 ( .A(n1573), .B(n5779), .C(n882), .D(n5824), .Y(n7115) );
  AOI22X1 U6850 ( .A(n6007), .B(n10502), .C(n409), .D(n5778), .Y(n7113) );
  AOI22X1 U6851 ( .A(n3844), .B(n5828), .C(n3202), .D(n5827), .Y(n7118) );
  AOI22X1 U6852 ( .A(n1059), .B(n5786), .C(n1316), .D(n6125), .Y(n7116) );
  NOR3X1 U6853 ( .A(n7119), .B(n4139), .C(n4336), .Y(n7120) );
  NAND3X1 U6854 ( .A(n7122), .B(n3077), .C(n7120), .Y(n7123) );
  AOI22X1 U6855 ( .A(n2944), .B(n6141), .C(n1846), .D(n6149), .Y(n7128) );
  AOI22X1 U6856 ( .A(n1621), .B(n5784), .C(n5975), .D(n6112), .Y(n7127) );
  AOI22X1 U6857 ( .A(n2849), .B(n6110), .C(n2528), .D(n6115), .Y(n7125) );
  NAND3X1 U6858 ( .A(n2406), .B(n3003), .C(n7126), .Y(n7129) );
  AOI22X1 U6859 ( .A(n3813), .B(n6108), .C(n3492), .D(n6106), .Y(n7135) );
  AOI22X1 U6860 ( .A(n1365), .B(n5772), .C(n851), .D(n5771), .Y(n7132) );
  NAND3X1 U6861 ( .A(n5334), .B(n5380), .C(n7133), .Y(n7205) );
  AOI22X1 U6862 ( .A(n5792), .B(n6288), .C(n7167), .D(n5944), .Y(n7137) );
  AOI22X1 U6863 ( .A(n7070), .B(n6286), .C(n7284), .D(n5938), .Y(n7136) );
  AOI22X1 U6864 ( .A(n7140), .B(n4762), .C(n3371), .D(n5158), .Y(n7145) );
  MUX2X1 U6865 ( .B(n6290), .A(n5948), .S(n6169), .Y(n7141) );
  MUX2X1 U6866 ( .B(n5949), .A(n6290), .S(n7284), .Y(n7142) );
  AOI22X1 U6867 ( .A(n5745), .B(n7430), .C(n5795), .D(n5258), .Y(n7143) );
  OAI21X1 U6868 ( .A(n6156), .B(n5731), .C(n5449), .Y(n10491) );
  OAI21X1 U6869 ( .A(n5715), .B(n5400), .C(n4697), .Y(n10505) );
  OAI21X1 U6870 ( .A(n7408), .B(n7150), .C(n1926), .Y(n7155) );
  NAND3X1 U6871 ( .A(n5841), .B(n7491), .C(n5188), .Y(n7154) );
  OAI21X1 U6872 ( .A(n5937), .B(n6091), .C(n6089), .Y(n7152) );
  NOR3X1 U6873 ( .A(n3748), .B(n7155), .C(n4340), .Y(n7197) );
  AOI22X1 U6874 ( .A(n5888), .B(n6285), .C(shift_amount[3]), .D(n6284), .Y(
        n7156) );
  AOI22X1 U6875 ( .A(n6625), .B(n4875), .C(n10500), .D(n5043), .Y(n7166) );
  AOI22X1 U6876 ( .A(n3524), .B(n6092), .C(n3845), .D(n6096), .Y(n7164) );
  NAND3X1 U6877 ( .A(n2407), .B(n3080), .C(n3395), .Y(n7177) );
  NAND3X1 U6878 ( .A(n2721), .B(n3081), .C(n5725), .Y(n7170) );
  AOI21X1 U6879 ( .A(n7284), .B(n5936), .C(n2342), .Y(n7422) );
  AOI22X1 U6880 ( .A(n4898), .B(n7285), .C(n7171), .D(n6161), .Y(n7175) );
  AOI22X1 U6881 ( .A(n7022), .B(n5059), .C(n7404), .D(n6626), .Y(n7173) );
  NAND3X1 U6882 ( .A(n2408), .B(n3082), .C(n3396), .Y(n7176) );
  MUX2X1 U6883 ( .B(n6090), .A(n6067), .S(n6173), .Y(n7178) );
  MUX2X1 U6884 ( .B(n6088), .A(n5353), .S(n5938), .Y(n7182) );
  AOI22X1 U6885 ( .A(n803), .B(n6137), .C(n5918), .D(n9969), .Y(n7180) );
  NAND3X1 U6886 ( .A(n7182), .B(n3084), .C(n3397), .Y(n7187) );
  AOI22X1 U6887 ( .A(n731), .B(n5790), .C(n2240), .D(n6104), .Y(n7185) );
  AOI22X1 U6888 ( .A(n2882), .B(n5829), .C(n482), .D(n5839), .Y(n7183) );
  NAND3X1 U6889 ( .A(n2409), .B(n3085), .C(n3398), .Y(n7186) );
  AOI22X1 U6890 ( .A(n883), .B(n5824), .C(n6290), .D(n9500), .Y(n7190) );
  AOI22X1 U6891 ( .A(n410), .B(n6117), .C(n562), .D(n5823), .Y(n7188) );
  AOI22X1 U6892 ( .A(n3203), .B(n5827), .C(n1799), .D(n6121), .Y(n7193) );
  AOI22X1 U6893 ( .A(n1317), .B(n6125), .C(n1574), .D(n6123), .Y(n7191) );
  NOR3X1 U6894 ( .A(n7194), .B(n4143), .C(n4343), .Y(n7195) );
  NAND3X1 U6895 ( .A(n7197), .B(n3083), .C(n7195), .Y(n7198) );
  AOI22X1 U6896 ( .A(n2945), .B(n6141), .C(n1847), .D(n6149), .Y(n7203) );
  AOI22X1 U6897 ( .A(n1622), .B(n5784), .C(n5978), .D(n6112), .Y(n7202) );
  AOI22X1 U6898 ( .A(n2850), .B(n5780), .C(n2529), .D(n5781), .Y(n7200) );
  NAND3X1 U6899 ( .A(n2410), .B(n3004), .C(n7201), .Y(n7204) );
  AOI22X1 U6900 ( .A(n3814), .B(n5775), .C(n3493), .D(n5774), .Y(n7210) );
  AOI22X1 U6901 ( .A(n1366), .B(n6139), .C(n852), .D(n5771), .Y(n7207) );
  NAND3X1 U6902 ( .A(n5374), .B(n5427), .C(n7208), .Y(n7271) );
  AOI22X1 U6903 ( .A(n7172), .B(n5183), .C(n7022), .D(n5110), .Y(n7220) );
  AOI22X1 U6904 ( .A(n10500), .B(n5068), .C(n6627), .D(n4979), .Y(n7219) );
  AOI22X1 U6905 ( .A(n3525), .B(n5830), .C(n3846), .D(n6096), .Y(n7217) );
  AOI22X1 U6906 ( .A(n3204), .B(n5827), .C(n1800), .D(n6121), .Y(n7216) );
  AOI21X1 U6907 ( .A(n5858), .B(n7221), .C(n5763), .Y(n7227) );
  AOI22X1 U6908 ( .A(n6971), .B(n5834), .C(n7490), .D(n5715), .Y(n7223) );
  NOR3X1 U6909 ( .A(n4948), .B(n9500), .C(n5745), .Y(n7225) );
  NAND3X1 U6910 ( .A(n2699), .B(n3086), .C(n7225), .Y(n7228) );
  AOI22X1 U6911 ( .A(n5949), .B(n2774), .C(n5795), .D(n5260), .Y(n7232) );
  AOI22X1 U6912 ( .A(n5792), .B(n5934), .C(n7167), .D(n5931), .Y(n7229) );
  AOI22X1 U6913 ( .A(n7285), .B(n4883), .C(n6866), .D(n5107), .Y(n7231) );
  OAI21X1 U6914 ( .A(n6286), .B(n6091), .C(n6089), .Y(n7234) );
  AOI21X1 U6915 ( .A(n6175), .B(n7234), .C(n7233), .Y(n7246) );
  NAND3X1 U6916 ( .A(n4726), .B(n7238), .C(n4967), .Y(n7476) );
  AOI22X1 U6917 ( .A(n5792), .B(n5945), .C(n7167), .D(n6290), .Y(n7240) );
  NAND3X1 U6918 ( .A(n2722), .B(n4773), .C(n3399), .Y(n7243) );
  AOI22X1 U6919 ( .A(n4899), .B(n5628), .C(n3359), .D(n5158), .Y(n7244) );
  NOR3X1 U6920 ( .A(n3752), .B(n4235), .C(n4377), .Y(n7263) );
  AOI22X1 U6921 ( .A(n1061), .B(n5786), .C(n1318), .D(n6125), .Y(n7252) );
  AOI22X1 U6922 ( .A(n1575), .B(n5779), .C(n884), .D(n5824), .Y(n7251) );
  AOI22X1 U6923 ( .A(n5285), .B(n10502), .C(n411), .D(n5778), .Y(n7249) );
  AOI22X1 U6924 ( .A(n563), .B(n5823), .C(n732), .D(n5790), .Y(n7248) );
  NAND3X1 U6925 ( .A(n5471), .B(n5559), .C(n7250), .Y(n7261) );
  MUX2X1 U6926 ( .B(n6090), .A(n6067), .S(n6175), .Y(n7253) );
  MUX2X1 U6927 ( .B(n6088), .A(n5288), .S(n5940), .Y(n7257) );
  AOI22X1 U6928 ( .A(n804), .B(n6137), .C(n17), .D(n9969), .Y(n7255) );
  AOI22X1 U6929 ( .A(n2241), .B(n5838), .C(n2562), .D(n6102), .Y(n7259) );
  AOI22X1 U6930 ( .A(n2883), .B(n5829), .C(n483), .D(n5839), .Y(n7258) );
  NOR3X1 U6931 ( .A(n3757), .B(n4147), .C(n4593), .Y(n7262) );
  AOI22X1 U6932 ( .A(n2977), .B(n6141), .C(n1848), .D(n6149), .Y(n7269) );
  AOI22X1 U6933 ( .A(n1623), .B(n5784), .C(n6303), .D(n6112), .Y(n7268) );
  AOI22X1 U6934 ( .A(n2851), .B(n6110), .C(n2530), .D(n6115), .Y(n7266) );
  NAND3X1 U6935 ( .A(n2411), .B(n3005), .C(n7267), .Y(n7270) );
  AOI22X1 U6936 ( .A(n3815), .B(n6108), .C(n3494), .D(n6106), .Y(n7276) );
  AOI22X1 U6937 ( .A(n1367), .B(n6139), .C(n853), .D(n5771), .Y(n7273) );
  NAND3X1 U6938 ( .A(n5473), .B(n5548), .C(n7274), .Y(n7333) );
  AOI22X1 U6939 ( .A(n885), .B(n5824), .C(n6016), .D(n10502), .Y(n7278) );
  AOI22X1 U6940 ( .A(n412), .B(n6117), .C(n564), .D(n5823), .Y(n7277) );
  AOI22X1 U6941 ( .A(n3205), .B(n6100), .C(n1801), .D(n6121), .Y(n7281) );
  AOI22X1 U6942 ( .A(n1319), .B(n6125), .C(n1576), .D(n6123), .Y(n7279) );
  NAND3X1 U6943 ( .A(n5416), .B(n5610), .C(n5552), .Y(n7282) );
  OAI21X1 U6944 ( .A(n5568), .B(n5638), .C(n5732), .Y(n7413) );
  MUX2X1 U6945 ( .B(n6090), .A(n6067), .S(n6177), .Y(n7286) );
  NAND3X1 U6946 ( .A(n7371), .B(n7286), .C(n7369), .Y(n7287) );
  MUX2X1 U6947 ( .B(n6088), .A(n2788), .S(n5942), .Y(n7290) );
  AOI22X1 U6948 ( .A(n805), .B(n6137), .C(n66), .D(n9969), .Y(n7288) );
  NAND3X1 U6949 ( .A(n7290), .B(n5560), .C(n5491), .Y(n7295) );
  AOI22X1 U6950 ( .A(n733), .B(n5790), .C(n2242), .D(n6104), .Y(n7293) );
  AOI22X1 U6951 ( .A(n2884), .B(n5829), .C(n484), .D(n5839), .Y(n7291) );
  NAND3X1 U6952 ( .A(n2412), .B(n3087), .C(n3400), .Y(n7294) );
  AOI21X1 U6953 ( .A(n7070), .B(n7285), .C(n5749), .Y(n7296) );
  OAI21X1 U6954 ( .A(n5763), .B(n5654), .C(n5949), .Y(n7301) );
  OAI21X1 U6955 ( .A(n10375), .B(n5745), .C(n5948), .Y(n7299) );
  NAND3X1 U6956 ( .A(n7301), .B(n5582), .C(n7299), .Y(n7345) );
  AOI21X1 U6957 ( .A(n6286), .B(n5226), .C(n4717), .Y(n7315) );
  AOI21X1 U6958 ( .A(n5792), .B(n7285), .C(n5751), .Y(n7302) );
  AOI21X1 U6959 ( .A(n7167), .B(n7285), .C(n5750), .Y(n7304) );
  AOI22X1 U6960 ( .A(n5937), .B(n5239), .C(n5933), .D(n5242), .Y(n7314) );
  OAI21X1 U6961 ( .A(n6288), .B(n6091), .C(n6089), .Y(n7306) );
  AOI22X1 U6962 ( .A(n5932), .B(n2776), .C(n6177), .D(n7306), .Y(n7312) );
  AOI22X1 U6963 ( .A(n5214), .B(n6073), .C(n5158), .D(n4826), .Y(n7311) );
  AOI22X1 U6964 ( .A(n7022), .B(n4909), .C(n10500), .D(n4976), .Y(n7317) );
  AOI22X1 U6965 ( .A(n3526), .B(n6092), .C(n3847), .D(n6096), .Y(n7316) );
  AOI22X1 U6966 ( .A(n5743), .B(n5803), .C(n5795), .D(n5162), .Y(n7321) );
  AOI22X1 U6967 ( .A(n6866), .B(n5235), .C(n7172), .D(n5095), .Y(n7319) );
  NOR3X1 U6968 ( .A(n3758), .B(n4236), .C(n4381), .Y(n7323) );
  NAND3X1 U6969 ( .A(n2723), .B(n3088), .C(n7323), .Y(n7326) );
  AOI22X1 U6970 ( .A(n2946), .B(n6141), .C(n1849), .D(n6149), .Y(n7331) );
  AOI22X1 U6971 ( .A(n1624), .B(n5784), .C(n6305), .D(n6112), .Y(n7330) );
  AOI22X1 U6972 ( .A(n2852), .B(n5780), .C(n2531), .D(n5781), .Y(n7328) );
  NAND3X1 U6973 ( .A(n2413), .B(n3006), .C(n7329), .Y(n7332) );
  AOI22X1 U6974 ( .A(n3816), .B(n5775), .C(n3495), .D(n5774), .Y(n7338) );
  AOI22X1 U6975 ( .A(n1368), .B(n6139), .C(n854), .D(n5771), .Y(n7335) );
  NAND3X1 U6976 ( .A(n5349), .B(n5485), .C(n7336), .Y(n7398) );
  AOI22X1 U6977 ( .A(n5941), .B(n5239), .C(n5937), .D(n5242), .Y(n7344) );
  OAI21X1 U6978 ( .A(n9500), .B(n7339), .C(n5934), .Y(n7343) );
  OAI21X1 U6979 ( .A(n5944), .B(n6091), .C(n6089), .Y(n7341) );
  AOI22X1 U6980 ( .A(n6179), .B(n7341), .C(n5791), .D(n7340), .Y(n7342) );
  NAND3X1 U6981 ( .A(n2414), .B(n7343), .C(n3401), .Y(n7350) );
  NAND3X1 U6982 ( .A(n7070), .B(n5932), .C(n5747), .Y(n7348) );
  AOI22X1 U6983 ( .A(n5808), .B(n7346), .C(n5942), .D(n5226), .Y(n7347) );
  NAND3X1 U6984 ( .A(n7418), .B(n3052), .C(n3402), .Y(n7349) );
  AOI22X1 U6985 ( .A(n7351), .B(n5718), .C(n7022), .D(n4912), .Y(n7357) );
  AOI22X1 U6986 ( .A(n10500), .B(n7354), .C(n3527), .D(n6092), .Y(n7355) );
  NAND3X1 U6987 ( .A(n2415), .B(n3089), .C(n3403), .Y(n7368) );
  AOI22X1 U6988 ( .A(n7360), .B(n7358), .C(n5841), .D(n7359), .Y(n7366) );
  AOI22X1 U6989 ( .A(n5822), .B(n7363), .C(n7147), .D(n7362), .Y(n7364) );
  NAND3X1 U6990 ( .A(n2416), .B(n3090), .C(n3404), .Y(n7367) );
  MUX2X1 U6991 ( .B(n6090), .A(n6067), .S(n6179), .Y(n7370) );
  NAND3X1 U6992 ( .A(n7371), .B(n7370), .C(n7369), .Y(n7372) );
  MUX2X1 U6993 ( .B(n6088), .A(n2789), .S(n5945), .Y(n7375) );
  AOI22X1 U6994 ( .A(n806), .B(n6137), .C(n5925), .D(n9969), .Y(n7373) );
  NAND3X1 U6995 ( .A(n7375), .B(n3092), .C(n3405), .Y(n7380) );
  AOI22X1 U6996 ( .A(n734), .B(n5790), .C(n2243), .D(n6104), .Y(n7378) );
  AOI22X1 U6997 ( .A(n2885), .B(n5829), .C(n485), .D(n5839), .Y(n7376) );
  NAND3X1 U6998 ( .A(n2417), .B(n3093), .C(n3406), .Y(n7379) );
  OR2X2 U6999 ( .A(n1991), .B(n2114), .Y(n7387) );
  AOI22X1 U7000 ( .A(n1577), .B(n5779), .C(n886), .D(n5824), .Y(n7383) );
  AOI22X1 U7001 ( .A(n413), .B(n5778), .C(n565), .D(n5823), .Y(n7381) );
  AOI22X1 U7002 ( .A(n3848), .B(n5828), .C(n3206), .D(n5827), .Y(n7386) );
  AOI22X1 U7003 ( .A(n1063), .B(n5786), .C(n1320), .D(n5785), .Y(n7384) );
  NOR3X1 U7004 ( .A(n7387), .B(n4151), .C(n4385), .Y(n7388) );
  NAND3X1 U7005 ( .A(n2724), .B(n3091), .C(n7388), .Y(n7391) );
  AOI22X1 U7006 ( .A(n2948), .B(n6141), .C(n1850), .D(n6149), .Y(n7396) );
  AOI22X1 U7007 ( .A(n1625), .B(n5784), .C(oprA[34]), .D(n6112), .Y(n7395) );
  AOI22X1 U7008 ( .A(n2853), .B(n5780), .C(n2532), .D(n6115), .Y(n7393) );
  NAND3X1 U7009 ( .A(n2419), .B(n3007), .C(n7394), .Y(n7397) );
  OR2X2 U7010 ( .A(n1988), .B(n107), .Y(result[50]) );
  AOI22X1 U7011 ( .A(n3817), .B(n5775), .C(n3496), .D(n5774), .Y(n7403) );
  AOI22X1 U7012 ( .A(n1369), .B(n5772), .C(n855), .D(n5771), .Y(n7400) );
  NAND3X1 U7013 ( .A(n5412), .B(n5615), .C(n7401), .Y(n7464) );
  AOI22X1 U7014 ( .A(n3528), .B(n5830), .C(n2244), .D(n5838), .Y(n7444) );
  AOI22X1 U7015 ( .A(n7358), .B(n5704), .C(n7404), .D(n7351), .Y(n7406) );
  OAI21X1 U7016 ( .A(n7408), .B(n4797), .C(n1869), .Y(n7409) );
  AOI21X1 U7017 ( .A(n5795), .B(n5059), .C(n7409), .Y(n7412) );
  AOI22X1 U7018 ( .A(n5803), .B(n5258), .C(n7022), .D(n4860), .Y(n7411) );
  AOI22X1 U7019 ( .A(n5940), .B(n5242), .C(n6288), .D(n5239), .Y(n7410) );
  MUX2X1 U7020 ( .B(n6091), .A(n6068), .S(n6181), .Y(n7414) );
  NOR3X1 U7021 ( .A(n4846), .B(n7414), .C(n7413), .Y(n7416) );
  MUX2X1 U7022 ( .B(n10522), .A(n7416), .S(n5947), .Y(n7437) );
  AOI22X1 U7023 ( .A(n8485), .B(n7417), .C(n7172), .D(n5043), .Y(n7419) );
  AOI21X1 U7024 ( .A(n10500), .B(n4875), .C(n2366), .Y(n7436) );
  AOI22X1 U7025 ( .A(n4898), .B(n5747), .C(n6926), .D(n5841), .Y(n7435) );
  OAI21X1 U7026 ( .A(n6290), .B(n6091), .C(n6089), .Y(n7425) );
  AOI22X1 U7027 ( .A(n5926), .B(n6094), .C(n5938), .D(n9500), .Y(n7423) );
  OAI21X1 U7028 ( .A(n6099), .B(n6338), .C(n1870), .Y(n7424) );
  AOI21X1 U7029 ( .A(n6181), .B(n7425), .C(n7424), .Y(n7426) );
  OAI21X1 U7030 ( .A(n7428), .B(n7427), .C(n1900), .Y(n7429) );
  AOI21X1 U7031 ( .A(n7138), .B(n7430), .C(n7429), .Y(n7432) );
  NAND3X1 U7032 ( .A(n5864), .B(n10487), .C(n6161), .Y(n7431) );
  AOI21X1 U7033 ( .A(n5944), .B(n5226), .C(n2367), .Y(n7434) );
  NOR3X1 U7034 ( .A(n3763), .B(n7437), .C(n4389), .Y(n7440) );
  AOI22X1 U7035 ( .A(n3849), .B(n5828), .C(n3207), .D(n6100), .Y(n7438) );
  NAND3X1 U7036 ( .A(n7440), .B(n3094), .C(n3407), .Y(n7441) );
  AOI21X1 U7037 ( .A(n2886), .B(n6086), .C(n2343), .Y(n7443) );
  NAND3X1 U7038 ( .A(n2420), .B(n3053), .C(n3657), .Y(n7445) );
  AOI21X1 U7039 ( .A(n887), .B(n5824), .C(n2344), .Y(n7448) );
  NAND3X1 U7040 ( .A(n2700), .B(n3095), .C(n3658), .Y(n7449) );
  AOI21X1 U7041 ( .A(n1112), .B(n5826), .C(n2345), .Y(n7452) );
  NAND3X1 U7042 ( .A(n2701), .B(n3096), .C(n5689), .Y(n7453) );
  AOI21X1 U7043 ( .A(n486), .B(n5839), .C(n120), .Y(n7456) );
  AOI22X1 U7044 ( .A(n1064), .B(n5786), .C(n807), .D(n5825), .Y(n7454) );
  NAND3X1 U7045 ( .A(n2702), .B(n3097), .C(n3408), .Y(n7457) );
  AOI22X1 U7046 ( .A(n2949), .B(n6141), .C(n1851), .D(n6149), .Y(n7462) );
  AOI22X1 U7047 ( .A(n1626), .B(n5784), .C(n6308), .D(n6112), .Y(n7461) );
  AOI22X1 U7048 ( .A(n2854), .B(n5780), .C(n2533), .D(n5781), .Y(n7459) );
  NAND3X1 U7049 ( .A(n2421), .B(n3008), .C(n7460), .Y(n7463) );
  AOI22X1 U7050 ( .A(n3818), .B(n5775), .C(n3497), .D(n5774), .Y(n7469) );
  AOI22X1 U7051 ( .A(n1370), .B(n6139), .C(n856), .D(n5771), .Y(n7466) );
  NAND3X1 U7052 ( .A(n5535), .B(n5680), .C(n7467), .Y(n7516) );
  AOI22X1 U7053 ( .A(n1322), .B(n6125), .C(n487), .D(n5839), .Y(n7508) );
  AOI22X1 U7054 ( .A(n5747), .B(n4883), .C(n5795), .D(n5110), .Y(n7474) );
  AOI22X1 U7055 ( .A(n7172), .B(n5068), .C(n7022), .D(n4979), .Y(n7473) );
  AOI22X1 U7056 ( .A(n3529), .B(n5830), .C(n3850), .D(n6096), .Y(n7471) );
  AOI22X1 U7057 ( .A(n4899), .B(n10574), .C(n5803), .D(n5260), .Y(n7477) );
  OAI21X1 U7058 ( .A(n7475), .B(n5644), .C(n1871), .Y(n7482) );
  AOI22X1 U7059 ( .A(n6290), .B(n5226), .C(n5944), .D(n5239), .Y(n7480) );
  OAI21X1 U7060 ( .A(n5949), .B(n6091), .C(n6089), .Y(n7478) );
  AOI22X1 U7061 ( .A(n6288), .B(n5242), .C(n6183), .D(n7478), .Y(n7479) );
  NOR3X1 U7062 ( .A(n3768), .B(n7482), .C(n4594), .Y(n7505) );
  AOI22X1 U7063 ( .A(n1804), .B(n6121), .C(n1579), .D(n6123), .Y(n7487) );
  AOI22X1 U7064 ( .A(n888), .B(n5824), .C(n5941), .D(n9500), .Y(n7486) );
  OAI21X1 U7065 ( .A(n6340), .B(n6099), .C(n5331), .Y(n7484) );
  AOI21X1 U7066 ( .A(n567), .B(n5823), .C(n7484), .Y(n7485) );
  AOI22X1 U7067 ( .A(n5929), .B(n6094), .C(n1113), .D(n6127), .Y(n7498) );
  AOI21X1 U7068 ( .A(n7221), .B(n5841), .C(n7488), .Y(n7495) );
  MUX2X1 U7069 ( .B(n6090), .A(n6067), .S(n6183), .Y(n7494) );
  AOI21X1 U7070 ( .A(n6971), .B(n7222), .C(n9576), .Y(n7489) );
  NAND3X1 U7071 ( .A(n5364), .B(n5400), .C(n3638), .Y(n10555) );
  NOR3X1 U7072 ( .A(n5265), .B(n5263), .C(n4855), .Y(n7493) );
  NAND3X1 U7073 ( .A(n2703), .B(n7494), .C(n7493), .Y(n7496) );
  MUX2X1 U7074 ( .B(n6088), .A(n2790), .S(n5948), .Y(n7497) );
  AOI22X1 U7075 ( .A(n736), .B(n5790), .C(n2245), .D(n5838), .Y(n7500) );
  AOI22X1 U7076 ( .A(n2566), .B(n6102), .C(n2887), .D(n6086), .Y(n7499) );
  NOR3X1 U7077 ( .A(n73), .B(n4237), .C(n4595), .Y(n7504) );
  NAND3X1 U7078 ( .A(n2422), .B(n5686), .C(n3639), .Y(n7509) );
  AOI22X1 U7079 ( .A(n2951), .B(n6141), .C(n1852), .D(n5783), .Y(n7514) );
  AOI22X1 U7080 ( .A(n1627), .B(n5784), .C(n5989), .D(n10480), .Y(n7513) );
  AOI22X1 U7081 ( .A(n2855), .B(n5780), .C(n2534), .D(n6115), .Y(n7511) );
  NAND3X1 U7082 ( .A(n124), .B(n5436), .C(n7512), .Y(n7515) );
  AOI22X1 U7083 ( .A(n3819), .B(n5775), .C(n3498), .D(n6106), .Y(n7521) );
  AOI22X1 U7084 ( .A(n1371), .B(n6139), .C(n857), .D(n5771), .Y(n7518) );
  NAND3X1 U7085 ( .A(n2423), .B(n5354), .C(n7519), .Y(n7575) );
  NAND3X1 U7086 ( .A(n4729), .B(n4775), .C(n4831), .Y(n7523) );
  NAND3X1 U7087 ( .A(n4730), .B(n7522), .C(n4968), .Y(n7805) );
  MUX2X1 U7088 ( .B(n2765), .A(n4963), .S(n6189), .Y(n7524) );
  AOI22X1 U7089 ( .A(n5767), .B(n6308), .C(n7586), .D(n5989), .Y(n7526) );
  AOI22X1 U7090 ( .A(n7611), .B(n5983), .C(n7550), .D(n5981), .Y(n7525) );
  AOI22X1 U7091 ( .A(n5767), .B(n6301), .C(n7586), .D(n5980), .Y(n7527) );
  AOI22X1 U7092 ( .A(n7755), .B(n5254), .C(n7988), .D(n5113), .Y(n7528) );
  OAI21X1 U7093 ( .A(n6191), .B(n7524), .C(n1872), .Y(n7531) );
  AOI22X1 U7094 ( .A(n5975), .B(n9632), .C(n6301), .D(n9626), .Y(n7529) );
  AOI22X1 U7095 ( .A(n7531), .B(n9647), .C(n9774), .D(n5143), .Y(n7536) );
  AOI22X1 U7096 ( .A(n3530), .B(n6092), .C(n3851), .D(n6096), .Y(n7535) );
  AOI22X1 U7097 ( .A(n3209), .B(n6100), .C(n1773), .D(n6121), .Y(n7533) );
  AOI22X1 U7098 ( .A(n1034), .B(n5786), .C(n1291), .D(n5785), .Y(n7532) );
  AOI22X1 U7099 ( .A(n4952), .B(n10087), .C(n7538), .D(n5733), .Y(n7543) );
  OAI21X1 U7100 ( .A(n6189), .B(n10104), .C(n5006), .Y(n7541) );
  AOI22X1 U7101 ( .A(n5984), .B(n9632), .C(n6308), .D(n9626), .Y(n7540) );
  AOI22X1 U7102 ( .A(n6080), .B(n5988), .C(n6305), .D(n6083), .Y(n7539) );
  AOI22X1 U7103 ( .A(n5744), .B(n7541), .C(n5742), .D(n5215), .Y(n7542) );
  AOI22X1 U7104 ( .A(n5961), .B(n9793), .C(n5957), .D(n6065), .Y(n7546) );
  OAI21X1 U7105 ( .A(n5952), .B(n6091), .C(n6089), .Y(n7544) );
  AOI22X1 U7106 ( .A(n5953), .B(n6066), .C(n6185), .D(n7544), .Y(n7545) );
  NOR3X1 U7107 ( .A(n3902), .B(n4238), .C(n4596), .Y(n7567) );
  AOI22X1 U7108 ( .A(n2567), .B(n6102), .C(n2888), .D(n5829), .Y(n7559) );
  AOI22X1 U7109 ( .A(n456), .B(n5839), .C(n777), .D(n5825), .Y(n7558) );
  AOI22X1 U7110 ( .A(n5974), .B(n6094), .C(n1114), .D(n6127), .Y(n7556) );
  NAND3X1 U7111 ( .A(n4731), .B(n5724), .C(n6085), .Y(n7549) );
  MUX2X1 U7112 ( .B(n6091), .A(n6068), .S(n6185), .Y(n7552) );
  OAI21X1 U7113 ( .A(n4753), .B(n5009), .C(n6070), .Y(n7551) );
  NAND3X1 U7114 ( .A(n8433), .B(n5736), .C(n3659), .Y(n7554) );
  MUX2X1 U7115 ( .B(n6088), .A(n2791), .S(n5952), .Y(n7555) );
  AOI22X1 U7116 ( .A(n400), .B(n5778), .C(n568), .D(n5823), .Y(n7561) );
  AOI22X1 U7117 ( .A(n721), .B(n5790), .C(n2246), .D(n5838), .Y(n7560) );
  AOI22X1 U7118 ( .A(n1548), .B(n5779), .C(n889), .D(n5824), .Y(n7563) );
  AOI22X1 U7119 ( .A(n5965), .B(n9500), .C(n6098), .D(n59), .Y(n7562) );
  NOR3X1 U7120 ( .A(n3907), .B(n4239), .C(n4597), .Y(n7566) );
  AOI22X1 U7121 ( .A(n2978), .B(n6141), .C(n1853), .D(n5783), .Y(n7573) );
  AOI22X1 U7122 ( .A(n1628), .B(n5784), .C(n5911), .D(n10480), .Y(n7572) );
  AOI22X1 U7123 ( .A(n2856), .B(n5780), .C(n2535), .D(n6115), .Y(n7570) );
  NAND3X1 U7124 ( .A(n2425), .B(n5387), .C(n7571), .Y(n7574) );
  AOI22X1 U7125 ( .A(n3820), .B(n6108), .C(n3499), .D(n5774), .Y(n7580) );
  AOI22X1 U7126 ( .A(n1372), .B(n6139), .C(n858), .D(n6145), .Y(n7577) );
  NAND3X1 U7127 ( .A(n2426), .B(n5378), .C(n7578), .Y(n7649) );
  MUX2X1 U7128 ( .B(n5953), .A(n5952), .S(n6185), .Y(n7581) );
  AOI21X1 U7129 ( .A(n7550), .B(n5953), .C(n7747), .Y(n7582) );
  NAND3X1 U7130 ( .A(n4732), .B(n4776), .C(n3640), .Y(n7583) );
  AOI22X1 U7131 ( .A(n8097), .B(n4941), .C(n3360), .D(n5210), .Y(n7589) );
  AOI21X1 U7132 ( .A(n7550), .B(n6295), .C(n2368), .Y(n7610) );
  NAND3X1 U7133 ( .A(n4837), .B(n4774), .C(n3660), .Y(n7616) );
  AOI22X1 U7134 ( .A(n5767), .B(n6303), .C(n7586), .D(n5982), .Y(n7587) );
  AOI22X1 U7135 ( .A(n5759), .B(n7875), .C(n5755), .D(n5116), .Y(n7588) );
  AOI22X1 U7136 ( .A(n5964), .B(n9793), .C(n5961), .D(n6065), .Y(n7594) );
  OAI21X1 U7137 ( .A(n5953), .B(n6091), .C(n6089), .Y(n7591) );
  OAI21X1 U7138 ( .A(n6064), .B(n6293), .C(n5466), .Y(n7864) );
  AOI22X1 U7139 ( .A(n6187), .B(n7591), .C(n5862), .D(n9916), .Y(n7592) );
  NAND3X1 U7140 ( .A(n2427), .B(n3098), .C(n3409), .Y(n7595) );
  AOI21X1 U7141 ( .A(n6308), .B(n6077), .C(n5634), .Y(n7598) );
  OAI21X1 U7142 ( .A(n6311), .B(n6082), .C(n5633), .Y(n8379) );
  OAI21X1 U7143 ( .A(n6311), .B(n6153), .C(n5633), .Y(n8378) );
  OAI21X1 U7144 ( .A(n7600), .B(n5731), .C(n1927), .Y(n8369) );
  AOI21X1 U7145 ( .A(n6083), .B(n6295), .C(n2369), .Y(n7604) );
  OAI21X1 U7146 ( .A(n6296), .B(n6078), .C(n4838), .Y(n7602) );
  AOI22X1 U7147 ( .A(n6731), .B(n8369), .C(n7876), .D(n10375), .Y(n7606) );
  NAND3X1 U7148 ( .A(n4838), .B(n6062), .C(n3661), .Y(n7613) );
  AOI22X1 U7149 ( .A(n8968), .B(n4942), .C(n3531), .D(n6092), .Y(n7605) );
  AOI22X1 U7150 ( .A(n7611), .B(n6308), .C(n7550), .D(n5984), .Y(n7609) );
  AOI22X1 U7151 ( .A(n5767), .B(n10487), .C(n6187), .D(n7491), .Y(n7607) );
  OAI21X1 U7152 ( .A(n5766), .B(n3354), .C(n7608), .Y(n8376) );
  OAI21X1 U7153 ( .A(n5969), .B(n4799), .C(n4837), .Y(n7612) );
  AOI22X1 U7154 ( .A(n7755), .B(n8376), .C(n7748), .D(n7874), .Y(n7619) );
  AOI21X1 U7155 ( .A(n6305), .B(n6079), .C(n8130), .Y(n7614) );
  AOI22X1 U7156 ( .A(n9774), .B(n5071), .C(n7732), .D(n4867), .Y(n7617) );
  NAND3X1 U7157 ( .A(n2428), .B(n3099), .C(n3410), .Y(n7620) );
  MUX2X1 U7158 ( .B(n6090), .A(n6067), .S(n6187), .Y(n7622) );
  NAND3X1 U7159 ( .A(n7622), .B(n6069), .C(n9803), .Y(n7623) );
  MUX2X1 U7160 ( .B(n6088), .A(n5476), .S(n5955), .Y(n7626) );
  AOI22X1 U7161 ( .A(n778), .B(n6137), .C(n5976), .D(n9969), .Y(n7624) );
  NAND3X1 U7162 ( .A(n7626), .B(n3101), .C(n3411), .Y(n7631) );
  AOI22X1 U7163 ( .A(n722), .B(n5790), .C(n2247), .D(n5838), .Y(n7629) );
  AOI22X1 U7164 ( .A(n2889), .B(n5829), .C(n457), .D(n5839), .Y(n7627) );
  NAND3X1 U7165 ( .A(n2429), .B(n3102), .C(n3412), .Y(n7630) );
  AOI22X1 U7166 ( .A(n45), .B(n9500), .C(n6098), .D(n6026), .Y(n7633) );
  AOI22X1 U7167 ( .A(n401), .B(n5778), .C(n569), .D(n5823), .Y(n7632) );
  AOI22X1 U7168 ( .A(n3852), .B(n5828), .C(n3210), .D(n5827), .Y(n7636) );
  AOI22X1 U7169 ( .A(n1292), .B(n6125), .C(n890), .D(n5824), .Y(n7634) );
  NOR3X1 U7170 ( .A(n7638), .B(n4240), .C(n4394), .Y(n7639) );
  NAND3X1 U7171 ( .A(n2725), .B(n3100), .C(n7639), .Y(n7642) );
  AOI22X1 U7172 ( .A(n2952), .B(n6141), .C(n1854), .D(n5783), .Y(n7647) );
  AOI22X1 U7173 ( .A(n1629), .B(n5784), .C(n5916), .D(n10480), .Y(n7646) );
  AOI22X1 U7174 ( .A(n2857), .B(n5780), .C(n2536), .D(n6115), .Y(n7644) );
  NAND3X1 U7175 ( .A(n2430), .B(n3009), .C(n7645), .Y(n7648) );
  AOI22X1 U7176 ( .A(n3821), .B(n5775), .C(n3500), .D(n5774), .Y(n7654) );
  AOI22X1 U7177 ( .A(n1373), .B(n6139), .C(n859), .D(n6145), .Y(n7651) );
  NAND3X1 U7178 ( .A(n2431), .B(n5425), .C(n7652), .Y(n7724) );
  AOI22X1 U7179 ( .A(n5955), .B(n9632), .C(n5952), .D(n9626), .Y(n7655) );
  OAI21X1 U7180 ( .A(n6064), .B(n6294), .C(n1873), .Y(n8418) );
  OAI21X1 U7181 ( .A(n6189), .B(n9846), .C(n5503), .Y(n7985) );
  AOI22X1 U7182 ( .A(n8418), .B(n6072), .C(n7985), .D(n5205), .Y(n7667) );
  NAND3X1 U7183 ( .A(n4734), .B(n4777), .C(n3662), .Y(n7661) );
  MUX2X1 U7184 ( .B(n5967), .A(n6298), .S(n6185), .Y(n7662) );
  AOI22X1 U7185 ( .A(n5980), .B(n9632), .C(n6305), .D(n9626), .Y(n7664) );
  AOI22X1 U7186 ( .A(n5983), .B(n6080), .C(n5977), .D(n6083), .Y(n7663) );
  AOI22X1 U7187 ( .A(n5759), .B(n7691), .C(n8954), .D(n5651), .Y(n7665) );
  NAND3X1 U7188 ( .A(n2432), .B(n3103), .C(n3413), .Y(n7676) );
  AOI22X1 U7189 ( .A(n5767), .B(n6305), .C(n7586), .D(n5983), .Y(n7668) );
  NAND3X1 U7190 ( .A(n7988), .B(n7491), .C(n5191), .Y(n7670) );
  OAI21X1 U7191 ( .A(n9703), .B(n6295), .C(n1901), .Y(n7671) );
  AOI21X1 U7192 ( .A(n5964), .B(n6065), .C(n7671), .Y(n7674) );
  OAI21X1 U7193 ( .A(n5958), .B(n6091), .C(n6089), .Y(n7672) );
  AOI22X1 U7194 ( .A(n5960), .B(n6066), .C(n6189), .D(n7672), .Y(n7673) );
  MUX2X1 U7195 ( .B(n5988), .A(n6308), .S(n9688), .Y(n8174) );
  MUX2X1 U7196 ( .B(n5970), .A(n5969), .S(n9688), .Y(n7677) );
  AOI22X1 U7197 ( .A(n6730), .B(n8426), .C(n10375), .D(n7932), .Y(n7682) );
  MUX2X1 U7198 ( .B(n6296), .A(n5970), .S(n5888), .Y(n7678) );
  AOI21X1 U7199 ( .A(n5973), .B(n9626), .C(n5648), .Y(n7679) );
  OAI21X1 U7200 ( .A(n6062), .B(n6300), .C(n1902), .Y(n7926) );
  AOI22X1 U7201 ( .A(n3532), .B(n6092), .C(n3853), .D(n6096), .Y(n7680) );
  NAND3X1 U7202 ( .A(n2433), .B(n3104), .C(n3414), .Y(n7696) );
  MUX2X1 U7203 ( .B(n6308), .A(n5988), .S(n5886), .Y(n7683) );
  MUX2X1 U7204 ( .B(n5651), .A(n5573), .S(n5890), .Y(n7684) );
  MUX2X1 U7205 ( .B(n6297), .A(n5968), .S(n7550), .Y(n7685) );
  AOI22X1 U7206 ( .A(n8172), .B(n5770), .C(n7748), .D(n7931), .Y(n7694) );
  MUX2X1 U7207 ( .B(n6311), .A(n6309), .S(n7550), .Y(n7686) );
  MUX2X1 U7208 ( .B(n6310), .A(n6311), .S(n6185), .Y(n7687) );
  MUX2X1 U7209 ( .B(n171), .A(n5707), .S(n6189), .Y(n7688) );
  OAI21X1 U7210 ( .A(n6190), .B(n5636), .C(n1928), .Y(n8167) );
  AOI22X1 U7211 ( .A(n5648), .B(n6721), .C(n7732), .D(n4982), .Y(n7692) );
  NAND3X1 U7212 ( .A(n2434), .B(n3105), .C(n3415), .Y(n7695) );
  MUX2X1 U7213 ( .B(n6090), .A(n6067), .S(n6189), .Y(n7697) );
  NAND3X1 U7214 ( .A(n7697), .B(n6069), .C(n9803), .Y(n7698) );
  MUX2X1 U7215 ( .B(n6088), .A(n5337), .S(n5957), .Y(n7701) );
  AOI22X1 U7216 ( .A(n779), .B(n6137), .C(n6301), .D(n9969), .Y(n7699) );
  NAND3X1 U7217 ( .A(n7701), .B(n3107), .C(n3416), .Y(n7706) );
  AOI22X1 U7218 ( .A(n723), .B(n5790), .C(n2248), .D(n6104), .Y(n7704) );
  AOI22X1 U7219 ( .A(n2890), .B(n5829), .C(n458), .D(n6131), .Y(n7702) );
  NAND3X1 U7220 ( .A(n2435), .B(n3108), .C(n3417), .Y(n7705) );
  AOI22X1 U7221 ( .A(n891), .B(n5824), .C(n6296), .D(n9500), .Y(n7709) );
  AOI22X1 U7222 ( .A(n402), .B(n5778), .C(n570), .D(n5823), .Y(n7707) );
  AOI22X1 U7223 ( .A(n3211), .B(n6100), .C(n1775), .D(n6121), .Y(n7712) );
  AOI22X1 U7224 ( .A(n1293), .B(n5785), .C(n1550), .D(n6123), .Y(n7710) );
  NOR3X1 U7225 ( .A(n7713), .B(n4155), .C(n4398), .Y(n7714) );
  NAND3X1 U7226 ( .A(n2726), .B(n3106), .C(n7714), .Y(n7717) );
  AOI22X1 U7227 ( .A(n2953), .B(n6141), .C(n1855), .D(n5783), .Y(n7722) );
  AOI22X1 U7228 ( .A(n1630), .B(n5784), .C(n5918), .D(n10480), .Y(n7721) );
  AOI22X1 U7229 ( .A(n2858), .B(n5780), .C(n2537), .D(n6115), .Y(n7719) );
  NAND3X1 U7230 ( .A(n2436), .B(n3010), .C(n7720), .Y(n7723) );
  AOI22X1 U7231 ( .A(n3822), .B(n5775), .C(n3501), .D(n5774), .Y(n7729) );
  AOI22X1 U7232 ( .A(n1374), .B(n6139), .C(n860), .D(n5771), .Y(n7726) );
  NAND3X1 U7233 ( .A(n2437), .B(n5481), .C(n7727), .Y(n7786) );
  AOI21X1 U7234 ( .A(n6301), .B(n6079), .C(n7978), .Y(n7730) );
  AOI22X1 U7235 ( .A(n8968), .B(n4886), .C(n3533), .D(n6092), .Y(n7743) );
  AOI22X1 U7236 ( .A(n3854), .B(n5828), .C(n3212), .D(n6100), .Y(n7742) );
  AOI21X1 U7237 ( .A(n7586), .B(n6301), .C(n8126), .Y(n7731) );
  NAND3X1 U7238 ( .A(n6191), .B(n5988), .C(n7491), .Y(n8316) );
  OAI21X1 U7239 ( .A(n155), .B(n5569), .C(n4858), .Y(n7740) );
  AOI22X1 U7240 ( .A(n6305), .B(n9632), .C(n5984), .D(n9626), .Y(n7733) );
  AOI22X1 U7241 ( .A(n5767), .B(n5983), .C(n7586), .D(n5987), .Y(n7736) );
  AOI22X1 U7242 ( .A(n5759), .B(n7735), .C(n5755), .D(n5119), .Y(n7738) );
  OAI21X1 U7243 ( .A(n159), .B(n5655), .C(n1874), .Y(n7739) );
  AOI22X1 U7244 ( .A(n5958), .B(n6077), .C(n5955), .D(n6081), .Y(n7745) );
  AOI22X1 U7245 ( .A(n5952), .B(n6079), .C(n5961), .D(n6083), .Y(n7744) );
  AOI22X1 U7246 ( .A(n5767), .B(n5953), .C(n7586), .D(n5952), .Y(n7746) );
  AOI22X1 U7247 ( .A(n5184), .B(n5628), .C(n7985), .D(n5245), .Y(n7754) );
  NAND3X1 U7248 ( .A(n4735), .B(n4778), .C(n3663), .Y(n7751) );
  AOI22X1 U7249 ( .A(n5970), .B(n2777), .C(n3362), .D(n5210), .Y(n7753) );
  OAI21X1 U7250 ( .A(n4754), .B(n5030), .C(n9791), .Y(n7756) );
  AOI22X1 U7251 ( .A(n5989), .B(n7756), .C(n5968), .D(n9793), .Y(n7760) );
  OAI21X1 U7252 ( .A(n5960), .B(n6091), .C(n6089), .Y(n7757) );
  AOI22X1 U7253 ( .A(n5965), .B(n6066), .C(n6191), .D(n7757), .Y(n7758) );
  NOR3X1 U7254 ( .A(n3912), .B(n4241), .C(n4402), .Y(n7778) );
  AOI22X1 U7255 ( .A(n2249), .B(n6104), .C(n2570), .D(n6102), .Y(n7769) );
  AOI22X1 U7256 ( .A(n2891), .B(n5829), .C(n459), .D(n5839), .Y(n7768) );
  AOI22X1 U7257 ( .A(n780), .B(n6137), .C(n6303), .D(n9969), .Y(n7766) );
  MUX2X1 U7258 ( .B(n6091), .A(n6068), .S(n6191), .Y(n7762) );
  NOR3X1 U7259 ( .A(n5728), .B(n9731), .C(n7762), .Y(n7763) );
  MUX2X1 U7260 ( .B(n10522), .A(n7763), .S(n5961), .Y(n7764) );
  AOI21X1 U7261 ( .A(n1117), .B(n5826), .C(n7764), .Y(n7765) );
  NAND3X1 U7262 ( .A(n5541), .B(n5483), .C(n7767), .Y(n7776) );
  AOI22X1 U7263 ( .A(n6098), .B(n6032), .C(n403), .D(n5778), .Y(n7771) );
  AOI22X1 U7264 ( .A(n571), .B(n6135), .C(n724), .D(n5790), .Y(n7770) );
  AOI22X1 U7265 ( .A(n1776), .B(n5777), .C(n1037), .D(n6129), .Y(n7774) );
  AOI22X1 U7266 ( .A(n1551), .B(n5779), .C(n892), .D(n5824), .Y(n7772) );
  NOR3X1 U7267 ( .A(n3916), .B(n4242), .C(n4406), .Y(n7777) );
  AOI22X1 U7268 ( .A(n2979), .B(n6141), .C(n1856), .D(n5783), .Y(n7784) );
  AOI22X1 U7269 ( .A(n1631), .B(n5784), .C(n17), .D(n10480), .Y(n7783) );
  AOI22X1 U7270 ( .A(n2859), .B(n5780), .C(n2538), .D(n6115), .Y(n7781) );
  NAND3X1 U7271 ( .A(n2438), .B(n3011), .C(n7782), .Y(n7785) );
  AOI22X1 U7272 ( .A(n3823), .B(n5775), .C(n3502), .D(n5774), .Y(n7791) );
  AOI22X1 U7273 ( .A(n1375), .B(n6139), .C(n861), .D(n5771), .Y(n7788) );
  NAND3X1 U7274 ( .A(n2439), .B(n3109), .C(n7789), .Y(n7837) );
  AOI22X1 U7275 ( .A(n5755), .B(n5254), .C(n9774), .D(n5215), .Y(n7796) );
  AOI22X1 U7276 ( .A(n7732), .B(n5113), .C(n8968), .D(n5143), .Y(n7795) );
  AOI22X1 U7277 ( .A(n3534), .B(n5830), .C(n3855), .D(n6096), .Y(n7793) );
  AOI22X1 U7278 ( .A(n3213), .B(n5827), .C(n1777), .D(n6121), .Y(n7792) );
  AOI22X1 U7279 ( .A(n5961), .B(n6077), .C(n5957), .D(n6081), .Y(n7797) );
  AOI21X1 U7280 ( .A(n7586), .B(n5955), .C(n7800), .Y(n7801) );
  AOI22X1 U7281 ( .A(n5065), .B(n6072), .C(n7985), .D(n5122), .Y(n7807) );
  OAI21X1 U7282 ( .A(n9846), .B(n6190), .C(n5501), .Y(n7980) );
  AOI22X1 U7283 ( .A(n5744), .B(n7980), .C(n5210), .D(n4963), .Y(n7806) );
  OAI21X1 U7284 ( .A(n10375), .B(n7748), .C(n6297), .Y(n7808) );
  NAND3X1 U7285 ( .A(n2727), .B(n4858), .C(n7808), .Y(n7860) );
  OAI21X1 U7286 ( .A(n5965), .B(n6091), .C(n6089), .Y(n7811) );
  AOI22X1 U7287 ( .A(n6193), .B(n7811), .C(n4952), .D(n6073), .Y(n7812) );
  NOR3X1 U7288 ( .A(n3917), .B(n4243), .C(n4410), .Y(n7829) );
  AOI22X1 U7289 ( .A(n1038), .B(n5786), .C(n1295), .D(n5785), .Y(n7819) );
  AOI22X1 U7290 ( .A(n1552), .B(n5779), .C(n893), .D(n6133), .Y(n7818) );
  AOI22X1 U7291 ( .A(n6098), .B(n5885), .C(n404), .D(n6117), .Y(n7816) );
  AOI22X1 U7292 ( .A(n572), .B(n6135), .C(n725), .D(n5790), .Y(n7815) );
  MUX2X1 U7293 ( .B(n6090), .A(n6067), .S(n6193), .Y(n7820) );
  MUX2X1 U7294 ( .B(n6088), .A(n5291), .S(n5965), .Y(n7824) );
  AOI22X1 U7295 ( .A(n781), .B(n6137), .C(n6305), .D(n9969), .Y(n7822) );
  AOI22X1 U7296 ( .A(n2250), .B(n6104), .C(n2571), .D(n5831), .Y(n7826) );
  AOI22X1 U7297 ( .A(n2892), .B(n5829), .C(n460), .D(n5839), .Y(n7825) );
  NOR3X1 U7298 ( .A(n3922), .B(n4159), .C(n4598), .Y(n7828) );
  AOI22X1 U7299 ( .A(n2980), .B(n6141), .C(n1857), .D(n5783), .Y(n7835) );
  AOI22X1 U7300 ( .A(n1632), .B(n5784), .C(n67), .D(n10480), .Y(n7834) );
  AOI22X1 U7301 ( .A(n2860), .B(n5780), .C(n2539), .D(n6115), .Y(n7832) );
  NAND3X1 U7302 ( .A(n2440), .B(n3012), .C(n7833), .Y(n7836) );
  AOI22X1 U7303 ( .A(n3824), .B(n5775), .C(n3503), .D(n5774), .Y(n7842) );
  AOI22X1 U7304 ( .A(n1376), .B(n6139), .C(n862), .D(n5771), .Y(n7839) );
  NAND3X1 U7305 ( .A(n2441), .B(n3110), .C(n7840), .Y(n7902) );
  AOI22X1 U7306 ( .A(n5955), .B(n9500), .C(n6098), .D(n6034), .Y(n7844) );
  AOI22X1 U7307 ( .A(n405), .B(n5778), .C(n573), .D(n5823), .Y(n7843) );
  AOI22X1 U7308 ( .A(n1778), .B(n5777), .C(n1039), .D(n5786), .Y(n7847) );
  AOI22X1 U7309 ( .A(n1553), .B(n5779), .C(n894), .D(n5824), .Y(n7845) );
  NAND3X1 U7310 ( .A(n2442), .B(n5612), .C(n3418), .Y(n7848) );
  MUX2X1 U7311 ( .B(n6090), .A(n6067), .S(n6195), .Y(n7850) );
  MUX2X1 U7312 ( .B(n6088), .A(n5303), .S(n5966), .Y(n7854) );
  AOI22X1 U7313 ( .A(n782), .B(n6137), .C(n5984), .D(n9969), .Y(n7852) );
  NAND3X1 U7314 ( .A(n7854), .B(n5439), .C(n3419), .Y(n7859) );
  AOI22X1 U7315 ( .A(n726), .B(n5790), .C(n2251), .D(n6104), .Y(n7857) );
  AOI22X1 U7316 ( .A(n2893), .B(n5829), .C(n461), .D(n5839), .Y(n7855) );
  NAND3X1 U7317 ( .A(n2443), .B(n3111), .C(n3420), .Y(n7858) );
  OAI21X1 U7318 ( .A(n5966), .B(n6091), .C(n6089), .Y(n7861) );
  AOI21X1 U7319 ( .A(n6195), .B(n7861), .C(n4718), .Y(n7882) );
  AOI22X1 U7320 ( .A(n5965), .B(n6077), .C(n5960), .D(n6081), .Y(n7863) );
  AOI22X1 U7321 ( .A(n5958), .B(n6079), .C(n5966), .D(n6083), .Y(n7862) );
  MUX2X1 U7322 ( .B(n8127), .A(n7865), .S(n5889), .Y(n8356) );
  AOI21X1 U7323 ( .A(n7550), .B(n5966), .C(n5810), .Y(n7866) );
  MUX2X1 U7324 ( .B(n4903), .A(n5705), .S(n6189), .Y(n7870) );
  AOI22X1 U7325 ( .A(n8356), .B(n9916), .C(n8363), .D(n4941), .Y(n7881) );
  AOI22X1 U7326 ( .A(n7875), .B(n7872), .C(n7874), .D(n7873), .Y(n7879) );
  AOI22X1 U7327 ( .A(n7877), .B(n5822), .C(n7876), .D(n7147), .Y(n7878) );
  AOI22X1 U7328 ( .A(n8968), .B(n5071), .C(n3535), .D(n6092), .Y(n7884) );
  AOI22X1 U7329 ( .A(n3856), .B(n5828), .C(n3214), .D(n6100), .Y(n7883) );
  AOI22X1 U7330 ( .A(n7988), .B(n8376), .C(n7732), .D(n5116), .Y(n7890) );
  AOI22X1 U7331 ( .A(n5833), .B(n8369), .C(n6791), .D(n4942), .Y(n7888) );
  NOR3X1 U7332 ( .A(n3927), .B(n4244), .C(n4413), .Y(n7892) );
  NAND3X1 U7333 ( .A(n2728), .B(n3112), .C(n7892), .Y(n7895) );
  AOI22X1 U7334 ( .A(n2954), .B(n6141), .C(n1858), .D(n5783), .Y(n7900) );
  AOI22X1 U7335 ( .A(n1633), .B(n5784), .C(n5924), .D(n10480), .Y(n7899) );
  AOI22X1 U7336 ( .A(n2861), .B(n5780), .C(n2540), .D(n6115), .Y(n7897) );
  NAND3X1 U7337 ( .A(n2444), .B(n3013), .C(n7898), .Y(n7901) );
  AOI22X1 U7338 ( .A(n3825), .B(n5775), .C(n3504), .D(n5774), .Y(n7907) );
  AOI22X1 U7339 ( .A(n1377), .B(n6139), .C(n863), .D(n5771), .Y(n7904) );
  NAND3X1 U7340 ( .A(n2445), .B(n3113), .C(n7905), .Y(n7965) );
  AOI22X1 U7341 ( .A(n1554), .B(n5779), .C(n895), .D(n6133), .Y(n7910) );
  AOI22X1 U7342 ( .A(n6098), .B(n6037), .C(n406), .D(n6117), .Y(n7908) );
  NAND3X1 U7343 ( .A(n2446), .B(n3114), .C(n3421), .Y(n7915) );
  AOI22X1 U7344 ( .A(n3857), .B(n5828), .C(n3215), .D(n5827), .Y(n7913) );
  AOI22X1 U7345 ( .A(n1040), .B(n5786), .C(n1297), .D(n5785), .Y(n7911) );
  NAND3X1 U7346 ( .A(n5531), .B(n5676), .C(n5621), .Y(n7914) );
  AOI22X1 U7347 ( .A(n574), .B(n6135), .C(n727), .D(n5790), .Y(n7918) );
  AOI22X1 U7348 ( .A(n2573), .B(n6102), .C(n2894), .D(n5829), .Y(n7916) );
  MUX2X1 U7349 ( .B(n6090), .A(n6067), .S(n6197), .Y(n7919) );
  MUX2X1 U7350 ( .B(n5832), .A(n5539), .S(n6296), .Y(n7922) );
  AOI22X1 U7351 ( .A(n462), .B(n5839), .C(n783), .D(n6137), .Y(n7923) );
  OAI21X1 U7352 ( .A(n6095), .B(n6309), .C(n5408), .Y(n7924) );
  NOR3X1 U7353 ( .A(n3932), .B(n4245), .C(n7924), .Y(n7956) );
  AOI22X1 U7354 ( .A(n7732), .B(n5191), .C(n7885), .D(n4982), .Y(n7929) );
  AOI22X1 U7355 ( .A(n8968), .B(n5651), .C(n3536), .D(n6092), .Y(n7927) );
  NAND3X1 U7356 ( .A(n2447), .B(n3115), .C(n3422), .Y(n7938) );
  AOI22X1 U7357 ( .A(n5861), .B(n5770), .C(n7691), .D(n7872), .Y(n7936) );
  AOI22X1 U7358 ( .A(n5648), .B(n5822), .C(n7147), .D(n7932), .Y(n7934) );
  NAND3X1 U7359 ( .A(n2448), .B(n3116), .C(n3423), .Y(n7937) );
  AOI22X1 U7360 ( .A(n5960), .B(n6079), .C(n5969), .D(n6083), .Y(n7939) );
  AOI22X1 U7361 ( .A(n7980), .B(n5205), .C(n5101), .D(n6072), .Y(n7949) );
  AOI21X1 U7362 ( .A(n7550), .B(n6296), .C(n7942), .Y(n7943) );
  AOI22X1 U7363 ( .A(n7946), .B(n7988), .C(n8954), .D(n8426), .Y(n7947) );
  NAND3X1 U7364 ( .A(n6191), .B(n10487), .C(n5806), .Y(n7953) );
  OAI21X1 U7365 ( .A(n5968), .B(n6091), .C(n6089), .Y(n7951) );
  AOI22X1 U7366 ( .A(n6197), .B(n7951), .C(n8418), .D(n10574), .Y(n7952) );
  NOR3X1 U7367 ( .A(n7954), .B(n4163), .C(n4417), .Y(n7955) );
  NAND3X1 U7368 ( .A(n2729), .B(n7956), .C(n7955), .Y(n7958) );
  AOI22X1 U7369 ( .A(n2955), .B(n6141), .C(n1859), .D(n5783), .Y(n7963) );
  AOI22X1 U7370 ( .A(n1634), .B(n5784), .C(n5926), .D(n10480), .Y(n7962) );
  AOI22X1 U7371 ( .A(n2862), .B(n5780), .C(n2541), .D(n6115), .Y(n7960) );
  NAND3X1 U7372 ( .A(n2449), .B(n3014), .C(n7961), .Y(n7964) );
  AOI22X1 U7373 ( .A(n3826), .B(n5775), .C(n3505), .D(n5774), .Y(n7970) );
  AOI22X1 U7374 ( .A(n1378), .B(n6139), .C(n864), .D(n5771), .Y(n7967) );
  NAND3X1 U7375 ( .A(n2450), .B(n3117), .C(n7968), .Y(n8016) );
  AOI22X1 U7376 ( .A(n7732), .B(n5119), .C(n7885), .D(n4811), .Y(n7976) );
  AOI22X1 U7377 ( .A(n6791), .B(n4886), .C(n8968), .D(n5016), .Y(n7975) );
  AOI22X1 U7378 ( .A(n3537), .B(n5830), .C(n3858), .D(n6096), .Y(n7973) );
  AOI22X1 U7379 ( .A(n3216), .B(n5827), .C(n1780), .D(n6121), .Y(n7972) );
  AOI22X1 U7380 ( .A(n5969), .B(n6077), .C(n45), .D(n6081), .Y(n7977) );
  AOI22X1 U7381 ( .A(n7980), .B(n5245), .C(n5152), .D(n5628), .Y(n7987) );
  AOI21X1 U7382 ( .A(n7611), .B(n6296), .C(n7735), .Y(n7981) );
  AOI22X1 U7383 ( .A(n7985), .B(n5083), .C(n7735), .D(n7872), .Y(n7986) );
  OAI21X1 U7384 ( .A(n4755), .B(n5030), .C(n10033), .Y(n7989) );
  OAI21X1 U7385 ( .A(n5970), .B(n6091), .C(n6089), .Y(n7990) );
  AOI22X1 U7386 ( .A(n6199), .B(n7990), .C(n5184), .D(n10574), .Y(n7991) );
  NOR3X1 U7387 ( .A(n3936), .B(n4246), .C(n4421), .Y(n8008) );
  AOI22X1 U7388 ( .A(n1041), .B(n5786), .C(n1298), .D(n5785), .Y(n7998) );
  AOI22X1 U7389 ( .A(n1555), .B(n5779), .C(n896), .D(n6133), .Y(n7997) );
  AOI22X1 U7390 ( .A(n5960), .B(n9500), .C(n6098), .D(n6039), .Y(n7995) );
  AOI22X1 U7391 ( .A(n407), .B(n5778), .C(n575), .D(n5823), .Y(n7994) );
  MUX2X1 U7392 ( .B(n6090), .A(n6067), .S(n6199), .Y(n7999) );
  MUX2X1 U7393 ( .B(n5832), .A(n2938), .S(n5970), .Y(n8003) );
  AOI22X1 U7394 ( .A(n463), .B(n5839), .C(n784), .D(n5825), .Y(n8001) );
  AOI22X1 U7395 ( .A(n728), .B(n5790), .C(n2253), .D(n6104), .Y(n8005) );
  AOI22X1 U7396 ( .A(n2574), .B(n6102), .C(n2895), .D(n6086), .Y(n8004) );
  NOR3X1 U7397 ( .A(n3941), .B(n4167), .C(n4599), .Y(n8007) );
  AOI22X1 U7398 ( .A(n2981), .B(n6141), .C(n1860), .D(n5783), .Y(n8014) );
  AOI22X1 U7399 ( .A(n1635), .B(n6147), .C(n5929), .D(n6112), .Y(n8013) );
  AOI22X1 U7400 ( .A(n2863), .B(n5780), .C(n2542), .D(n6115), .Y(n8011) );
  NAND3X1 U7401 ( .A(n125), .B(n3015), .C(n8012), .Y(n8015) );
  AOI22X1 U7402 ( .A(n3827), .B(n5775), .C(n3506), .D(n5774), .Y(n8021) );
  AOI22X1 U7403 ( .A(n1379), .B(n6139), .C(n865), .D(n5771), .Y(n8018) );
  NAND3X1 U7404 ( .A(n2451), .B(n5543), .C(n8019), .Y(n8073) );
  AOI21X1 U7405 ( .A(n45), .B(n6079), .C(n8022), .Y(n8023) );
  AOI22X1 U7406 ( .A(n5951), .B(n10072), .C(n6625), .D(n4984), .Y(n8034) );
  AOI21X1 U7407 ( .A(n7611), .B(n5970), .C(n8026), .Y(n8027) );
  AOI22X1 U7408 ( .A(n10500), .B(n5065), .C(n7656), .D(n4915), .Y(n8033) );
  AOI22X1 U7409 ( .A(n3538), .B(n5830), .C(n3859), .D(n6096), .Y(n8031) );
  AOI22X1 U7410 ( .A(n3217), .B(n6100), .C(n1781), .D(n6121), .Y(n8030) );
  AOI22X1 U7411 ( .A(n5744), .B(n5796), .C(n7732), .D(n5254), .Y(n8037) );
  AOI22X1 U7412 ( .A(n8035), .B(n5122), .C(n7885), .D(n5113), .Y(n8036) );
  OAI21X1 U7413 ( .A(n5974), .B(n6091), .C(n6089), .Y(n8038) );
  OAI21X1 U7414 ( .A(n6311), .B(n5729), .C(n5518), .Y(n8175) );
  AOI21X1 U7415 ( .A(n6201), .B(n8038), .C(n8175), .Y(n8047) );
  OAI21X1 U7416 ( .A(n6304), .B(n5726), .C(n5596), .Y(n8040) );
  AOI21X1 U7417 ( .A(n8102), .B(n5975), .C(n8040), .Y(n8043) );
  AOI22X1 U7418 ( .A(n5787), .B(n6308), .C(n8163), .D(n5988), .Y(n8042) );
  AOI22X1 U7419 ( .A(n8102), .B(n5984), .C(n8299), .D(n5981), .Y(n8041) );
  MUX2X1 U7420 ( .B(n2766), .A(n8324), .S(n6205), .Y(n8044) );
  AOI22X1 U7421 ( .A(n5143), .B(n6073), .C(n8044), .D(n5733), .Y(n8045) );
  NOR3X1 U7422 ( .A(n3946), .B(n4247), .C(n4424), .Y(n8065) );
  AOI22X1 U7423 ( .A(n1042), .B(n5786), .C(n1299), .D(n5785), .Y(n8053) );
  AOI22X1 U7424 ( .A(n1556), .B(n5779), .C(n897), .D(n5824), .Y(n8052) );
  AOI22X1 U7425 ( .A(n6305), .B(n9500), .C(n6042), .D(n10502), .Y(n8050) );
  AOI22X1 U7426 ( .A(n392), .B(n5778), .C(n576), .D(n5823), .Y(n8049) );
  NAND3X1 U7427 ( .A(n8299), .B(n5589), .C(n6206), .Y(n8054) );
  MUX2X1 U7428 ( .B(n6091), .A(n6068), .S(n6201), .Y(n8055) );
  AOI21X1 U7429 ( .A(n8156), .B(n8299), .C(n8055), .Y(n8056) );
  NAND3X1 U7430 ( .A(n8497), .B(n6085), .C(n3641), .Y(n8057) );
  MUX2X1 U7431 ( .B(n5832), .A(n2792), .S(n5974), .Y(n8060) );
  AOI22X1 U7432 ( .A(n464), .B(n5839), .C(n785), .D(n6137), .Y(n8058) );
  AOI22X1 U7433 ( .A(n713), .B(n5790), .C(n2254), .D(n5838), .Y(n8062) );
  AOI22X1 U7434 ( .A(n2575), .B(n6102), .C(n2896), .D(n5829), .Y(n8061) );
  NOR3X1 U7435 ( .A(n3951), .B(n4171), .C(n4600), .Y(n8064) );
  AOI22X1 U7436 ( .A(n2982), .B(n6141), .C(n1861), .D(n5783), .Y(n8071) );
  AOI22X1 U7437 ( .A(n1636), .B(n6147), .C(n5932), .D(n10480), .Y(n8070) );
  AOI22X1 U7438 ( .A(n2864), .B(n6110), .C(n2543), .D(n6115), .Y(n8068) );
  NAND3X1 U7439 ( .A(n2452), .B(n3016), .C(n8069), .Y(n8072) );
  AOI22X1 U7440 ( .A(n3828), .B(n5775), .C(n3507), .D(n5774), .Y(n8078) );
  AOI22X1 U7441 ( .A(n1380), .B(n6139), .C(n866), .D(n5771), .Y(n8075) );
  NAND3X1 U7442 ( .A(n2453), .B(n3118), .C(n8076), .Y(n8148) );
  AOI22X1 U7443 ( .A(n898), .B(n5824), .C(n5983), .D(n9500), .Y(n8081) );
  AOI22X1 U7444 ( .A(n393), .B(n5778), .C(n577), .D(n5823), .Y(n8079) );
  NAND3X1 U7445 ( .A(n2454), .B(n3119), .C(n3424), .Y(n8086) );
  AOI22X1 U7446 ( .A(n3218), .B(n5827), .C(n1782), .D(n6121), .Y(n8084) );
  AOI22X1 U7447 ( .A(n1300), .B(n5785), .C(n1557), .D(n6123), .Y(n8082) );
  NAND3X1 U7448 ( .A(n2455), .B(n5608), .C(n5383), .Y(n8085) );
  MUX2X1 U7449 ( .B(n6090), .A(n6067), .S(n6203), .Y(n8087) );
  MUX2X1 U7450 ( .B(n5832), .A(n5310), .S(n5976), .Y(n8091) );
  AOI22X1 U7451 ( .A(n786), .B(n5825), .C(n5953), .D(n9969), .Y(n8089) );
  NAND3X1 U7452 ( .A(n8091), .B(n3120), .C(n3425), .Y(n8096) );
  AOI22X1 U7453 ( .A(n714), .B(n5790), .C(n2255), .D(n5838), .Y(n8094) );
  AOI22X1 U7454 ( .A(n2897), .B(n5829), .C(n465), .D(n5839), .Y(n8092) );
  NAND3X1 U7455 ( .A(n2456), .B(n3121), .C(n3426), .Y(n8095) );
  AOI21X1 U7456 ( .A(n5787), .B(n6303), .C(n8244), .Y(n8098) );
  OAI21X1 U7457 ( .A(n6306), .B(n5726), .C(n1903), .Y(n8113) );
  NAND3X1 U7458 ( .A(n5974), .B(n5819), .C(n8102), .Y(n8099) );
  OAI21X1 U7459 ( .A(n10104), .B(n4801), .C(n1904), .Y(n8100) );
  AOI21X1 U7460 ( .A(n10291), .B(n8113), .C(n8100), .Y(n8108) );
  AOI21X1 U7461 ( .A(n8299), .B(n6307), .C(n2370), .Y(n8105) );
  OAI21X1 U7462 ( .A(n6308), .B(n4800), .C(n4839), .Y(n8103) );
  NAND3X1 U7463 ( .A(n4839), .B(n5726), .C(n3664), .Y(n8106) );
  AOI22X1 U7464 ( .A(n8377), .B(n10290), .C(n8375), .D(n10291), .Y(n8107) );
  MUX2X1 U7465 ( .B(n2767), .A(n2783), .S(n6205), .Y(n8109) );
  NOR3X1 U7466 ( .A(n4122), .B(n8109), .C(n8175), .Y(n8122) );
  OAI21X1 U7467 ( .A(n5976), .B(n6091), .C(n6089), .Y(n8111) );
  AOI22X1 U7468 ( .A(n6203), .B(n8111), .C(n5071), .D(n6073), .Y(n8121) );
  OAI21X1 U7469 ( .A(n8112), .B(n8113), .C(n8156), .Y(n8114) );
  OAI21X1 U7470 ( .A(n8116), .B(n5699), .C(n8114), .Y(n8117) );
  AOI21X1 U7471 ( .A(n5862), .B(n5791), .C(n8117), .Y(n8119) );
  AOI22X1 U7472 ( .A(n6721), .B(n8379), .C(n8035), .D(n4903), .Y(n8118) );
  NAND3X1 U7473 ( .A(n8122), .B(n3017), .C(n8120), .Y(n8137) );
  AOI21X1 U7474 ( .A(n5767), .B(n6297), .C(n8123), .Y(n8124) );
  AOI22X1 U7475 ( .A(n10500), .B(n4763), .C(n7656), .D(n4987), .Y(n8129) );
  AOI22X1 U7476 ( .A(n3539), .B(n5830), .C(n3860), .D(n5828), .Y(n8128) );
  AOI22X1 U7477 ( .A(n7885), .B(n5116), .C(n5834), .D(n8369), .Y(n8135) );
  AOI21X1 U7478 ( .A(n6297), .B(n9626), .C(n5712), .Y(n8132) );
  OAI21X1 U7479 ( .A(n6062), .B(n5967), .C(n1905), .Y(n8370) );
  AOI22X1 U7480 ( .A(n6625), .B(n8370), .C(n10375), .D(n8378), .Y(n8133) );
  NOR3X1 U7481 ( .A(n3956), .B(n4248), .C(n4428), .Y(n8138) );
  NAND3X1 U7482 ( .A(n2730), .B(n3122), .C(n8138), .Y(n8141) );
  AOI22X1 U7483 ( .A(n2956), .B(n6141), .C(n1862), .D(n5783), .Y(n8146) );
  AOI22X1 U7484 ( .A(n1637), .B(n5784), .C(n5934), .D(n10480), .Y(n8145) );
  AOI22X1 U7485 ( .A(n2865), .B(n5780), .C(n2544), .D(n6115), .Y(n8143) );
  NAND3X1 U7486 ( .A(n2457), .B(n3018), .C(n8144), .Y(n8147) );
  AOI22X1 U7487 ( .A(n3829), .B(n5775), .C(n3508), .D(n6106), .Y(n8153) );
  AOI22X1 U7488 ( .A(n1381), .B(n6139), .C(n867), .D(n6145), .Y(n8150) );
  NAND3X1 U7489 ( .A(n2458), .B(n3123), .C(n8151), .Y(n8222) );
  AOI22X1 U7490 ( .A(n5787), .B(n6305), .C(n8163), .D(n5984), .Y(n8155) );
  AOI22X1 U7491 ( .A(n8102), .B(n6303), .C(n8299), .D(n6301), .Y(n8154) );
  MUX2X1 U7492 ( .B(n5989), .A(n6308), .S(n8299), .Y(n8157) );
  MUX2X1 U7493 ( .B(n6308), .A(n5989), .S(n6201), .Y(n8158) );
  AOI22X1 U7494 ( .A(n5709), .B(n10291), .C(n6090), .D(n6302), .Y(n8159) );
  NAND3X1 U7495 ( .A(n2731), .B(n6089), .C(n3427), .Y(n8161) );
  AOI22X1 U7496 ( .A(n2983), .B(n5104), .C(n6205), .D(n3372), .Y(n8170) );
  NAND3X1 U7497 ( .A(n2732), .B(n3124), .C(n5726), .Y(n8166) );
  AOI21X1 U7498 ( .A(n8299), .B(n6302), .C(n2346), .Y(n8419) );
  AOI22X1 U7499 ( .A(n4900), .B(n8300), .C(n8167), .D(n6192), .Y(n8168) );
  OAI21X1 U7500 ( .A(n8171), .B(n8174), .C(n1929), .Y(n8179) );
  NAND3X1 U7501 ( .A(n5799), .B(n7491), .C(n5191), .Y(n8178) );
  NOR3X1 U7502 ( .A(n3957), .B(n8179), .C(n4432), .Y(n8214) );
  AOI22X1 U7503 ( .A(n7656), .B(n4918), .C(n3540), .D(n6092), .Y(n8186) );
  AOI22X1 U7504 ( .A(n3861), .B(n5828), .C(n3219), .D(n6100), .Y(n8185) );
  AOI22X1 U7505 ( .A(n8035), .B(n5056), .C(n7172), .D(n8418), .Y(n8192) );
  AOI22X1 U7506 ( .A(n5887), .B(n6300), .C(shift_amount[3]), .D(n6299), .Y(
        n8187) );
  AOI22X1 U7507 ( .A(n6625), .B(n4943), .C(n10500), .D(n5101), .Y(n8190) );
  NAND3X1 U7508 ( .A(n2459), .B(n3125), .C(n3428), .Y(n8193) );
  MUX2X1 U7509 ( .B(n6090), .A(n6067), .S(n6205), .Y(n8195) );
  MUX2X1 U7510 ( .B(n5832), .A(n5376), .S(n5978), .Y(n8199) );
  AOI22X1 U7511 ( .A(n787), .B(n5825), .C(n5957), .D(n9969), .Y(n8197) );
  NAND3X1 U7512 ( .A(n8199), .B(n3127), .C(n3429), .Y(n8204) );
  AOI22X1 U7513 ( .A(n715), .B(n6119), .C(n2256), .D(n6104), .Y(n8202) );
  AOI22X1 U7514 ( .A(n2898), .B(n5829), .C(n466), .D(n5839), .Y(n8200) );
  NAND3X1 U7515 ( .A(n2460), .B(n3128), .C(n3430), .Y(n8203) );
  AOI22X1 U7516 ( .A(n6308), .B(n9500), .C(n21), .D(n10502), .Y(n8206) );
  AOI22X1 U7517 ( .A(n394), .B(n5778), .C(n578), .D(n5823), .Y(n8205) );
  AOI22X1 U7518 ( .A(n1783), .B(n5777), .C(n1044), .D(n6129), .Y(n8209) );
  AOI22X1 U7519 ( .A(n1558), .B(n5779), .C(n899), .D(n5824), .Y(n8207) );
  NOR3X1 U7520 ( .A(n8211), .B(n4249), .C(n4435), .Y(n8212) );
  NAND3X1 U7521 ( .A(n8214), .B(n3126), .C(n8212), .Y(n8215) );
  AOI22X1 U7522 ( .A(n2957), .B(n6141), .C(n1863), .D(n5783), .Y(n8220) );
  AOI22X1 U7523 ( .A(n1638), .B(n5784), .C(n5938), .D(n6112), .Y(n8219) );
  AOI22X1 U7524 ( .A(n2866), .B(n5780), .C(n2545), .D(n6115), .Y(n8217) );
  NAND3X1 U7525 ( .A(n2461), .B(n3019), .C(n8218), .Y(n8221) );
  AOI22X1 U7526 ( .A(n3830), .B(n6108), .C(n3509), .D(n6106), .Y(n8227) );
  AOI22X1 U7527 ( .A(n1382), .B(n6139), .C(n868), .D(n6145), .Y(n8224) );
  AND2X2 U7528 ( .A(n332), .B(n1671), .Y(n8225) );
  NAND3X1 U7529 ( .A(n2462), .B(n3257), .C(n8225), .Y(n8286) );
  AOI22X1 U7530 ( .A(n8035), .B(n5083), .C(n7885), .D(n5119), .Y(n8237) );
  AOI22X1 U7531 ( .A(n7172), .B(n5184), .C(n10500), .D(n5152), .Y(n8236) );
  AOI22X1 U7532 ( .A(n7656), .B(n4889), .C(n3541), .D(n6092), .Y(n8234) );
  AOI22X1 U7533 ( .A(n3862), .B(n5828), .C(n3220), .D(n6100), .Y(n8233) );
  OAI21X1 U7534 ( .A(n5656), .B(n5514), .C(n5588), .Y(n8242) );
  NAND3X1 U7535 ( .A(n2733), .B(n5444), .C(n5756), .Y(n8241) );
  AOI22X1 U7536 ( .A(n5761), .B(n8242), .C(n5989), .D(n3373), .Y(n8246) );
  AOI22X1 U7537 ( .A(n5787), .B(n5976), .C(n8163), .D(n5973), .Y(n8243) );
  AOI22X1 U7538 ( .A(n5796), .B(n5245), .C(n8300), .D(n4921), .Y(n8245) );
  OAI21X1 U7539 ( .A(n6303), .B(n6091), .C(n6089), .Y(n8248) );
  AOI21X1 U7540 ( .A(n6207), .B(n8248), .C(n8247), .Y(n8260) );
  NAND3X1 U7541 ( .A(n4733), .B(n8252), .C(n4969), .Y(n8483) );
  AOI22X1 U7542 ( .A(n5787), .B(n5983), .C(n8163), .D(n5986), .Y(n8254) );
  NAND3X1 U7543 ( .A(n2734), .B(n4779), .C(n3431), .Y(n8257) );
  AOI22X1 U7544 ( .A(n4901), .B(n5628), .C(n3363), .D(n5104), .Y(n8258) );
  NOR3X1 U7545 ( .A(n3961), .B(n4250), .C(n4439), .Y(n8278) );
  AOI22X1 U7546 ( .A(n2257), .B(n5838), .C(n2578), .D(n6102), .Y(n8269) );
  AOI22X1 U7547 ( .A(n2899), .B(n5829), .C(n467), .D(n5839), .Y(n8268) );
  AOI22X1 U7548 ( .A(n788), .B(n5825), .C(n5961), .D(n9969), .Y(n8266) );
  MUX2X1 U7549 ( .B(n6091), .A(n6068), .S(n6207), .Y(n8262) );
  MUX2X1 U7550 ( .B(n10522), .A(n2939), .S(n5980), .Y(n8264) );
  AOI21X1 U7551 ( .A(n1125), .B(n5826), .C(n8264), .Y(n8265) );
  NAND3X1 U7552 ( .A(n2463), .B(n3020), .C(n8267), .Y(n8276) );
  AOI22X1 U7553 ( .A(n6098), .B(n6351), .C(n395), .D(n6117), .Y(n8271) );
  AOI22X1 U7554 ( .A(n579), .B(n6135), .C(n716), .D(n5790), .Y(n8270) );
  AOI22X1 U7555 ( .A(n1784), .B(n5777), .C(n1045), .D(n5786), .Y(n8274) );
  AOI22X1 U7556 ( .A(n1559), .B(n5779), .C(n900), .D(n5824), .Y(n8272) );
  NOR3X1 U7557 ( .A(n3966), .B(n4251), .C(n4443), .Y(n8277) );
  AOI22X1 U7558 ( .A(n2984), .B(n6141), .C(n1864), .D(n5783), .Y(n8284) );
  AOI22X1 U7559 ( .A(n1639), .B(n5784), .C(n5941), .D(n6112), .Y(n8283) );
  AOI22X1 U7560 ( .A(n2867), .B(n5780), .C(n2546), .D(n6115), .Y(n8281) );
  NAND3X1 U7561 ( .A(n2465), .B(n3021), .C(n8282), .Y(n8285) );
  AOI22X1 U7562 ( .A(n3831), .B(n6108), .C(n3510), .D(n6106), .Y(n8291) );
  AOI22X1 U7563 ( .A(n1383), .B(n5772), .C(n869), .D(n5771), .Y(n8288) );
  AND2X2 U7564 ( .A(n338), .B(n1673), .Y(n8289) );
  NAND3X1 U7565 ( .A(n2466), .B(n3258), .C(n8289), .Y(n8349) );
  AOI22X1 U7566 ( .A(n901), .B(n5824), .C(n6055), .D(n10502), .Y(n8293) );
  AOI22X1 U7567 ( .A(n396), .B(n5778), .C(n580), .D(n5823), .Y(n8292) );
  AOI22X1 U7568 ( .A(n3221), .B(n5827), .C(n1785), .D(n5777), .Y(n8296) );
  AOI22X1 U7569 ( .A(n1303), .B(n5785), .C(n1560), .D(n6123), .Y(n8294) );
  NAND3X1 U7570 ( .A(n2467), .B(n3259), .C(n3432), .Y(n8297) );
  OAI21X1 U7571 ( .A(n5443), .B(n5514), .C(n5732), .Y(n8301) );
  MUX2X1 U7572 ( .B(n6090), .A(n6067), .S(n6209), .Y(n8302) );
  NAND3X1 U7573 ( .A(n8435), .B(n8302), .C(n8433), .Y(n8303) );
  MUX2X1 U7574 ( .B(n5832), .A(n2793), .S(n5981), .Y(n8306) );
  AOI22X1 U7575 ( .A(n789), .B(n5825), .C(n5965), .D(n9969), .Y(n8304) );
  NAND3X1 U7576 ( .A(n8306), .B(n3260), .C(n3433), .Y(n8311) );
  AOI22X1 U7577 ( .A(n717), .B(n5790), .C(n2258), .D(n6104), .Y(n8309) );
  AOI22X1 U7578 ( .A(n2900), .B(n5829), .C(n468), .D(n5839), .Y(n8307) );
  NAND3X1 U7579 ( .A(n2468), .B(n3261), .C(n3434), .Y(n8310) );
  AOI21X1 U7580 ( .A(n8102), .B(n8300), .C(n5749), .Y(n8312) );
  OAI21X1 U7581 ( .A(n8314), .B(n5654), .C(n5988), .Y(n8317) );
  AOI22X1 U7582 ( .A(n5761), .B(n10290), .C(n10375), .D(n5989), .Y(n8315) );
  NAND3X1 U7583 ( .A(n8317), .B(n5518), .C(n3435), .Y(n8361) );
  AOI21X1 U7584 ( .A(n6303), .B(n5229), .C(n4720), .Y(n8331) );
  AOI21X1 U7585 ( .A(n5787), .B(n8300), .C(n5751), .Y(n8318) );
  AOI21X1 U7586 ( .A(n8163), .B(n8300), .C(n5750), .Y(n8320) );
  AOI22X1 U7587 ( .A(n6301), .B(n5248), .C(n5975), .D(n5251), .Y(n8330) );
  OAI21X1 U7588 ( .A(n6305), .B(n6091), .C(n6089), .Y(n8322) );
  AOI22X1 U7589 ( .A(n5973), .B(n2778), .C(n6209), .D(n8322), .Y(n8328) );
  AOI22X1 U7590 ( .A(n5215), .B(n6073), .C(n5104), .D(n4827), .Y(n8327) );
  AOI22X1 U7591 ( .A(n7172), .B(n5065), .C(n10500), .D(n4984), .Y(n8333) );
  AOI22X1 U7592 ( .A(n3542), .B(n5830), .C(n3863), .D(n5828), .Y(n8332) );
  AOI22X1 U7593 ( .A(n5744), .B(n5802), .C(n5796), .D(n5122), .Y(n8337) );
  AOI22X1 U7594 ( .A(n8035), .B(n4915), .C(n7885), .D(n5254), .Y(n8335) );
  NOR3X1 U7595 ( .A(n3967), .B(n4252), .C(n4447), .Y(n8339) );
  NAND3X1 U7596 ( .A(n2735), .B(n3262), .C(n8339), .Y(n8342) );
  AOI22X1 U7597 ( .A(n2958), .B(n6141), .C(n1865), .D(n5783), .Y(n8347) );
  AOI22X1 U7598 ( .A(n1640), .B(n6147), .C(n6288), .D(n6112), .Y(n8346) );
  AOI22X1 U7599 ( .A(n2868), .B(n5780), .C(n2547), .D(n6115), .Y(n8344) );
  NAND3X1 U7600 ( .A(n2469), .B(n3022), .C(n8345), .Y(n8348) );
  AOI22X1 U7601 ( .A(n3832), .B(n6108), .C(n3511), .D(n6106), .Y(n8354) );
  AOI22X1 U7602 ( .A(n1384), .B(n5772), .C(n870), .D(n6145), .Y(n8351) );
  NAND3X1 U7603 ( .A(n2470), .B(n3263), .C(n8352), .Y(n8412) );
  AOI22X1 U7604 ( .A(n6303), .B(n5248), .C(n5978), .D(n5251), .Y(n8360) );
  OAI21X1 U7605 ( .A(n9500), .B(n8355), .C(n5975), .Y(n8359) );
  OAI21X1 U7606 ( .A(n5983), .B(n6091), .C(n6089), .Y(n8357) );
  AOI22X1 U7607 ( .A(n6211), .B(n8357), .C(n5791), .D(n8356), .Y(n8358) );
  NAND3X1 U7608 ( .A(n2471), .B(n8359), .C(n3436), .Y(n8367) );
  NAND3X1 U7609 ( .A(n8102), .B(n5973), .C(n5748), .Y(n8365) );
  AOI22X1 U7610 ( .A(n8362), .B(n8363), .C(n6305), .D(n5229), .Y(n8364) );
  NAND3X1 U7611 ( .A(n4719), .B(n3054), .C(n3437), .Y(n8366) );
  AOI22X1 U7612 ( .A(n7351), .B(n5712), .C(n8035), .D(n4987), .Y(n8373) );
  AOI22X1 U7613 ( .A(n10500), .B(n8370), .C(n3543), .D(n6092), .Y(n8371) );
  NAND3X1 U7614 ( .A(n2472), .B(n3264), .C(n3438), .Y(n8384) );
  AOI22X1 U7615 ( .A(n5799), .B(n8376), .C(n8375), .D(n8374), .Y(n8382) );
  AOI22X1 U7616 ( .A(n5822), .B(n8379), .C(n7147), .D(n8378), .Y(n8380) );
  NAND3X1 U7617 ( .A(n2473), .B(n3265), .C(n3439), .Y(n8383) );
  MUX2X1 U7618 ( .B(n6090), .A(n6067), .S(n6211), .Y(n8385) );
  NAND3X1 U7619 ( .A(n8435), .B(n8385), .C(n8433), .Y(n8386) );
  MUX2X1 U7620 ( .B(n5832), .A(n2794), .S(n5985), .Y(n8389) );
  AOI22X1 U7621 ( .A(n790), .B(n5825), .C(n5966), .D(n9969), .Y(n8387) );
  NAND3X1 U7622 ( .A(n8389), .B(n3267), .C(n3440), .Y(n8394) );
  AOI22X1 U7623 ( .A(n718), .B(n6119), .C(n2259), .D(n6104), .Y(n8392) );
  AOI22X1 U7624 ( .A(n2901), .B(n6086), .C(n469), .D(n5839), .Y(n8390) );
  NAND3X1 U7625 ( .A(n2474), .B(n3268), .C(n3441), .Y(n8393) );
  AOI22X1 U7626 ( .A(n1561), .B(n5779), .C(n902), .D(n5824), .Y(n8397) );
  AOI22X1 U7627 ( .A(n397), .B(n5778), .C(n581), .D(n6135), .Y(n8395) );
  AOI22X1 U7628 ( .A(n3864), .B(n5828), .C(n3222), .D(n5827), .Y(n8400) );
  AOI22X1 U7629 ( .A(n1047), .B(n5786), .C(n1304), .D(n5785), .Y(n8398) );
  NOR3X1 U7630 ( .A(n8401), .B(n4175), .C(n4451), .Y(n8402) );
  NAND3X1 U7631 ( .A(n2736), .B(n3266), .C(n8402), .Y(n8405) );
  AOI22X1 U7632 ( .A(n137), .B(n6141), .C(n1866), .D(n5783), .Y(n8410) );
  AOI22X1 U7633 ( .A(n1641), .B(n5784), .C(n5945), .D(n6112), .Y(n8409) );
  AOI22X1 U7634 ( .A(n2869), .B(n6110), .C(n2548), .D(n6115), .Y(n8407) );
  NAND3X1 U7635 ( .A(n8408), .B(n3024), .C(n126), .Y(n8411) );
  OR2X2 U7636 ( .A(n103), .B(n112), .Y(result[34]) );
  AOI22X1 U7637 ( .A(n871), .B(n5771), .C(n550), .D(n5773), .Y(n8470) );
  AOI22X1 U7638 ( .A(n8374), .B(n5709), .C(n8156), .D(n8413), .Y(n8417) );
  AOI22X1 U7639 ( .A(n8415), .B(n7351), .C(n8035), .D(n4918), .Y(n8416) );
  AOI22X1 U7640 ( .A(n7946), .B(n5799), .C(n5802), .D(n5205), .Y(n8422) );
  AOI22X1 U7641 ( .A(n4900), .B(n5748), .C(n5796), .D(n5056), .Y(n8420) );
  NAND3X1 U7642 ( .A(n2475), .B(n3269), .C(n3442), .Y(n8423) );
  OAI21X1 U7643 ( .A(n6308), .B(n6091), .C(n6089), .Y(n8425) );
  AOI22X1 U7644 ( .A(n5980), .B(n5251), .C(n6213), .D(n8425), .Y(n8428) );
  AOI22X1 U7645 ( .A(n8426), .B(n10505), .C(n5861), .D(n10491), .Y(n8427) );
  NAND3X1 U7646 ( .A(n5806), .B(n10487), .C(n6192), .Y(n8430) );
  AOI22X1 U7647 ( .A(n5983), .B(n5229), .C(n6305), .D(n5248), .Y(n8429) );
  NOR3X1 U7648 ( .A(n8432), .B(n4253), .C(n4455), .Y(n8456) );
  MUX2X1 U7649 ( .B(n6090), .A(n6067), .S(n6213), .Y(n8434) );
  NAND3X1 U7650 ( .A(n8435), .B(n8434), .C(n8433), .Y(n8436) );
  MUX2X1 U7651 ( .B(n5832), .A(n2795), .S(n6308), .Y(n8439) );
  AOI22X1 U7652 ( .A(n2581), .B(n6102), .C(n2902), .D(n5829), .Y(n8437) );
  NAND3X1 U7653 ( .A(n8439), .B(n3270), .C(n3443), .Y(n8444) );
  AOI22X1 U7654 ( .A(n6098), .B(n6356), .C(n398), .D(n5778), .Y(n8442) );
  AOI22X1 U7655 ( .A(n719), .B(n6119), .C(n2260), .D(n5838), .Y(n8440) );
  NAND3X1 U7656 ( .A(n2476), .B(n3271), .C(n3444), .Y(n8443) );
  AOI22X1 U7657 ( .A(n1787), .B(n5777), .C(n1562), .D(n6123), .Y(n8446) );
  AOI22X1 U7658 ( .A(n903), .B(n5824), .C(n5978), .D(n9500), .Y(n8445) );
  AOI22X1 U7659 ( .A(n7172), .B(n5101), .C(n10500), .D(n4943), .Y(n8450) );
  AOI22X1 U7660 ( .A(n3865), .B(n5828), .C(n3223), .D(n6100), .Y(n8448) );
  NAND3X1 U7661 ( .A(n2477), .B(n5683), .C(n5624), .Y(n8451) );
  NOR3X1 U7662 ( .A(n8453), .B(n4254), .C(n4459), .Y(n8455) );
  AOI22X1 U7663 ( .A(n791), .B(n5825), .C(n1128), .D(n5826), .Y(n8454) );
  NAND3X1 U7664 ( .A(n8456), .B(n8455), .C(n5690), .Y(n8460) );
  AOI22X1 U7665 ( .A(n1048), .B(n5786), .C(n1305), .D(n5785), .Y(n8458) );
  AOI22X1 U7666 ( .A(n1385), .B(n5772), .C(n3833), .D(n5775), .Y(n8465) );
  AOI22X1 U7667 ( .A(n2549), .B(n6115), .C(n2870), .D(n6110), .Y(n8464) );
  AOI22X1 U7668 ( .A(n6290), .B(n6112), .C(n3191), .D(n5776), .Y(n8462) );
  AOI22X1 U7669 ( .A(n3512), .B(n6106), .C(n2228), .D(n6113), .Y(n8461) );
  NAND3X1 U7670 ( .A(n128), .B(n3025), .C(n8463), .Y(n8466) );
  AOI22X1 U7671 ( .A(n1642), .B(n6147), .C(n5783), .D(n1867), .Y(n8468) );
  NAND3X1 U7672 ( .A(n127), .B(n142), .C(n8469), .Y(n10615) );
  AOI22X1 U7673 ( .A(n1643), .B(n5784), .C(n5783), .D(n1868), .Y(n8520) );
  AOI22X1 U7674 ( .A(n2229), .B(n6113), .C(n2550), .D(n6115), .Y(n8475) );
  AOI22X1 U7675 ( .A(n2871), .B(n6110), .C(n3192), .D(n5776), .Y(n8474) );
  OAI21X1 U7676 ( .A(n5722), .B(n6292), .C(n5406), .Y(n8472) );
  AOI21X1 U7677 ( .A(n3513), .B(n6106), .C(n8472), .Y(n8473) );
  NAND3X1 U7678 ( .A(n2479), .B(n3026), .C(n3642), .Y(n8476) );
  AOI22X1 U7679 ( .A(n471), .B(n5839), .C(n792), .D(n5825), .Y(n8514) );
  AOI22X1 U7680 ( .A(n5748), .B(n4921), .C(n5796), .D(n5083), .Y(n8481) );
  AOI22X1 U7681 ( .A(n8035), .B(n4889), .C(n7172), .D(n5152), .Y(n8480) );
  AOI22X1 U7682 ( .A(n3545), .B(n5830), .C(n3866), .D(n6096), .Y(n8478) );
  AOI22X1 U7683 ( .A(n4901), .B(n10574), .C(n5802), .D(n5245), .Y(n8484) );
  OAI21X1 U7684 ( .A(n8482), .B(n5644), .C(n1875), .Y(n8490) );
  AOI22X1 U7685 ( .A(n6308), .B(n5229), .C(n5984), .D(n5248), .Y(n8488) );
  OAI21X1 U7686 ( .A(n5989), .B(n6091), .C(n6089), .Y(n8486) );
  AOI22X1 U7687 ( .A(n6305), .B(n5251), .C(n6215), .D(n8486), .Y(n8487) );
  NOR3X1 U7688 ( .A(n3972), .B(n8490), .C(n4601), .Y(n8510) );
  AOI22X1 U7689 ( .A(n1788), .B(n5777), .C(n1563), .D(n5779), .Y(n8495) );
  AOI22X1 U7690 ( .A(n904), .B(n5824), .C(n6303), .D(n9500), .Y(n8494) );
  OAI21X1 U7691 ( .A(n6099), .B(n6359), .C(n5407), .Y(n8492) );
  AOI21X1 U7692 ( .A(n583), .B(n5823), .C(n8492), .Y(n8493) );
  AOI22X1 U7693 ( .A(n2903), .B(n6086), .C(n5970), .D(n9969), .Y(n8503) );
  AOI21X1 U7694 ( .A(n8238), .B(n5799), .C(n8496), .Y(n8500) );
  MUX2X1 U7695 ( .B(n6090), .A(n6067), .S(n6215), .Y(n8499) );
  NOR3X1 U7696 ( .A(n5265), .B(n5263), .C(n4856), .Y(n8498) );
  NAND3X1 U7697 ( .A(n2704), .B(n8499), .C(n8498), .Y(n8501) );
  MUX2X1 U7698 ( .B(n5832), .A(n2796), .S(n5988), .Y(n8502) );
  AOI22X1 U7699 ( .A(n720), .B(n6119), .C(n2261), .D(n6104), .Y(n8505) );
  NOR3X1 U7700 ( .A(n3977), .B(n4255), .C(n4602), .Y(n8509) );
  NAND3X1 U7701 ( .A(n8510), .B(n3665), .C(n8509), .Y(n8511) );
  AOI21X1 U7702 ( .A(n1306), .B(n6125), .C(n121), .Y(n8512) );
  NAND3X1 U7703 ( .A(n2480), .B(n3272), .C(n3643), .Y(n8515) );
  AOI22X1 U7704 ( .A(n5773), .B(n551), .C(n872), .D(n6145), .Y(n8518) );
  NAND3X1 U7705 ( .A(n2478), .B(n8519), .C(n143), .Y(n10614) );
  AOI22X1 U7706 ( .A(n3771), .B(n6108), .C(n3450), .D(n6106), .Y(n8525) );
  AOI22X1 U7707 ( .A(n1323), .B(n5772), .C(n809), .D(n5771), .Y(n8522) );
  NAND3X1 U7708 ( .A(n2481), .B(n5305), .C(n8523), .Y(n8579) );
  NAND3X1 U7709 ( .A(n4736), .B(n4781), .C(n4832), .Y(n8527) );
  NAND3X1 U7710 ( .A(n4871), .B(n8526), .C(n4970), .Y(n8812) );
  MUX2X1 U7711 ( .B(n2768), .A(n4964), .S(n5907), .Y(n8528) );
  AOI22X1 U7712 ( .A(n5768), .B(n6337), .C(n8588), .D(n5271), .Y(n8530) );
  AOI22X1 U7713 ( .A(n8610), .B(n6018), .C(n8554), .D(n6016), .Y(n8529) );
  AOI22X1 U7714 ( .A(n5768), .B(n6008), .C(n8588), .D(n5285), .Y(n8531) );
  AOI22X1 U7715 ( .A(n8762), .B(n5236), .C(n8999), .D(n5086), .Y(n8532) );
  OAI21X1 U7716 ( .A(n5883), .B(n8528), .C(n1876), .Y(n8535) );
  AOI22X1 U7717 ( .A(n10), .B(n6077), .C(n6332), .D(n6081), .Y(n8533) );
  AOI22X1 U7718 ( .A(n8535), .B(n9647), .C(n9774), .D(n5146), .Y(n8540) );
  AOI22X1 U7719 ( .A(n3546), .B(n5830), .C(n3867), .D(n6096), .Y(n8539) );
  AOI22X1 U7720 ( .A(n3225), .B(n5827), .C(n1757), .D(n5777), .Y(n8537) );
  AOI22X1 U7721 ( .A(n1018), .B(n5786), .C(n1275), .D(n5785), .Y(n8536) );
  AOI22X1 U7722 ( .A(n4955), .B(n10087), .C(n8542), .D(n5733), .Y(n8547) );
  OAI21X1 U7723 ( .A(n5908), .B(n10104), .C(n5174), .Y(n8545) );
  AOI22X1 U7724 ( .A(n6018), .B(n6077), .C(n5282), .D(n6081), .Y(n8544) );
  AOI22X1 U7725 ( .A(n6079), .B(n5272), .C(n5286), .D(n6083), .Y(n8543) );
  AOI22X1 U7726 ( .A(n5740), .B(n8545), .C(n5742), .D(n5216), .Y(n8546) );
  AOI22X1 U7727 ( .A(n5276), .B(n9793), .C(n6315), .D(n6065), .Y(n8550) );
  OAI21X1 U7728 ( .A(n5880), .B(n6091), .C(n6089), .Y(n8548) );
  AOI22X1 U7729 ( .A(n5993), .B(n6066), .C(n5267), .D(n8548), .Y(n8549) );
  NOR3X1 U7730 ( .A(n3982), .B(n4256), .C(n4603), .Y(n8571) );
  AOI22X1 U7731 ( .A(n2583), .B(n6102), .C(n2904), .D(n5829), .Y(n8563) );
  AOI22X1 U7732 ( .A(n440), .B(n6131), .C(n761), .D(n5825), .Y(n8562) );
  AOI22X1 U7733 ( .A(n6004), .B(n6094), .C(n1066), .D(n5826), .Y(n8560) );
  NAND3X1 U7734 ( .A(n4737), .B(n5724), .C(n6085), .Y(n8553) );
  MUX2X1 U7735 ( .B(n6091), .A(n6068), .S(n5267), .Y(n8556) );
  OAI21X1 U7736 ( .A(n151), .B(n5010), .C(n6070), .Y(n8555) );
  NAND3X1 U7737 ( .A(n9441), .B(n5736), .C(n3666), .Y(n8558) );
  MUX2X1 U7738 ( .B(n5832), .A(n2797), .S(n5991), .Y(n8559) );
  AOI22X1 U7739 ( .A(n384), .B(n5778), .C(n584), .D(n5823), .Y(n8565) );
  AOI22X1 U7740 ( .A(n705), .B(n5790), .C(n2262), .D(n5838), .Y(n8564) );
  AOI22X1 U7741 ( .A(n1532), .B(n5779), .C(n905), .D(n6133), .Y(n8567) );
  AOI22X1 U7742 ( .A(n27), .B(n9500), .C(n5912), .D(n10502), .Y(n8566) );
  NOR3X1 U7743 ( .A(n3987), .B(n4257), .C(n4604), .Y(n8570) );
  AOI22X1 U7744 ( .A(n2985), .B(n6141), .C(n1805), .D(n5783), .Y(n8577) );
  AOI22X1 U7745 ( .A(n1580), .B(n6147), .C(n59), .D(n6112), .Y(n8576) );
  AOI22X1 U7746 ( .A(n2808), .B(n6110), .C(n2487), .D(n6115), .Y(n8574) );
  NAND3X1 U7747 ( .A(n2482), .B(n3027), .C(n8575), .Y(n8578) );
  AOI22X1 U7748 ( .A(n3451), .B(n6106), .C(n3130), .D(n5776), .Y(n8582) );
  AOI22X1 U7749 ( .A(n810), .B(n5771), .C(n489), .D(n5773), .Y(n8580) );
  NAND3X1 U7750 ( .A(n2483), .B(n3273), .C(n3445), .Y(n8651) );
  AOI22X1 U7751 ( .A(n2488), .B(n5781), .C(n2167), .D(n6113), .Y(n8649) );
  MUX2X1 U7752 ( .B(n5992), .A(n5879), .S(n5267), .Y(n8583) );
  AOI21X1 U7753 ( .A(n8554), .B(n5993), .C(n8754), .Y(n8584) );
  NAND3X1 U7754 ( .A(n4738), .B(n4782), .C(n3644), .Y(n8585) );
  AOI22X1 U7755 ( .A(n9109), .B(n4944), .C(n3364), .D(n5256), .Y(n8591) );
  AOI21X1 U7756 ( .A(n8554), .B(n72), .C(n2371), .Y(n8609) );
  NAND3X1 U7757 ( .A(n4840), .B(n4780), .C(n3667), .Y(n8618) );
  AOI22X1 U7758 ( .A(n5768), .B(n5269), .C(n8588), .D(n5286), .Y(n8589) );
  AOI22X1 U7759 ( .A(n5737), .B(n8881), .C(n5752), .D(n5165), .Y(n8590) );
  AOI22X1 U7760 ( .A(n43), .B(n9793), .C(n5276), .D(n6065), .Y(n8596) );
  OAI21X1 U7761 ( .A(n5993), .B(n6091), .C(n6089), .Y(n8593) );
  OAI21X1 U7762 ( .A(n6064), .B(n6313), .C(n5346), .Y(n8871) );
  AOI22X1 U7763 ( .A(n6217), .B(n8593), .C(n5837), .D(n9916), .Y(n8594) );
  NAND3X1 U7764 ( .A(n2485), .B(n3274), .C(n3446), .Y(n8597) );
  AOI21X1 U7765 ( .A(n6337), .B(n9632), .C(n5396), .Y(n8600) );
  OAI21X1 U7766 ( .A(n6340), .B(n6082), .C(n5395), .Y(n9389) );
  OAI21X1 U7767 ( .A(n6340), .B(n6153), .C(n5395), .Y(n9388) );
  OAI21X1 U7768 ( .A(n8602), .B(n5731), .C(n1930), .Y(n9379) );
  AOI21X1 U7769 ( .A(n6083), .B(n72), .C(n2372), .Y(n8606) );
  OAI21X1 U7770 ( .A(n6322), .B(n6078), .C(n4841), .Y(n8604) );
  AOI22X1 U7771 ( .A(n6731), .B(n9379), .C(n8882), .D(n10375), .Y(n8608) );
  NAND3X1 U7772 ( .A(n4841), .B(n6062), .C(n3668), .Y(n8615) );
  AOI22X1 U7773 ( .A(n8968), .B(n4945), .C(n3547), .D(n6092), .Y(n8607) );
  OAI21X1 U7774 ( .A(n6322), .B(n4802), .C(n4840), .Y(n8611) );
  AOI22X1 U7775 ( .A(n8610), .B(n6337), .C(n8554), .D(n6018), .Y(n8614) );
  AOI22X1 U7776 ( .A(n5768), .B(n10487), .C(n6217), .D(n7491), .Y(n8612) );
  OAI21X1 U7777 ( .A(n5766), .B(n3355), .C(n8613), .Y(n9386) );
  AOI22X1 U7778 ( .A(n8755), .B(n8880), .C(n8762), .D(n9386), .Y(n8621) );
  AOI21X1 U7779 ( .A(n5286), .B(n5800), .C(n9142), .Y(n8616) );
  AOI22X1 U7780 ( .A(n9774), .B(n5074), .C(n8738), .D(n4868), .Y(n8619) );
  NAND3X1 U7781 ( .A(n2486), .B(n3275), .C(n3447), .Y(n8622) );
  MUX2X1 U7782 ( .B(n6090), .A(n6067), .S(n6217), .Y(n8624) );
  NAND3X1 U7783 ( .A(n8624), .B(n6069), .C(n9803), .Y(n8625) );
  MUX2X1 U7784 ( .B(n5832), .A(n5603), .S(n5992), .Y(n8628) );
  AOI22X1 U7785 ( .A(n762), .B(n5825), .C(n10), .D(n9969), .Y(n8626) );
  NAND3X1 U7786 ( .A(n8628), .B(n3277), .C(n3448), .Y(n8633) );
  AOI22X1 U7787 ( .A(n706), .B(n6119), .C(n2263), .D(n6104), .Y(n8631) );
  AOI22X1 U7788 ( .A(n2905), .B(n6086), .C(n441), .D(n5839), .Y(n8629) );
  NAND3X1 U7789 ( .A(n2615), .B(n3278), .C(n3449), .Y(n8632) );
  AOI22X1 U7790 ( .A(n6319), .B(n9500), .C(n5915), .D(n10502), .Y(n8635) );
  AOI22X1 U7791 ( .A(n385), .B(n6117), .C(n585), .D(n6135), .Y(n8634) );
  AOI22X1 U7792 ( .A(n3868), .B(n5828), .C(n3226), .D(n6100), .Y(n8638) );
  AOI22X1 U7793 ( .A(n1276), .B(n5785), .C(n906), .D(n6133), .Y(n8636) );
  NOR3X1 U7794 ( .A(n8640), .B(n4258), .C(n4460), .Y(n8641) );
  NAND3X1 U7795 ( .A(n2737), .B(n3276), .C(n8641), .Y(n8644) );
  OAI21X1 U7796 ( .A(n5722), .B(n6341), .C(n1931), .Y(n8646) );
  AOI21X1 U7797 ( .A(n2809), .B(n6110), .C(n8646), .Y(n8647) );
  NAND3X1 U7798 ( .A(n2484), .B(n5681), .C(n3645), .Y(n8650) );
  AOI22X1 U7799 ( .A(n2906), .B(n6086), .C(n490), .D(n5849), .Y(n8656) );
  OAI21X1 U7800 ( .A(n5583), .B(n6343), .C(n5431), .Y(n8653) );
  AOI21X1 U7801 ( .A(n1582), .B(n5846), .C(n8653), .Y(n8654) );
  AOI22X1 U7802 ( .A(n707), .B(n6119), .C(n2264), .D(n6104), .Y(n8658) );
  AOI22X1 U7803 ( .A(n5283), .B(n9500), .C(n5918), .D(n10502), .Y(n8660) );
  AOI22X1 U7804 ( .A(n386), .B(n6117), .C(n586), .D(n6135), .Y(n8659) );
  NOR3X1 U7805 ( .A(n3992), .B(n4259), .C(n4605), .Y(n8729) );
  AOI22X1 U7806 ( .A(n2810), .B(n5835), .C(n442), .D(n5839), .Y(n8669) );
  AOI22X1 U7807 ( .A(n6008), .B(n6094), .C(n1068), .D(n5826), .Y(n8666) );
  MUX2X1 U7808 ( .B(n6090), .A(n6067), .S(n5907), .Y(n8663) );
  NAND3X1 U7809 ( .A(n8663), .B(n6069), .C(n9803), .Y(n8664) );
  MUX2X1 U7810 ( .B(n5832), .A(n2798), .S(n5995), .Y(n8665) );
  NAND3X1 U7811 ( .A(n5414), .B(n5544), .C(n8667), .Y(n8676) );
  AOI22X1 U7812 ( .A(n3773), .B(n5845), .C(n2168), .D(n5843), .Y(n8671) );
  AOI22X1 U7813 ( .A(n1807), .B(n5842), .C(n3131), .D(n5844), .Y(n8673) );
  NOR3X1 U7814 ( .A(n3996), .B(n4260), .C(n4606), .Y(n8728) );
  OAI21X1 U7815 ( .A(n5907), .B(n9846), .C(n5394), .Y(n8996) );
  OAI21X1 U7816 ( .A(n5995), .B(n6091), .C(n6089), .Y(n8681) );
  AOI22X1 U7817 ( .A(n5993), .B(n6077), .C(n5991), .D(n6081), .Y(n8680) );
  OAI21X1 U7818 ( .A(n6064), .B(n6316), .C(n1877), .Y(n9458) );
  AOI22X1 U7819 ( .A(n5907), .B(n8681), .C(n9458), .D(n6072), .Y(n8682) );
  OAI21X1 U7820 ( .A(n167), .B(n8683), .C(n1878), .Y(n8690) );
  AOI22X1 U7821 ( .A(n5768), .B(n5286), .C(n8588), .D(n6018), .Y(n8684) );
  NAND3X1 U7822 ( .A(n8999), .B(n7491), .C(n5194), .Y(n8687) );
  AOI22X1 U7823 ( .A(n27), .B(n6065), .C(n5276), .D(n6066), .Y(n8686) );
  NAND3X1 U7824 ( .A(n2738), .B(n3055), .C(n3578), .Y(n8689) );
  MUX2X1 U7825 ( .B(n6340), .A(n6338), .S(n8554), .Y(n8691) );
  MUX2X1 U7826 ( .B(n6338), .A(n6340), .S(n5267), .Y(n8692) );
  MUX2X1 U7827 ( .B(n172), .A(n5642), .S(n5908), .Y(n8693) );
  OAI21X1 U7828 ( .A(n6219), .B(n5570), .C(n1932), .Y(n9179) );
  AOI22X1 U7829 ( .A(n5269), .B(n6077), .C(n5286), .D(n9626), .Y(n8696) );
  AOI22X1 U7830 ( .A(n6018), .B(n6079), .C(n6008), .D(n6083), .Y(n8695) );
  MUX2X1 U7831 ( .B(n6337), .A(n5272), .S(n5887), .Y(n8697) );
  MUX2X1 U7832 ( .B(n5579), .A(n5509), .S(n5890), .Y(n8698) );
  AOI22X1 U7833 ( .A(n8954), .B(n5579), .C(n9183), .D(n5770), .Y(n8699) );
  OAI21X1 U7834 ( .A(n8700), .B(n6221), .C(n1879), .Y(n8707) );
  MUX2X1 U7835 ( .B(n5274), .A(n6322), .S(n8554), .Y(n8947) );
  NAND3X1 U7836 ( .A(n4740), .B(n4783), .C(n3669), .Y(n8704) );
  MUX2X1 U7837 ( .B(n6324), .A(n6326), .S(n5267), .Y(n8703) );
  AOI22X1 U7838 ( .A(n2959), .B(n5256), .C(n5737), .D(n8717), .Y(n8705) );
  OAI21X1 U7839 ( .A(n8947), .B(n5711), .C(n1880), .Y(n8706) );
  AOI22X1 U7840 ( .A(n3227), .B(n6100), .C(n1759), .D(n5777), .Y(n8714) );
  AOI22X1 U7841 ( .A(n1277), .B(n5785), .C(n1534), .D(n5779), .Y(n8711) );
  MUX2X1 U7842 ( .B(n6322), .A(n6003), .S(n5888), .Y(n8715) );
  AOI22X1 U7843 ( .A(n5717), .B(n6721), .C(n8738), .D(n4990), .Y(n8725) );
  MUX2X1 U7844 ( .B(n6024), .A(n6337), .S(n9688), .Y(n9185) );
  MUX2X1 U7845 ( .B(n6003), .A(n5283), .S(n9688), .Y(n8718) );
  AOI22X1 U7846 ( .A(n6730), .B(n9461), .C(n10375), .D(n8964), .Y(n8724) );
  AOI21X1 U7847 ( .A(n6328), .B(n9626), .C(n5717), .Y(n8719) );
  OAI21X1 U7848 ( .A(n6062), .B(n6331), .C(n1906), .Y(n8966) );
  OAI21X1 U7849 ( .A(n8721), .B(n5520), .C(n1933), .Y(n8722) );
  AOI21X1 U7850 ( .A(n3869), .B(n6096), .C(n8722), .Y(n8723) );
  NOR3X1 U7851 ( .A(n4123), .B(n4179), .C(n4464), .Y(n8727) );
  NAND3X1 U7852 ( .A(n8729), .B(n8728), .C(n8727), .Y(n8730) );
  AOI22X1 U7853 ( .A(n3774), .B(n6108), .C(n3453), .D(n6106), .Y(n8735) );
  AOI22X1 U7854 ( .A(n1326), .B(n5772), .C(n812), .D(n5771), .Y(n8732) );
  NAND3X1 U7855 ( .A(n2616), .B(n5312), .C(n8733), .Y(n8793) );
  AOI21X1 U7856 ( .A(n6008), .B(n5800), .C(n8990), .Y(n8736) );
  AOI22X1 U7857 ( .A(n8968), .B(n4892), .C(n3549), .D(n6092), .Y(n8750) );
  AOI22X1 U7858 ( .A(n3870), .B(n6096), .C(n3228), .D(n5827), .Y(n8749) );
  AOI21X1 U7859 ( .A(n8588), .B(n6332), .C(n9138), .Y(n8737) );
  NAND3X1 U7860 ( .A(n5883), .B(n5271), .C(n7491), .Y(n9326) );
  OAI21X1 U7861 ( .A(n8739), .B(n5506), .C(n4698), .Y(n8747) );
  AOI22X1 U7862 ( .A(n5286), .B(n6077), .C(n6018), .D(n6081), .Y(n8740) );
  AOI22X1 U7863 ( .A(n5768), .B(n6018), .C(n8588), .D(n6022), .Y(n8743) );
  AOI22X1 U7864 ( .A(n5737), .B(n8742), .C(n5752), .D(n5089), .Y(n8745) );
  OAI21X1 U7865 ( .A(n160), .B(n5655), .C(n1881), .Y(n8746) );
  AOI22X1 U7866 ( .A(n6315), .B(n6077), .C(n5992), .D(n6081), .Y(n8752) );
  AOI22X1 U7867 ( .A(n5991), .B(n6079), .C(n5276), .D(n6083), .Y(n8751) );
  AOI22X1 U7868 ( .A(n5768), .B(n5993), .C(n8588), .D(n5880), .Y(n8753) );
  AOI22X1 U7869 ( .A(n5238), .B(n5628), .C(n8996), .D(n5200), .Y(n8761) );
  NAND3X1 U7870 ( .A(n4741), .B(n4784), .C(n3670), .Y(n8758) );
  AOI22X1 U7871 ( .A(n5274), .B(n2779), .C(n3365), .D(n5256), .Y(n8760) );
  OAI21X1 U7872 ( .A(n4756), .B(n5031), .C(n9791), .Y(n8763) );
  AOI22X1 U7873 ( .A(n5271), .B(n8763), .C(n6322), .D(n9793), .Y(n8767) );
  OAI21X1 U7874 ( .A(n5276), .B(n6091), .C(n6089), .Y(n8764) );
  AOI22X1 U7875 ( .A(n43), .B(n6066), .C(n6220), .D(n8764), .Y(n8765) );
  NOR3X1 U7876 ( .A(n3997), .B(n4261), .C(n4469), .Y(n8785) );
  AOI22X1 U7877 ( .A(n2265), .B(n5838), .C(n2586), .D(n6102), .Y(n8776) );
  AOI22X1 U7878 ( .A(n2907), .B(n6086), .C(n443), .D(n5839), .Y(n8775) );
  AOI22X1 U7879 ( .A(n764), .B(n5825), .C(n5285), .D(n9969), .Y(n8773) );
  MUX2X1 U7880 ( .B(n6091), .A(n6068), .S(n5883), .Y(n8769) );
  NOR3X1 U7881 ( .A(n5728), .B(n9731), .C(n8769), .Y(n8770) );
  MUX2X1 U7882 ( .B(n10522), .A(n8770), .S(n5276), .Y(n8771) );
  AOI21X1 U7883 ( .A(n1069), .B(n6127), .C(n8771), .Y(n8772) );
  NAND3X1 U7884 ( .A(n5350), .B(n5547), .C(n8774), .Y(n8783) );
  AOI22X1 U7885 ( .A(n5922), .B(n10502), .C(n387), .D(n5778), .Y(n8778) );
  AOI22X1 U7886 ( .A(n587), .B(n5823), .C(n708), .D(n6119), .Y(n8777) );
  AOI22X1 U7887 ( .A(n1760), .B(n5777), .C(n1021), .D(n6129), .Y(n8781) );
  AOI22X1 U7888 ( .A(n1535), .B(n5779), .C(n908), .D(n5824), .Y(n8779) );
  NOR3X1 U7889 ( .A(n4001), .B(n4262), .C(n4473), .Y(n8784) );
  AOI22X1 U7890 ( .A(n2986), .B(n6141), .C(n1808), .D(n5783), .Y(n8791) );
  AOI22X1 U7891 ( .A(n1583), .B(n6147), .C(n6032), .D(n6112), .Y(n8790) );
  AOI22X1 U7892 ( .A(n2811), .B(n6110), .C(n2490), .D(n6115), .Y(n8788) );
  NAND3X1 U7893 ( .A(n2617), .B(n3028), .C(n8789), .Y(n8792) );
  AOI22X1 U7894 ( .A(n3775), .B(n6108), .C(n3454), .D(n6106), .Y(n8798) );
  AOI22X1 U7895 ( .A(n1327), .B(n5772), .C(n813), .D(n6145), .Y(n8795) );
  NAND3X1 U7896 ( .A(n2618), .B(n5320), .C(n8796), .Y(n8845) );
  AOI22X1 U7897 ( .A(n5752), .B(n5236), .C(n9774), .D(n5216), .Y(n8803) );
  AOI22X1 U7898 ( .A(n8738), .B(n5086), .C(n8968), .D(n5146), .Y(n8802) );
  AOI22X1 U7899 ( .A(n3550), .B(n5830), .C(n3871), .D(n6096), .Y(n8800) );
  AOI22X1 U7900 ( .A(n3229), .B(n5827), .C(n1761), .D(n6121), .Y(n8799) );
  AOI22X1 U7901 ( .A(n5276), .B(n6077), .C(n5995), .D(n6081), .Y(n8804) );
  AOI21X1 U7902 ( .A(n8588), .B(n5992), .C(n8807), .Y(n8808) );
  AOI22X1 U7903 ( .A(n5098), .B(n5628), .C(n8996), .D(n5168), .Y(n8814) );
  OAI21X1 U7904 ( .A(n9846), .B(n6219), .C(n5441), .Y(n8992) );
  AOI22X1 U7905 ( .A(n5740), .B(n8992), .C(n5256), .D(n4964), .Y(n8813) );
  OAI21X1 U7906 ( .A(n10375), .B(n8755), .C(n6325), .Y(n8815) );
  OAI21X1 U7907 ( .A(n27), .B(n6091), .C(n6089), .Y(n8818) );
  AOI22X1 U7908 ( .A(n6222), .B(n8818), .C(n4955), .D(n6073), .Y(n8819) );
  NOR3X1 U7909 ( .A(n4002), .B(n4263), .C(n4477), .Y(n8837) );
  AOI22X1 U7910 ( .A(n1022), .B(n5786), .C(n1279), .D(n5785), .Y(n8826) );
  AOI22X1 U7911 ( .A(n1536), .B(n5779), .C(n909), .D(n5824), .Y(n8825) );
  AOI22X1 U7912 ( .A(n66), .B(n10502), .C(n388), .D(n6117), .Y(n8823) );
  AOI22X1 U7913 ( .A(n588), .B(n6135), .C(n709), .D(n5790), .Y(n8822) );
  NAND3X1 U7914 ( .A(n2619), .B(n5499), .C(n8824), .Y(n8835) );
  MUX2X1 U7915 ( .B(n6090), .A(n6067), .S(n6222), .Y(n8827) );
  MUX2X1 U7916 ( .B(n6088), .A(n5295), .S(n27), .Y(n8831) );
  AOI22X1 U7917 ( .A(n765), .B(n5825), .C(n6016), .D(n9969), .Y(n8829) );
  AOI22X1 U7918 ( .A(n2266), .B(n6104), .C(n2587), .D(n6102), .Y(n8833) );
  AOI22X1 U7919 ( .A(n2908), .B(n6086), .C(n444), .D(n5839), .Y(n8832) );
  NOR3X1 U7920 ( .A(n4007), .B(n4183), .C(n4607), .Y(n8836) );
  AOI22X1 U7921 ( .A(n2987), .B(n6141), .C(n1809), .D(n5783), .Y(n8843) );
  AOI22X1 U7922 ( .A(n1584), .B(n6147), .C(n5885), .D(n6112), .Y(n8842) );
  AOI22X1 U7923 ( .A(n2812), .B(n6110), .C(n2491), .D(n5781), .Y(n8840) );
  NAND3X1 U7924 ( .A(n2620), .B(n3029), .C(n8841), .Y(n8844) );
  AOI22X1 U7925 ( .A(n3776), .B(n6108), .C(n3455), .D(n6106), .Y(n8850) );
  AOI22X1 U7926 ( .A(n1328), .B(n5772), .C(n814), .D(n5771), .Y(n8847) );
  NAND3X1 U7927 ( .A(n2621), .B(n5328), .C(n8848), .Y(n8908) );
  AOI22X1 U7928 ( .A(n5992), .B(n9500), .C(n5924), .D(n10502), .Y(n8852) );
  AOI22X1 U7929 ( .A(n389), .B(n6117), .C(n589), .D(n6135), .Y(n8851) );
  AOI22X1 U7930 ( .A(n1762), .B(n5777), .C(n1023), .D(n6129), .Y(n8855) );
  AOI22X1 U7931 ( .A(n1537), .B(n5779), .C(n910), .D(n6133), .Y(n8853) );
  NAND3X1 U7932 ( .A(n2622), .B(n5678), .C(n3579), .Y(n8856) );
  MUX2X1 U7933 ( .B(n6090), .A(n6067), .S(n6224), .Y(n8858) );
  MUX2X1 U7934 ( .B(n6088), .A(n5318), .S(n6319), .Y(n8862) );
  AOI22X1 U7935 ( .A(n766), .B(n5825), .C(n6018), .D(n9969), .Y(n8860) );
  NAND3X1 U7936 ( .A(n8862), .B(n3279), .C(n3580), .Y(n8867) );
  AOI22X1 U7937 ( .A(n710), .B(n6119), .C(n2267), .D(n5838), .Y(n8865) );
  AOI22X1 U7938 ( .A(n2909), .B(n6086), .C(n445), .D(n5839), .Y(n8863) );
  NAND3X1 U7939 ( .A(n2623), .B(n3280), .C(n5688), .Y(n8866) );
  OAI21X1 U7940 ( .A(n6000), .B(n6091), .C(n6089), .Y(n8868) );
  AOI21X1 U7941 ( .A(n6224), .B(n8868), .C(n5039), .Y(n8888) );
  AOI22X1 U7942 ( .A(n43), .B(n6077), .C(n5276), .D(n9626), .Y(n8870) );
  AOI22X1 U7943 ( .A(n5995), .B(n6079), .C(n6319), .D(n9688), .Y(n8869) );
  MUX2X1 U7944 ( .B(n9139), .A(n8872), .S(n5889), .Y(n9366) );
  AOI21X1 U7945 ( .A(n8554), .B(n6000), .C(n5809), .Y(n8873) );
  MUX2X1 U7946 ( .B(n4877), .A(n5639), .S(n5908), .Y(n8877) );
  AOI22X1 U7947 ( .A(n9366), .B(n9916), .C(n9372), .D(n4944), .Y(n8887) );
  AOI22X1 U7948 ( .A(n8881), .B(n8879), .C(n8880), .D(n8946), .Y(n8885) );
  AOI22X1 U7949 ( .A(n8883), .B(n5822), .C(n8882), .D(n7147), .Y(n8884) );
  AOI22X1 U7950 ( .A(n8968), .B(n5074), .C(n3551), .D(n6092), .Y(n8890) );
  AOI22X1 U7951 ( .A(n3872), .B(n6096), .C(n3230), .D(n5827), .Y(n8889) );
  AOI22X1 U7952 ( .A(n8999), .B(n9386), .C(n8738), .D(n5165), .Y(n8896) );
  AOI22X1 U7953 ( .A(n5833), .B(n9379), .C(n6791), .D(n4945), .Y(n8894) );
  NOR3X1 U7954 ( .A(n4008), .B(n4264), .C(n4480), .Y(n8898) );
  NAND3X1 U7955 ( .A(n2739), .B(n3281), .C(n8898), .Y(n8901) );
  AOI22X1 U7956 ( .A(n2960), .B(n6141), .C(n1810), .D(n5783), .Y(n8906) );
  AOI22X1 U7957 ( .A(n1585), .B(n5784), .C(n6034), .D(n6112), .Y(n8905) );
  AOI22X1 U7958 ( .A(n2813), .B(n5780), .C(n2492), .D(n5781), .Y(n8903) );
  NAND3X1 U7959 ( .A(n2624), .B(n3030), .C(n8904), .Y(n8907) );
  AOI22X1 U7960 ( .A(n2589), .B(n6102), .C(n2910), .D(n6086), .Y(n8914) );
  OAI21X1 U7961 ( .A(n5583), .B(n6344), .C(n1934), .Y(n8911) );
  AOI21X1 U7962 ( .A(n1329), .B(n5848), .C(n8911), .Y(n8912) );
  AOI22X1 U7963 ( .A(n590), .B(n6135), .C(n711), .D(n5790), .Y(n8916) );
  AOI22X1 U7964 ( .A(n911), .B(n5824), .C(n6315), .D(n9500), .Y(n8918) );
  AOI22X1 U7965 ( .A(n5926), .B(n6098), .C(n390), .D(n6117), .Y(n8917) );
  NOR3X1 U7966 ( .A(n4013), .B(n4265), .C(n4608), .Y(n8977) );
  AOI22X1 U7967 ( .A(n2814), .B(n5835), .C(n446), .D(n5839), .Y(n8927) );
  AOI22X1 U7968 ( .A(n5282), .B(n6094), .C(n1072), .D(n5826), .Y(n8924) );
  MUX2X1 U7969 ( .B(n6090), .A(n6067), .S(n56), .Y(n8921) );
  MUX2X1 U7970 ( .B(n5832), .A(n5479), .S(n6322), .Y(n8923) );
  NAND3X1 U7971 ( .A(n5325), .B(n5607), .C(n8925), .Y(n8934) );
  AOI22X1 U7972 ( .A(n3777), .B(n5845), .C(n2172), .D(n5843), .Y(n8929) );
  AOI22X1 U7973 ( .A(n1586), .B(n5846), .C(n1811), .D(n5842), .Y(n8931) );
  AOI22X1 U7974 ( .A(n3135), .B(n5844), .C(n3456), .D(n5847), .Y(n8930) );
  NOR3X1 U7975 ( .A(n4017), .B(n4266), .C(n4609), .Y(n8976) );
  AOI22X1 U7976 ( .A(n5276), .B(n6079), .C(n5283), .D(n6083), .Y(n8935) );
  AOI22X1 U7977 ( .A(n9458), .B(n10574), .C(n8992), .D(n5178), .Y(n8938) );
  OAI21X1 U7978 ( .A(n6071), .B(n165), .C(n1882), .Y(n8943) );
  AOI21X1 U7979 ( .A(n6090), .B(n6324), .C(n10564), .Y(n8941) );
  NAND3X1 U7980 ( .A(n5883), .B(n10487), .C(n5789), .Y(n8940) );
  OAI21X1 U7981 ( .A(n2761), .B(n71), .C(n1907), .Y(n8942) );
  NOR3X1 U7982 ( .A(n8943), .B(n8942), .C(n5039), .Y(n8958) );
  AOI22X1 U7983 ( .A(n5860), .B(n5770), .C(n8717), .D(n8879), .Y(n8945) );
  OAI21X1 U7984 ( .A(n8947), .B(n5174), .C(n1883), .Y(n8956) );
  AOI21X1 U7985 ( .A(n8554), .B(n6322), .C(n8948), .Y(n8949) );
  AOI22X1 U7986 ( .A(n8996), .B(n5033), .C(n8952), .D(n8999), .Y(n8953) );
  OAI21X1 U7987 ( .A(n9185), .B(n5578), .C(n1884), .Y(n8955) );
  AOI22X1 U7988 ( .A(n3873), .B(n5828), .C(n3231), .D(n5827), .Y(n8963) );
  AOI22X1 U7989 ( .A(n1024), .B(n5786), .C(n1281), .D(n5785), .Y(n8960) );
  NAND3X1 U7990 ( .A(n5601), .B(n5675), .C(n8961), .Y(n8973) );
  AOI22X1 U7991 ( .A(n5717), .B(n5822), .C(n7147), .D(n8964), .Y(n8972) );
  AOI22X1 U7992 ( .A(n8738), .B(n5194), .C(n8891), .D(n4990), .Y(n8971) );
  OAI21X1 U7993 ( .A(n9187), .B(n5520), .C(n1935), .Y(n8969) );
  AOI21X1 U7994 ( .A(n3552), .B(n5830), .C(n8969), .Y(n8970) );
  NOR3X1 U7995 ( .A(n4124), .B(n4187), .C(n4484), .Y(n8975) );
  NAND3X1 U7996 ( .A(n8977), .B(n8976), .C(n8975), .Y(n8978) );
  AOI22X1 U7997 ( .A(n3778), .B(n6108), .C(n3457), .D(n6106), .Y(n8983) );
  AOI22X1 U7998 ( .A(n1330), .B(n5772), .C(n816), .D(n5771), .Y(n8980) );
  NAND3X1 U7999 ( .A(n2625), .B(n5341), .C(n8981), .Y(n9027) );
  AOI22X1 U8000 ( .A(n8738), .B(n5089), .C(n8891), .D(n4815), .Y(n8988) );
  AOI22X1 U8001 ( .A(n6791), .B(n4892), .C(n8968), .D(n5019), .Y(n8987) );
  AOI22X1 U8002 ( .A(n3553), .B(n5830), .C(n3874), .D(n6096), .Y(n8985) );
  AOI22X1 U8003 ( .A(n3232), .B(n5827), .C(n1764), .D(n5777), .Y(n8984) );
  AOI22X1 U8004 ( .A(n6322), .B(n9632), .C(n6000), .D(n9626), .Y(n8989) );
  AOI22X1 U8005 ( .A(n8992), .B(n5200), .C(n5155), .D(n5628), .Y(n8998) );
  AOI21X1 U8006 ( .A(n8610), .B(n6322), .C(n8742), .Y(n8993) );
  AOI22X1 U8007 ( .A(n8996), .B(n5053), .C(n8742), .D(n8879), .Y(n8997) );
  OAI21X1 U8008 ( .A(n4757), .B(n5031), .C(n10033), .Y(n9000) );
  OAI21X1 U8009 ( .A(n6003), .B(n6091), .C(n6089), .Y(n9001) );
  AOI22X1 U8010 ( .A(n6228), .B(n9001), .C(n5238), .D(n10574), .Y(n9002) );
  NOR3X1 U8011 ( .A(n4018), .B(n4267), .C(n4489), .Y(n9019) );
  AOI22X1 U8012 ( .A(n1025), .B(n5786), .C(n1282), .D(n5785), .Y(n9009) );
  AOI22X1 U8013 ( .A(n1539), .B(n5779), .C(n912), .D(n6133), .Y(n9008) );
  AOI22X1 U8014 ( .A(n5276), .B(n9500), .C(n5929), .D(n10502), .Y(n9006) );
  AOI22X1 U8015 ( .A(n391), .B(n6117), .C(n591), .D(n6135), .Y(n9005) );
  MUX2X1 U8016 ( .B(n6090), .A(n6067), .S(n6228), .Y(n9010) );
  MUX2X1 U8017 ( .B(n6088), .A(n2940), .S(n5274), .Y(n9014) );
  AOI22X1 U8018 ( .A(n447), .B(n5839), .C(n768), .D(n6137), .Y(n9012) );
  AOI22X1 U8019 ( .A(n712), .B(n6119), .C(n2269), .D(n5838), .Y(n9016) );
  AOI22X1 U8020 ( .A(n2590), .B(n5831), .C(n2911), .D(n5829), .Y(n9015) );
  NOR3X1 U8021 ( .A(n4023), .B(n4188), .C(n4610), .Y(n9018) );
  AOI22X1 U8022 ( .A(n2988), .B(n6141), .C(n1812), .D(n5783), .Y(n9025) );
  AOI22X1 U8023 ( .A(n1587), .B(n6147), .C(n6039), .D(n6112), .Y(n9024) );
  AOI22X1 U8024 ( .A(n2815), .B(n6110), .C(n2494), .D(n6115), .Y(n9022) );
  NAND3X1 U8025 ( .A(n2626), .B(n3031), .C(n9023), .Y(n9026) );
  AOI22X1 U8026 ( .A(n3779), .B(n6108), .C(n3458), .D(n6106), .Y(n9032) );
  AOI22X1 U8027 ( .A(n1331), .B(n5772), .C(n817), .D(n6145), .Y(n9029) );
  NAND3X1 U8028 ( .A(n5335), .B(n5356), .C(n9030), .Y(n9085) );
  AOI21X1 U8029 ( .A(n6000), .B(n5800), .C(n9033), .Y(n9034) );
  AOI22X1 U8030 ( .A(n5879), .B(n10072), .C(n6625), .D(n4992), .Y(n9045) );
  AOI21X1 U8031 ( .A(n8610), .B(n6325), .C(n9037), .Y(n9038) );
  AOI22X1 U8032 ( .A(n10500), .B(n5098), .C(n8679), .D(n4924), .Y(n9044) );
  AOI22X1 U8033 ( .A(n3554), .B(n5830), .C(n3875), .D(n5828), .Y(n9042) );
  AOI22X1 U8034 ( .A(n3233), .B(n5827), .C(n1765), .D(n5777), .Y(n9041) );
  AOI22X1 U8035 ( .A(n5740), .B(n9460), .C(n8738), .D(n5236), .Y(n9048) );
  AOI22X1 U8036 ( .A(n8891), .B(n5086), .C(n9046), .D(n5168), .Y(n9047) );
  OAI21X1 U8037 ( .A(n6004), .B(n6091), .C(n6089), .Y(n9049) );
  OAI21X1 U8038 ( .A(n6340), .B(n5729), .C(n5452), .Y(n9186) );
  AOI21X1 U8039 ( .A(n46), .B(n9049), .C(n9186), .Y(n9058) );
  OAI21X1 U8040 ( .A(n6010), .B(n5727), .C(n5465), .Y(n9051) );
  AOI21X1 U8041 ( .A(n9114), .B(n6330), .C(n9051), .Y(n9054) );
  AOI22X1 U8042 ( .A(n5788), .B(n6337), .C(n9175), .D(n5272), .Y(n9053) );
  AOI22X1 U8043 ( .A(n9114), .B(n6018), .C(n9310), .D(n6016), .Y(n9052) );
  MUX2X1 U8044 ( .B(n2769), .A(n9334), .S(n6232), .Y(n9055) );
  AOI22X1 U8045 ( .A(n5146), .B(n6073), .C(n9055), .D(n5733), .Y(n9056) );
  NOR3X1 U8046 ( .A(n4028), .B(n4268), .C(n4492), .Y(n9077) );
  AOI22X1 U8047 ( .A(n1026), .B(n5786), .C(n1283), .D(n5785), .Y(n9064) );
  AOI22X1 U8048 ( .A(n1540), .B(n5779), .C(n913), .D(n6133), .Y(n9063) );
  AOI22X1 U8049 ( .A(n5286), .B(n9500), .C(n5931), .D(n10502), .Y(n9061) );
  AOI22X1 U8050 ( .A(n376), .B(n6117), .C(n592), .D(n5823), .Y(n9060) );
  NAND3X1 U8051 ( .A(n2627), .B(n5500), .C(n9062), .Y(n9075) );
  NAND3X1 U8052 ( .A(n9310), .B(n5589), .C(n6233), .Y(n9065) );
  MUX2X1 U8053 ( .B(n6091), .A(n6068), .S(n46), .Y(n9066) );
  AOI21X1 U8054 ( .A(n9168), .B(n9310), .C(n9066), .Y(n9067) );
  NAND3X1 U8055 ( .A(n9509), .B(n6085), .C(n3646), .Y(n9068) );
  MUX2X1 U8056 ( .B(n5832), .A(n2799), .S(n6004), .Y(n9071) );
  AOI22X1 U8057 ( .A(n448), .B(n6131), .C(n769), .D(n5825), .Y(n9069) );
  AOI22X1 U8058 ( .A(n697), .B(n6119), .C(n2270), .D(n6104), .Y(n9073) );
  AOI22X1 U8059 ( .A(n2591), .B(n5831), .C(n2912), .D(n5829), .Y(n9072) );
  NOR3X1 U8060 ( .A(n4033), .B(n4192), .C(n4611), .Y(n9076) );
  AOI22X1 U8061 ( .A(n2989), .B(n6141), .C(n1813), .D(n5783), .Y(n9083) );
  AOI22X1 U8062 ( .A(n1588), .B(n5784), .C(n6042), .D(n6112), .Y(n9082) );
  AOI22X1 U8063 ( .A(n2816), .B(n6110), .C(n2495), .D(n6115), .Y(n9080) );
  NAND3X1 U8064 ( .A(n2628), .B(n3032), .C(n9081), .Y(n9084) );
  AOI22X1 U8065 ( .A(n3780), .B(n6108), .C(n3459), .D(n5774), .Y(n9090) );
  AOI22X1 U8066 ( .A(n1332), .B(n5772), .C(n818), .D(n6145), .Y(n9087) );
  NAND3X1 U8067 ( .A(n5351), .B(n5381), .C(n9088), .Y(n9160) );
  AOI22X1 U8068 ( .A(n914), .B(n5824), .C(n6018), .D(n9500), .Y(n9093) );
  AOI22X1 U8069 ( .A(n377), .B(n6117), .C(n593), .D(n5823), .Y(n9091) );
  NAND3X1 U8070 ( .A(n5435), .B(n3282), .C(n3581), .Y(n9098) );
  AOI22X1 U8071 ( .A(n3234), .B(n5827), .C(n1766), .D(n5777), .Y(n9096) );
  AOI22X1 U8072 ( .A(n1284), .B(n5785), .C(n1541), .D(n6123), .Y(n9094) );
  NAND3X1 U8073 ( .A(n5532), .B(n5677), .C(n5622), .Y(n9097) );
  MUX2X1 U8074 ( .B(n6090), .A(n6067), .S(n20), .Y(n9099) );
  MUX2X1 U8075 ( .B(n5832), .A(n5326), .S(n10), .Y(n9103) );
  AOI22X1 U8076 ( .A(n770), .B(n5825), .C(n5993), .D(n9969), .Y(n9101) );
  NAND3X1 U8077 ( .A(n9103), .B(n3283), .C(n3582), .Y(n9108) );
  AOI22X1 U8078 ( .A(n698), .B(n6119), .C(n2271), .D(n6104), .Y(n9106) );
  AOI22X1 U8079 ( .A(n2913), .B(n5829), .C(n449), .D(n5839), .Y(n9104) );
  NAND3X1 U8080 ( .A(n2629), .B(n3284), .C(n3583), .Y(n9107) );
  AOI21X1 U8081 ( .A(n5788), .B(n6334), .C(n9255), .Y(n9110) );
  OAI21X1 U8082 ( .A(n6014), .B(n5727), .C(n1908), .Y(n9125) );
  NAND3X1 U8083 ( .A(n6004), .B(n5819), .C(n9114), .Y(n9111) );
  OAI21X1 U8084 ( .A(n10104), .B(n4804), .C(n1909), .Y(n9112) );
  AOI21X1 U8085 ( .A(n10291), .B(n9125), .C(n9112), .Y(n9120) );
  AOI21X1 U8086 ( .A(n9310), .B(n6336), .C(n2373), .Y(n9117) );
  OAI21X1 U8087 ( .A(n6337), .B(n4803), .C(n4842), .Y(n9115) );
  NAND3X1 U8088 ( .A(n4842), .B(n5727), .C(n3671), .Y(n9118) );
  AOI22X1 U8089 ( .A(n9387), .B(n10290), .C(n9385), .D(n10291), .Y(n9119) );
  MUX2X1 U8090 ( .B(n2770), .A(n2784), .S(n6232), .Y(n9121) );
  NOR3X1 U8091 ( .A(n4125), .B(n9121), .C(n9186), .Y(n9134) );
  OAI21X1 U8092 ( .A(n10), .B(n6091), .C(n6089), .Y(n9123) );
  AOI22X1 U8093 ( .A(n19), .B(n9123), .C(n5074), .D(n6073), .Y(n9133) );
  OAI21X1 U8094 ( .A(n9124), .B(n9125), .C(n9168), .Y(n9126) );
  OAI21X1 U8095 ( .A(n9128), .B(n5571), .C(n9126), .Y(n9129) );
  AOI21X1 U8096 ( .A(n5837), .B(n5791), .C(n9129), .Y(n9131) );
  AOI22X1 U8097 ( .A(n6721), .B(n9389), .C(n8891), .D(n5165), .Y(n9130) );
  NAND3X1 U8098 ( .A(n9134), .B(n3033), .C(n9132), .Y(n9149) );
  AOI21X1 U8099 ( .A(n5768), .B(n6325), .C(n9135), .Y(n9136) );
  AOI22X1 U8100 ( .A(n10500), .B(n4764), .C(n8679), .D(n4995), .Y(n9141) );
  AOI22X1 U8101 ( .A(n3555), .B(n6092), .C(n3876), .D(n6096), .Y(n9140) );
  AOI22X1 U8102 ( .A(n9046), .B(n4877), .C(n5834), .D(n9379), .Y(n9147) );
  AOI21X1 U8103 ( .A(n5274), .B(n9626), .C(n5714), .Y(n9144) );
  OAI21X1 U8104 ( .A(n6062), .B(n6324), .C(n1910), .Y(n9380) );
  AOI22X1 U8105 ( .A(n6625), .B(n9380), .C(n10375), .D(n9388), .Y(n9145) );
  NOR3X1 U8106 ( .A(n4034), .B(n4269), .C(n4496), .Y(n9150) );
  NAND3X1 U8107 ( .A(n2740), .B(n3285), .C(n9150), .Y(n9153) );
  AOI22X1 U8108 ( .A(n2961), .B(n6141), .C(n1814), .D(n6149), .Y(n9158) );
  AOI22X1 U8109 ( .A(n1589), .B(n5784), .C(n6046), .D(n6112), .Y(n9157) );
  AOI22X1 U8110 ( .A(n2817), .B(n6110), .C(n2496), .D(n5781), .Y(n9155) );
  NAND3X1 U8111 ( .A(n2630), .B(n3034), .C(n9156), .Y(n9159) );
  AOI22X1 U8112 ( .A(n3781), .B(n6108), .C(n3460), .D(n5774), .Y(n9165) );
  AOI22X1 U8113 ( .A(n1333), .B(n5772), .C(n819), .D(n6145), .Y(n9162) );
  NAND3X1 U8114 ( .A(n5371), .B(n5428), .C(n9163), .Y(n9234) );
  AOI22X1 U8115 ( .A(n5788), .B(n5286), .C(n9175), .D(n6018), .Y(n9167) );
  AOI22X1 U8116 ( .A(n9114), .B(n6011), .C(n9310), .D(n6008), .Y(n9166) );
  MUX2X1 U8117 ( .B(n5272), .A(n6337), .S(n9310), .Y(n9169) );
  MUX2X1 U8118 ( .B(n6337), .A(n5272), .S(n46), .Y(n9170) );
  AOI22X1 U8119 ( .A(n5708), .B(n10291), .C(n6090), .D(n6333), .Y(n9171) );
  NAND3X1 U8120 ( .A(n2741), .B(n6089), .C(n3584), .Y(n9173) );
  AOI22X1 U8121 ( .A(n2990), .B(n5105), .C(n6232), .D(n3374), .Y(n9182) );
  NAND3X1 U8122 ( .A(n2742), .B(n3286), .C(n5727), .Y(n9178) );
  AOI21X1 U8123 ( .A(n9310), .B(n6333), .C(n2349), .Y(n9457) );
  AOI22X1 U8124 ( .A(n4958), .B(n9309), .C(n9179), .D(n6221), .Y(n9180) );
  OAI21X1 U8125 ( .A(n8171), .B(n9185), .C(n5367), .Y(n9190) );
  NAND3X1 U8126 ( .A(n5798), .B(n7491), .C(n5194), .Y(n9189) );
  NOR3X1 U8127 ( .A(n4035), .B(n9190), .C(n4500), .Y(n9226) );
  AOI22X1 U8128 ( .A(n8679), .B(n4852), .C(n3556), .D(n5830), .Y(n9197) );
  AOI22X1 U8129 ( .A(n3877), .B(n5828), .C(n3235), .D(n5827), .Y(n9196) );
  AOI22X1 U8130 ( .A(n7172), .B(n9458), .C(n9046), .D(n5033), .Y(n9203) );
  AOI22X1 U8131 ( .A(n5888), .B(n6331), .C(shift_amount[3]), .D(n1), .Y(n9198)
         );
  AOI22X1 U8132 ( .A(n6625), .B(n4765), .C(n10500), .D(n5046), .Y(n9201) );
  NAND3X1 U8133 ( .A(n2631), .B(n3287), .C(n3585), .Y(n9204) );
  MUX2X1 U8134 ( .B(n6090), .A(n6067), .S(n6232), .Y(n9206) );
  MUX2X1 U8135 ( .B(n5832), .A(n5420), .S(n6008), .Y(n9210) );
  AOI22X1 U8136 ( .A(n771), .B(n5825), .C(n6315), .D(n9969), .Y(n9208) );
  NAND3X1 U8137 ( .A(n9210), .B(n3289), .C(n3586), .Y(n9215) );
  AOI22X1 U8138 ( .A(n699), .B(n6119), .C(n2272), .D(n5838), .Y(n9213) );
  AOI22X1 U8139 ( .A(n2914), .B(n5829), .C(n450), .D(n5839), .Y(n9211) );
  NAND3X1 U8140 ( .A(n2632), .B(n3290), .C(n3587), .Y(n9214) );
  AOI22X1 U8141 ( .A(n6337), .B(n9500), .C(n5938), .D(n10502), .Y(n9217) );
  AOI22X1 U8142 ( .A(n378), .B(n6117), .C(n594), .D(n5823), .Y(n9216) );
  AOI22X1 U8143 ( .A(n1767), .B(n5777), .C(n1028), .D(n5786), .Y(n9220) );
  AOI22X1 U8144 ( .A(n1542), .B(n5779), .C(n915), .D(n6133), .Y(n9218) );
  NAND3X1 U8145 ( .A(n2633), .B(n5379), .C(n5432), .Y(n9221) );
  NOR3X1 U8146 ( .A(n9223), .B(n4270), .C(n4503), .Y(n9224) );
  NAND3X1 U8147 ( .A(n9226), .B(n3288), .C(n9224), .Y(n9227) );
  AOI22X1 U8148 ( .A(n2962), .B(n6141), .C(n1815), .D(n5783), .Y(n9232) );
  AOI22X1 U8149 ( .A(n1590), .B(n5784), .C(n21), .D(n6112), .Y(n9231) );
  AOI22X1 U8150 ( .A(n2818), .B(n6110), .C(n2497), .D(n5781), .Y(n9229) );
  NAND3X1 U8151 ( .A(n2634), .B(n5558), .C(n9230), .Y(n9233) );
  AOI22X1 U8152 ( .A(n3782), .B(n6108), .C(n3461), .D(n5774), .Y(n9239) );
  AOI22X1 U8153 ( .A(n1334), .B(n5772), .C(n820), .D(n6145), .Y(n9236) );
  NAND3X1 U8154 ( .A(n5418), .B(n5486), .C(n9237), .Y(n9296) );
  AOI22X1 U8155 ( .A(n8891), .B(n5089), .C(n7172), .D(n5238), .Y(n9249) );
  AOI22X1 U8156 ( .A(n9046), .B(n5053), .C(n10500), .D(n5155), .Y(n9248) );
  AOI22X1 U8157 ( .A(n8679), .B(n4927), .C(n3557), .D(n6092), .Y(n9246) );
  AOI22X1 U8158 ( .A(n3878), .B(n6096), .C(n3236), .D(n5827), .Y(n9245) );
  OAI21X1 U8159 ( .A(n5656), .B(n5450), .C(n5588), .Y(n9253) );
  NAND3X1 U8160 ( .A(n2743), .B(n5398), .C(n5756), .Y(n9252) );
  AOI22X1 U8161 ( .A(n5762), .B(n9253), .C(n5272), .D(n3375), .Y(n9257) );
  AOI22X1 U8162 ( .A(n5788), .B(n5270), .C(n9175), .D(n6328), .Y(n9254) );
  AOI22X1 U8163 ( .A(n9460), .B(n5200), .C(n9309), .D(n4818), .Y(n9256) );
  OAI21X1 U8164 ( .A(n6334), .B(n6091), .C(n6089), .Y(n9259) );
  AOI21X1 U8165 ( .A(n6234), .B(n9259), .C(n9258), .Y(n9271) );
  NAND3X1 U8166 ( .A(n4739), .B(n9263), .C(n4971), .Y(n9492) );
  AOI22X1 U8167 ( .A(n5788), .B(n6018), .C(n9175), .D(n5282), .Y(n9265) );
  NAND3X1 U8168 ( .A(n2744), .B(n4873), .C(n3588), .Y(n9268) );
  AOI22X1 U8169 ( .A(n4902), .B(n5628), .C(n3366), .D(n5105), .Y(n9269) );
  NOR3X1 U8170 ( .A(n4039), .B(n4271), .C(n4504), .Y(n9288) );
  AOI22X1 U8171 ( .A(n2273), .B(n6104), .C(n2594), .D(n6102), .Y(n9280) );
  AOI22X1 U8172 ( .A(n2915), .B(n5829), .C(n451), .D(n5839), .Y(n9279) );
  AOI22X1 U8173 ( .A(n772), .B(n5825), .C(n5276), .D(n9969), .Y(n9277) );
  MUX2X1 U8174 ( .B(n6091), .A(n6068), .S(n6234), .Y(n9273) );
  MUX2X1 U8175 ( .B(n10522), .A(n5537), .S(n5269), .Y(n9275) );
  AOI21X1 U8176 ( .A(n1077), .B(n6127), .C(n9275), .Y(n9276) );
  AOI22X1 U8177 ( .A(n5941), .B(n6098), .C(n379), .D(n5778), .Y(n9282) );
  AOI22X1 U8178 ( .A(n595), .B(n6135), .C(n700), .D(n5790), .Y(n9281) );
  AOI22X1 U8179 ( .A(n1768), .B(n5777), .C(n1029), .D(n6129), .Y(n9285) );
  AOI22X1 U8180 ( .A(n1543), .B(n5779), .C(n916), .D(n6133), .Y(n9283) );
  NOR3X1 U8181 ( .A(n4044), .B(n4272), .C(n4508), .Y(n9287) );
  AOI22X1 U8182 ( .A(n2991), .B(n6141), .C(n1816), .D(n5783), .Y(n9294) );
  AOI22X1 U8183 ( .A(n1591), .B(n5784), .C(n6351), .D(n6112), .Y(n9293) );
  AOI22X1 U8184 ( .A(n2819), .B(n6110), .C(n2498), .D(n5781), .Y(n9291) );
  NAND3X1 U8185 ( .A(n2635), .B(n5343), .C(n9292), .Y(n9295) );
  AOI22X1 U8186 ( .A(n3783), .B(n6108), .C(n3462), .D(n6106), .Y(n9301) );
  AOI22X1 U8187 ( .A(n1335), .B(n5772), .C(n821), .D(n6145), .Y(n9298) );
  NAND3X1 U8188 ( .A(n5474), .B(n5549), .C(n9299), .Y(n9359) );
  AOI22X1 U8189 ( .A(n917), .B(n5824), .C(n5942), .D(n10502), .Y(n9303) );
  AOI22X1 U8190 ( .A(n380), .B(n6117), .C(n596), .D(n5823), .Y(n9302) );
  AOI22X1 U8191 ( .A(n3237), .B(n5827), .C(n1769), .D(n6121), .Y(n9306) );
  AOI22X1 U8192 ( .A(n1287), .B(n6125), .C(n1544), .D(n5779), .Y(n9304) );
  NAND3X1 U8193 ( .A(n5373), .B(n5684), .C(n5623), .Y(n9307) );
  OAI21X1 U8194 ( .A(n5450), .B(n5637), .C(n5732), .Y(n9311) );
  MUX2X1 U8195 ( .B(n6090), .A(n6067), .S(n5280), .Y(n9312) );
  NAND3X1 U8196 ( .A(n9443), .B(n9312), .C(n9441), .Y(n9313) );
  MUX2X1 U8197 ( .B(n5832), .A(n2800), .S(n5286), .Y(n9316) );
  AOI22X1 U8198 ( .A(n773), .B(n5825), .C(n43), .D(n9969), .Y(n9314) );
  NAND3X1 U8199 ( .A(n9316), .B(n5561), .C(n5493), .Y(n9321) );
  AOI22X1 U8200 ( .A(n701), .B(n6119), .C(n2274), .D(n5838), .Y(n9319) );
  AOI22X1 U8201 ( .A(n2916), .B(n6086), .C(n452), .D(n5839), .Y(n9317) );
  NAND3X1 U8202 ( .A(n2636), .B(n3291), .C(n3589), .Y(n9320) );
  AOI21X1 U8203 ( .A(n9309), .B(n9114), .C(n5749), .Y(n9322) );
  OAI21X1 U8204 ( .A(n9324), .B(n5654), .C(n5272), .Y(n9327) );
  AOI22X1 U8205 ( .A(n5762), .B(n10290), .C(n10375), .D(n5271), .Y(n9325) );
  NAND3X1 U8206 ( .A(n9327), .B(n5452), .C(n3590), .Y(n9454) );
  AOI21X1 U8207 ( .A(n6011), .B(n5185), .C(n5042), .Y(n9341) );
  AOI21X1 U8208 ( .A(n9309), .B(n5788), .C(n5751), .Y(n9328) );
  AOI21X1 U8209 ( .A(n9309), .B(n9175), .C(n5750), .Y(n9330) );
  AOI22X1 U8210 ( .A(n6332), .B(n5223), .C(n6007), .D(n5217), .Y(n9340) );
  OAI21X1 U8211 ( .A(n5286), .B(n6091), .C(n6089), .Y(n9332) );
  AOI22X1 U8212 ( .A(n6328), .B(n2780), .C(n5279), .D(n9332), .Y(n9338) );
  AOI22X1 U8213 ( .A(n5216), .B(n6073), .C(n5105), .D(n4828), .Y(n9337) );
  AOI22X1 U8214 ( .A(n9046), .B(n4924), .C(n10500), .D(n4992), .Y(n9343) );
  AOI22X1 U8215 ( .A(n3558), .B(n5830), .C(n3879), .D(n5828), .Y(n9342) );
  AOI22X1 U8216 ( .A(n5740), .B(n5805), .C(n9460), .D(n5168), .Y(n9347) );
  AOI22X1 U8217 ( .A(n8891), .B(n5236), .C(n7172), .D(n5098), .Y(n9345) );
  NOR3X1 U8218 ( .A(n4049), .B(n4273), .C(n4512), .Y(n9349) );
  NAND3X1 U8219 ( .A(n2745), .B(n3292), .C(n9349), .Y(n9352) );
  AOI22X1 U8220 ( .A(n2963), .B(n6141), .C(n1817), .D(n6149), .Y(n9357) );
  AOI22X1 U8221 ( .A(n1592), .B(n5784), .C(n6053), .D(n6112), .Y(n9356) );
  AOI22X1 U8222 ( .A(n2820), .B(n6110), .C(n2499), .D(n5781), .Y(n9354) );
  NAND3X1 U8223 ( .A(n2637), .B(n3035), .C(n9355), .Y(n9358) );
  AOI22X1 U8224 ( .A(n3784), .B(n5775), .C(n3463), .D(n6106), .Y(n9364) );
  AOI22X1 U8225 ( .A(n1336), .B(n5772), .C(n822), .D(n6145), .Y(n9361) );
  NAND3X1 U8226 ( .A(n5530), .B(n5616), .C(n9362), .Y(n9423) );
  AOI22X1 U8227 ( .A(n5285), .B(n5223), .C(n6008), .D(n5217), .Y(n9370) );
  OAI21X1 U8228 ( .A(n9500), .B(n9365), .C(n6330), .Y(n9369) );
  OAI21X1 U8229 ( .A(n6018), .B(n6091), .C(n6089), .Y(n9367) );
  AOI22X1 U8230 ( .A(n6237), .B(n9367), .C(n5791), .D(n9366), .Y(n9368) );
  NAND3X1 U8231 ( .A(n2638), .B(n9369), .C(n3591), .Y(n9377) );
  NAND3X1 U8232 ( .A(n9114), .B(n6004), .C(n9498), .Y(n9374) );
  AOI22X1 U8233 ( .A(n9371), .B(n9372), .C(n5286), .D(n5185), .Y(n9373) );
  NAND3X1 U8234 ( .A(n9375), .B(n3056), .C(n3592), .Y(n9376) );
  AOI22X1 U8235 ( .A(n7351), .B(n5714), .C(n9046), .D(n4995), .Y(n9383) );
  AOI22X1 U8236 ( .A(n10500), .B(n9380), .C(n3559), .D(n5830), .Y(n9381) );
  NAND3X1 U8237 ( .A(n2639), .B(n3293), .C(n3593), .Y(n9394) );
  AOI22X1 U8238 ( .A(n5798), .B(n9386), .C(n9385), .D(n9384), .Y(n9392) );
  AOI22X1 U8239 ( .A(n5822), .B(n9389), .C(n7147), .D(n9388), .Y(n9390) );
  NAND3X1 U8240 ( .A(n2640), .B(n3294), .C(n3594), .Y(n9393) );
  MUX2X1 U8241 ( .B(n6090), .A(n6067), .S(n6237), .Y(n9395) );
  NAND3X1 U8242 ( .A(n9443), .B(n9395), .C(n9441), .Y(n9396) );
  MUX2X1 U8243 ( .B(n5832), .A(n2801), .S(n6018), .Y(n9399) );
  AOI22X1 U8244 ( .A(n774), .B(n5825), .C(n6319), .D(n9969), .Y(n9397) );
  NAND3X1 U8245 ( .A(n9399), .B(n3296), .C(n3595), .Y(n9404) );
  AOI22X1 U8246 ( .A(n702), .B(n6119), .C(n2275), .D(n5838), .Y(n9402) );
  AOI22X1 U8247 ( .A(n2917), .B(n5829), .C(n453), .D(n5839), .Y(n9400) );
  NAND3X1 U8248 ( .A(n2641), .B(n3297), .C(n3597), .Y(n9403) );
  AOI22X1 U8249 ( .A(n1545), .B(n5779), .C(n918), .D(n6133), .Y(n9407) );
  AOI22X1 U8250 ( .A(n381), .B(n6117), .C(n597), .D(n5823), .Y(n9405) );
  AOI22X1 U8251 ( .A(n3880), .B(n6096), .C(n3238), .D(n5827), .Y(n9410) );
  AOI22X1 U8252 ( .A(n1031), .B(n6129), .C(n1288), .D(n5785), .Y(n9408) );
  NOR3X1 U8253 ( .A(n9412), .B(n4196), .C(n39), .Y(n9413) );
  NAND3X1 U8254 ( .A(n2746), .B(n3295), .C(n9413), .Y(n9416) );
  AOI22X1 U8255 ( .A(n138), .B(n6141), .C(n1818), .D(n5783), .Y(n9421) );
  AOI22X1 U8256 ( .A(n1593), .B(n5784), .C(n6354), .D(n6112), .Y(n9420) );
  AOI22X1 U8257 ( .A(n2821), .B(n6110), .C(n2500), .D(n5781), .Y(n9418) );
  NAND3X1 U8258 ( .A(n9419), .B(n3036), .C(n129), .Y(n9422) );
  OR2X2 U8259 ( .A(n2036), .B(n115), .Y(result[18]) );
  AOI22X1 U8260 ( .A(n2597), .B(n5831), .C(n2918), .D(n5829), .Y(n9428) );
  OAI21X1 U8261 ( .A(n6095), .B(n6324), .C(n5368), .Y(n9425) );
  AOI21X1 U8262 ( .A(n1080), .B(n5826), .C(n9425), .Y(n9426) );
  AOI22X1 U8263 ( .A(n598), .B(n6135), .C(n703), .D(n5790), .Y(n9430) );
  AOI22X1 U8264 ( .A(n919), .B(n5824), .C(n6008), .D(n9500), .Y(n9432) );
  AOI22X1 U8265 ( .A(n6290), .B(n10502), .C(n382), .D(n5778), .Y(n9431) );
  NOR3X1 U8266 ( .A(n74), .B(n4274), .C(n4612), .Y(n9485) );
  AOI22X1 U8267 ( .A(n3785), .B(n6108), .C(n3464), .D(n6106), .Y(n9440) );
  AOI22X1 U8268 ( .A(n1337), .B(n5772), .C(n823), .D(n5771), .Y(n9437) );
  MUX2X1 U8269 ( .B(n6090), .A(n6067), .S(n6239), .Y(n9442) );
  NAND3X1 U8270 ( .A(n9443), .B(n9442), .C(n9441), .Y(n9444) );
  MUX2X1 U8271 ( .B(n5832), .A(n2802), .S(n6022), .Y(n9447) );
  AOI22X1 U8272 ( .A(n1594), .B(n5784), .C(n6356), .D(n10480), .Y(n9445) );
  AOI22X1 U8273 ( .A(n2822), .B(n6110), .C(n2501), .D(n6115), .Y(n9449) );
  NOR3X1 U8274 ( .A(n4055), .B(n4200), .C(n4613), .Y(n9484) );
  AOI21X1 U8275 ( .A(n6090), .B(n6339), .C(n10564), .Y(n9452) );
  AOI22X1 U8276 ( .A(n5286), .B(n5223), .C(n5269), .D(n5217), .Y(n9451) );
  OAI21X1 U8277 ( .A(n2762), .B(n6240), .C(n1885), .Y(n9456) );
  NAND3X1 U8278 ( .A(n5789), .B(n10487), .C(n6221), .Y(n9453) );
  OAI21X1 U8279 ( .A(n169), .B(n6336), .C(n1911), .Y(n9455) );
  NOR3X1 U8280 ( .A(n9456), .B(n9455), .C(n5042), .Y(n9467) );
  AOI22X1 U8281 ( .A(n8485), .B(n9458), .C(n4958), .D(n9498), .Y(n9459) );
  OAI21X1 U8282 ( .A(n163), .B(n5701), .C(n1886), .Y(n9465) );
  AOI22X1 U8283 ( .A(n9461), .B(n10505), .C(n5860), .D(n10491), .Y(n9463) );
  AOI22X1 U8284 ( .A(n8952), .B(n5798), .C(n5805), .D(n5178), .Y(n9462) );
  AOI22X1 U8285 ( .A(n3881), .B(n5828), .C(n3239), .D(n5827), .Y(n9472) );
  AOI22X1 U8286 ( .A(n1032), .B(n5786), .C(n1289), .D(n5785), .Y(n9469) );
  NAND3X1 U8287 ( .A(n2642), .B(n3298), .C(n9470), .Y(n9481) );
  AOI22X1 U8288 ( .A(n9384), .B(n5708), .C(n9168), .D(n9473), .Y(n9480) );
  AOI22X1 U8289 ( .A(n152), .B(n7351), .C(n7172), .D(n5046), .Y(n9479) );
  OAI21X1 U8290 ( .A(n9475), .B(n5721), .C(n1936), .Y(n9477) );
  AOI21X1 U8291 ( .A(n3560), .B(n6092), .C(n9477), .Y(n9478) );
  NOR3X1 U8292 ( .A(n4126), .B(n145), .C(n4517), .Y(n9483) );
  NAND3X1 U8293 ( .A(n9485), .B(n9484), .C(n9483), .Y(n9486) );
  AOI22X1 U8294 ( .A(n3786), .B(n6108), .C(n3465), .D(n6106), .Y(n9491) );
  AOI22X1 U8295 ( .A(n1338), .B(n5772), .C(n824), .D(n6145), .Y(n9488) );
  NAND3X1 U8296 ( .A(n5602), .B(n5682), .C(n9489), .Y(n9543) );
  AOI22X1 U8297 ( .A(n3882), .B(n5828), .C(n2598), .D(n5831), .Y(n9520) );
  AOI22X1 U8298 ( .A(n4902), .B(n10574), .C(n9046), .D(n4927), .Y(n9495) );
  AOI22X1 U8299 ( .A(n6018), .B(n5223), .C(n6022), .D(n5185), .Y(n9493) );
  OAI21X1 U8300 ( .A(n156), .B(n5698), .C(n1937), .Y(n9507) );
  AOI22X1 U8301 ( .A(n5948), .B(n6098), .C(n6003), .D(n6094), .Y(n9499) );
  OAI21X1 U8302 ( .A(n5519), .B(n5273), .C(n1887), .Y(n9501) );
  AOI21X1 U8303 ( .A(n8485), .B(n5238), .C(n9501), .Y(n9506) );
  OAI21X1 U8304 ( .A(n5271), .B(n6091), .C(n6089), .Y(n9503) );
  AOI22X1 U8305 ( .A(n6241), .B(n9503), .C(n7172), .D(n5155), .Y(n9505) );
  NOR3X1 U8306 ( .A(n4059), .B(n9507), .C(n4522), .Y(n9516) );
  AOI21X1 U8307 ( .A(n9250), .B(n5798), .C(n9508), .Y(n9512) );
  MUX2X1 U8308 ( .B(n5818), .A(n6067), .S(n6241), .Y(n9511) );
  NOR3X1 U8309 ( .A(n5265), .B(n5263), .C(n4857), .Y(n9510) );
  NAND3X1 U8310 ( .A(n2705), .B(n9511), .C(n9510), .Y(n9513) );
  MUX2X1 U8311 ( .B(n5832), .A(n2803), .S(n5271), .Y(n9515) );
  NAND3X1 U8312 ( .A(n9516), .B(n9515), .C(n3672), .Y(n9517) );
  AOI21X1 U8313 ( .A(n3561), .B(n5830), .C(n2350), .Y(n9519) );
  AOI22X1 U8314 ( .A(n2919), .B(n5829), .C(n2277), .D(n5838), .Y(n9518) );
  NAND3X1 U8315 ( .A(n2643), .B(n3057), .C(n3598), .Y(n9521) );
  AOI21X1 U8316 ( .A(n599), .B(n5823), .C(n2351), .Y(n9524) );
  NAND3X1 U8317 ( .A(n2706), .B(n3299), .C(n3673), .Y(n9525) );
  AOI21X1 U8318 ( .A(n704), .B(n5790), .C(n2352), .Y(n9528) );
  NAND3X1 U8319 ( .A(n2707), .B(n3300), .C(n3674), .Y(n9529) );
  AOI21X1 U8320 ( .A(n1547), .B(n6123), .C(n2353), .Y(n9532) );
  NAND3X1 U8321 ( .A(n2708), .B(n3675), .C(n5685), .Y(n9533) );
  AOI21X1 U8322 ( .A(n1033), .B(n6129), .C(n122), .Y(n9535) );
  AOI22X1 U8323 ( .A(n140), .B(n6141), .C(n1820), .D(n5783), .Y(n9541) );
  AOI22X1 U8324 ( .A(n1595), .B(n5784), .C(n6061), .D(n10480), .Y(n9540) );
  AOI22X1 U8325 ( .A(n2823), .B(n6110), .C(n2502), .D(n5781), .Y(n9538) );
  NAND3X1 U8326 ( .A(n5437), .B(n130), .C(n9539), .Y(n9542) );
  OR2X2 U8327 ( .A(n2040), .B(n116), .Y(result[16]) );
  AOI22X1 U8328 ( .A(n3787), .B(n6108), .C(n3466), .D(n6106), .Y(n9548) );
  AOI22X1 U8329 ( .A(n1339), .B(n5772), .C(n825), .D(n6145), .Y(n9545) );
  NAND3X1 U8330 ( .A(n2644), .B(n5289), .C(n9546), .Y(n9603) );
  NAND3X1 U8331 ( .A(n4742), .B(n4786), .C(n4833), .Y(n9550) );
  NAND3X1 U8332 ( .A(n4743), .B(n9549), .C(n4972), .Y(n9847) );
  MUX2X1 U8333 ( .B(n2771), .A(n4965), .S(n6245), .Y(n9551) );
  AOI22X1 U8334 ( .A(n5769), .B(n6356), .C(n6060), .D(n9614), .Y(n9553) );
  AOI22X1 U8335 ( .A(n6354), .B(n9639), .C(n6055), .D(n9577), .Y(n9552) );
  AOI22X1 U8336 ( .A(n6049), .B(n5769), .C(n6351), .D(n9614), .Y(n9554) );
  AOI22X1 U8337 ( .A(n9792), .B(n5255), .C(n10034), .D(n5125), .Y(n9555) );
  OAI21X1 U8338 ( .A(n6247), .B(n9551), .C(n1888), .Y(n9558) );
  AOI22X1 U8339 ( .A(n5734), .B(n6077), .C(n21), .D(n6081), .Y(n9556) );
  AOI22X1 U8340 ( .A(n9558), .B(n9647), .C(n9774), .D(n5149), .Y(n9563) );
  AOI22X1 U8341 ( .A(n3562), .B(n6092), .C(n3883), .D(n5828), .Y(n9562) );
  AOI22X1 U8342 ( .A(n3241), .B(n5827), .C(n1741), .D(n5777), .Y(n9560) );
  AOI22X1 U8343 ( .A(n1002), .B(n5786), .C(n1259), .D(n5785), .Y(n9559) );
  AOI22X1 U8344 ( .A(n4959), .B(n10087), .C(n9565), .D(n5733), .Y(n9570) );
  OAI21X1 U8345 ( .A(n6245), .B(n10104), .C(n5007), .Y(n9568) );
  AOI22X1 U8346 ( .A(n6354), .B(n6077), .C(n6081), .D(n6356), .Y(n9567) );
  AOI22X1 U8347 ( .A(n6061), .B(n6079), .C(n6054), .D(n9688), .Y(n9566) );
  AOI22X1 U8348 ( .A(n5746), .B(n9568), .C(n5742), .D(n5207), .Y(n9569) );
  AOI22X1 U8349 ( .A(n6032), .B(n9793), .C(n6029), .D(n6065), .Y(n9573) );
  OAI21X1 U8350 ( .A(n59), .B(n6091), .C(n6089), .Y(n9571) );
  AOI22X1 U8351 ( .A(n6026), .B(n6066), .C(n70), .D(n9571), .Y(n9572) );
  NOR3X1 U8352 ( .A(n4063), .B(n4275), .C(n4614), .Y(n9595) );
  AOI22X1 U8353 ( .A(n2599), .B(n5831), .C(n2920), .D(n5829), .Y(n9586) );
  AOI22X1 U8354 ( .A(n424), .B(n6131), .C(n745), .D(n5825), .Y(n9585) );
  AOI22X1 U8355 ( .A(n6043), .B(n6094), .C(n1082), .D(n6127), .Y(n9583) );
  NAND3X1 U8356 ( .A(n4744), .B(n5724), .C(n6085), .Y(n10520) );
  MUX2X1 U8357 ( .B(n6091), .A(n6068), .S(n70), .Y(n9579) );
  OAI21X1 U8358 ( .A(n4758), .B(n5011), .C(n6070), .Y(n9578) );
  NAND3X1 U8359 ( .A(n5736), .B(n10447), .C(n3676), .Y(n9581) );
  MUX2X1 U8360 ( .B(n5832), .A(n2804), .S(n59), .Y(n9582) );
  NAND3X1 U8361 ( .A(n5489), .B(n3037), .C(n9584), .Y(n9593) );
  AOI22X1 U8362 ( .A(n368), .B(n6117), .C(n600), .D(n5823), .Y(n9588) );
  AOI22X1 U8363 ( .A(n689), .B(n5790), .C(n2278), .D(n6104), .Y(n9587) );
  AOI22X1 U8364 ( .A(n1516), .B(n5779), .C(n921), .D(n5824), .Y(n9590) );
  AOI22X1 U8365 ( .A(n9500), .B(n5885), .C(n5952), .D(n10502), .Y(n9589) );
  NOR3X1 U8366 ( .A(n4068), .B(n4276), .C(n4615), .Y(n9594) );
  AOI22X1 U8367 ( .A(n2992), .B(n6141), .C(n1821), .D(n5783), .Y(n9601) );
  AOI22X1 U8368 ( .A(n1596), .B(n6147), .C(n5879), .D(n6112), .Y(n9600) );
  AOI22X1 U8369 ( .A(n2824), .B(n6110), .C(n2503), .D(n5781), .Y(n9598) );
  NAND3X1 U8370 ( .A(n2645), .B(n5359), .C(n9599), .Y(n9602) );
  AOI22X1 U8371 ( .A(n3788), .B(n5775), .C(n3467), .D(n6106), .Y(n9608) );
  AOI22X1 U8372 ( .A(n1340), .B(n5772), .C(n826), .D(n6145), .Y(n9605) );
  NAND3X1 U8373 ( .A(n2646), .B(n5292), .C(n9606), .Y(n9681) );
  MUX2X1 U8374 ( .B(n6026), .A(n59), .S(n70), .Y(n9609) );
  AOI21X1 U8375 ( .A(n9577), .B(n6026), .C(n9783), .Y(n9610) );
  NAND3X1 U8376 ( .A(n4745), .B(n4787), .C(n3647), .Y(n9611) );
  AOI22X1 U8377 ( .A(n10149), .B(n4946), .C(n3367), .D(n5212), .Y(n9617) );
  AOI21X1 U8378 ( .A(n9577), .B(n6033), .C(n2374), .Y(n9638) );
  NAND3X1 U8379 ( .A(n4843), .B(n4785), .C(n3677), .Y(n9648) );
  AOI22X1 U8380 ( .A(n6351), .B(n5769), .C(n6055), .D(n9614), .Y(n9615) );
  AOI22X1 U8381 ( .A(n5757), .B(n9919), .C(n5754), .D(n5128), .Y(n9616) );
  AOI22X1 U8382 ( .A(n5885), .B(n9793), .C(n6032), .D(n6065), .Y(n9622) );
  OAI21X1 U8383 ( .A(n6026), .B(n6091), .C(n6089), .Y(n9619) );
  OAI21X1 U8384 ( .A(n6341), .B(n6063), .C(n5528), .Y(n9908) );
  AOI22X1 U8385 ( .A(n6243), .B(n9619), .C(n5836), .D(n9916), .Y(n9620) );
  NAND3X1 U8386 ( .A(n2647), .B(n3301), .C(n3599), .Y(n9623) );
  AOI21X1 U8387 ( .A(n6356), .B(n9632), .C(n2375), .Y(n9627) );
  OAI21X1 U8388 ( .A(n6082), .B(n6359), .C(n4723), .Y(n10441) );
  OAI21X1 U8389 ( .A(n6153), .B(n6359), .C(n4723), .Y(n10440) );
  OAI21X1 U8390 ( .A(n9630), .B(n5731), .C(n1938), .Y(n10431) );
  AOI21X1 U8391 ( .A(n6083), .B(n6033), .C(n2376), .Y(n9635) );
  OAI21X1 U8392 ( .A(n6037), .B(n6078), .C(n4844), .Y(n9633) );
  AOI22X1 U8393 ( .A(n6731), .B(n10431), .C(n9921), .D(n10375), .Y(n9637) );
  NAND3X1 U8394 ( .A(n4844), .B(n6062), .C(n3678), .Y(n9644) );
  AOI22X1 U8395 ( .A(n8968), .B(n4947), .C(n3563), .D(n6092), .Y(n9636) );
  OAI21X1 U8396 ( .A(n6037), .B(n4805), .C(n4843), .Y(n9640) );
  AOI22X1 U8397 ( .A(n6356), .B(n9639), .C(n6354), .D(n9577), .Y(n9643) );
  AOI22X1 U8398 ( .A(n10487), .B(n5769), .C(n7491), .D(n6243), .Y(n9641) );
  OAI21X1 U8399 ( .A(n5766), .B(n3356), .C(n9642), .Y(n10438) );
  AOI22X1 U8400 ( .A(n9784), .B(n9920), .C(n9792), .D(n10438), .Y(n9651) );
  AOI21X1 U8401 ( .A(n6054), .B(n5800), .C(n10182), .Y(n9645) );
  AOI22X1 U8402 ( .A(n9774), .B(n5077), .C(n9767), .D(n4869), .Y(n9649) );
  NAND3X1 U8403 ( .A(n2648), .B(n3302), .C(n3600), .Y(n9652) );
  MUX2X1 U8404 ( .B(n6090), .A(n6067), .S(n6243), .Y(n9654) );
  NAND3X1 U8405 ( .A(n9654), .B(n6070), .C(n9803), .Y(n9655) );
  MUX2X1 U8406 ( .B(n6088), .A(n5352), .S(n6026), .Y(n9658) );
  AOI22X1 U8407 ( .A(n746), .B(n5825), .C(n6046), .D(n9969), .Y(n9656) );
  NAND3X1 U8408 ( .A(n9658), .B(n3304), .C(n3601), .Y(n9663) );
  AOI22X1 U8409 ( .A(n690), .B(n6119), .C(n2279), .D(n5838), .Y(n9661) );
  AOI22X1 U8410 ( .A(n2921), .B(n6086), .C(n425), .D(n5839), .Y(n9659) );
  NAND3X1 U8411 ( .A(n2649), .B(n3305), .C(n3602), .Y(n9662) );
  AOI22X1 U8412 ( .A(n9500), .B(n6034), .C(n5955), .D(n10502), .Y(n9665) );
  AOI22X1 U8413 ( .A(n369), .B(n6117), .C(n601), .D(n5823), .Y(n9664) );
  AOI22X1 U8414 ( .A(n3884), .B(n5828), .C(n3242), .D(n5827), .Y(n9668) );
  AOI22X1 U8415 ( .A(n1260), .B(n5785), .C(n922), .D(n6133), .Y(n9666) );
  NOR3X1 U8416 ( .A(n9670), .B(n4277), .C(n4526), .Y(n9671) );
  NAND3X1 U8417 ( .A(n2747), .B(n3303), .C(n9671), .Y(n9674) );
  AOI22X1 U8418 ( .A(n2964), .B(n6141), .C(n1822), .D(n5783), .Y(n9679) );
  AOI22X1 U8419 ( .A(n1597), .B(n5784), .C(n5992), .D(n6112), .Y(n9678) );
  AOI22X1 U8420 ( .A(n2825), .B(n6110), .C(n2504), .D(n5781), .Y(n9676) );
  NAND3X1 U8421 ( .A(n2650), .B(n3038), .C(n9677), .Y(n9680) );
  AOI22X1 U8422 ( .A(n3789), .B(n6108), .C(n3468), .D(n5774), .Y(n9686) );
  AOI22X1 U8423 ( .A(n1341), .B(n5772), .C(n827), .D(n6145), .Y(n9683) );
  NAND3X1 U8424 ( .A(n2651), .B(n5296), .C(n9684), .Y(n9759) );
  AOI22X1 U8425 ( .A(n6026), .B(n6077), .C(n6081), .D(n59), .Y(n9687) );
  OAI21X1 U8426 ( .A(n6343), .B(n6063), .C(n1889), .Y(n10504) );
  OAI21X1 U8427 ( .A(n6245), .B(n9846), .C(n5442), .Y(n10030) );
  AOI22X1 U8428 ( .A(n6072), .B(n10504), .C(n10030), .D(n5203), .Y(n9699) );
  NAND3X1 U8429 ( .A(n4747), .B(n4788), .C(n3679), .Y(n9694) );
  MUX2X1 U8430 ( .B(n6344), .A(n6346), .S(n70), .Y(n9695) );
  MUX2X1 U8431 ( .B(n6039), .A(n6037), .S(n9577), .Y(n9696) );
  AOI22X1 U8432 ( .A(n5757), .B(n9725), .C(n9784), .D(n9977), .Y(n9697) );
  NAND3X1 U8433 ( .A(n2652), .B(n3306), .C(n3603), .Y(n9709) );
  AOI22X1 U8434 ( .A(n6054), .B(n5769), .C(n6354), .D(n9614), .Y(n9700) );
  NAND3X1 U8435 ( .A(n7491), .B(n10034), .C(n5197), .Y(n9702) );
  OAI21X1 U8436 ( .A(n9703), .B(n6033), .C(n1912), .Y(n9704) );
  AOI21X1 U8437 ( .A(n5885), .B(n6065), .C(n9704), .Y(n9707) );
  OAI21X1 U8438 ( .A(n6029), .B(n6091), .C(n6089), .Y(n9705) );
  AOI22X1 U8439 ( .A(n6032), .B(n6066), .C(n6245), .D(n9705), .Y(n9706) );
  MUX2X1 U8440 ( .B(n6060), .A(n6356), .S(n9688), .Y(n10224) );
  MUX2X1 U8441 ( .B(n6039), .A(n6037), .S(n9688), .Y(n9710) );
  AOI22X1 U8442 ( .A(n6730), .B(n10506), .C(n10375), .D(n9978), .Y(n9715) );
  MUX2X1 U8443 ( .B(n6037), .A(n6039), .S(n5886), .Y(n9711) );
  AOI21X1 U8444 ( .A(n6043), .B(n9626), .C(n5649), .Y(n9712) );
  OAI21X1 U8445 ( .A(n6062), .B(n6348), .C(n1913), .Y(n9972) );
  AOI22X1 U8446 ( .A(n3564), .B(n6092), .C(n3885), .D(n6096), .Y(n9713) );
  NAND3X1 U8447 ( .A(n2653), .B(n3307), .C(n3604), .Y(n9730) );
  AOI22X1 U8448 ( .A(n6351), .B(n6077), .C(n6054), .D(n6081), .Y(n9717) );
  AOI22X1 U8449 ( .A(n6354), .B(n6079), .C(n6049), .D(n9688), .Y(n9716) );
  MUX2X1 U8450 ( .B(n6356), .A(n6060), .S(n5887), .Y(n9718) );
  MUX2X1 U8451 ( .B(n5584), .A(n5448), .S(n5890), .Y(n9719) );
  AOI22X1 U8452 ( .A(n8954), .B(n5584), .C(n5770), .D(n10222), .Y(n9728) );
  MUX2X1 U8453 ( .B(n6359), .A(n6358), .S(n9577), .Y(n9720) );
  MUX2X1 U8454 ( .B(n6358), .A(n6359), .S(n70), .Y(n9721) );
  MUX2X1 U8455 ( .B(n173), .A(n5635), .S(n6245), .Y(n9722) );
  OAI21X1 U8456 ( .A(n6246), .B(n5702), .C(n1939), .Y(n10218) );
  AOI22X1 U8457 ( .A(n5649), .B(n6721), .C(n9767), .D(n4998), .Y(n9726) );
  NAND3X1 U8458 ( .A(n2654), .B(n3308), .C(n3605), .Y(n9729) );
  MUX2X1 U8459 ( .B(n6090), .A(n6067), .S(n6245), .Y(n9732) );
  NAND3X1 U8460 ( .A(n9732), .B(n6070), .C(n9803), .Y(n9733) );
  MUX2X1 U8461 ( .B(n6088), .A(n5375), .S(n6342), .Y(n9736) );
  AOI22X1 U8462 ( .A(n747), .B(n5825), .C(n6049), .D(n9969), .Y(n9734) );
  NAND3X1 U8463 ( .A(n9736), .B(n3310), .C(n3606), .Y(n9741) );
  AOI22X1 U8464 ( .A(n691), .B(n6119), .C(n2280), .D(n5838), .Y(n9739) );
  AOI22X1 U8465 ( .A(n2922), .B(n6086), .C(n426), .D(n5839), .Y(n9737) );
  NAND3X1 U8466 ( .A(n2655), .B(n3311), .C(n3607), .Y(n9740) );
  AOI22X1 U8467 ( .A(n923), .B(n5824), .C(n9500), .D(n6037), .Y(n9744) );
  AOI22X1 U8468 ( .A(n370), .B(n5778), .C(n602), .D(n5823), .Y(n9742) );
  AOI22X1 U8469 ( .A(n3243), .B(n5827), .C(n1743), .D(n5777), .Y(n9747) );
  AOI22X1 U8470 ( .A(n1261), .B(n5785), .C(n1518), .D(n6123), .Y(n9745) );
  NOR3X1 U8471 ( .A(n9748), .B(n4204), .C(n4530), .Y(n9749) );
  NAND3X1 U8472 ( .A(n2748), .B(n3309), .C(n9749), .Y(n9752) );
  AOI22X1 U8473 ( .A(n2965), .B(n6141), .C(n1823), .D(n6149), .Y(n9757) );
  AOI22X1 U8474 ( .A(n1598), .B(n5784), .C(n6315), .D(n10480), .Y(n9756) );
  AOI22X1 U8475 ( .A(n2826), .B(n6110), .C(n2505), .D(n5781), .Y(n9754) );
  NAND3X1 U8476 ( .A(n2656), .B(n5497), .C(n9755), .Y(n9758) );
  AOI22X1 U8477 ( .A(n3790), .B(n5775), .C(n3469), .D(n5774), .Y(n9764) );
  AOI22X1 U8478 ( .A(n1342), .B(n5772), .C(n828), .D(n6145), .Y(n9761) );
  NAND3X1 U8479 ( .A(n2657), .B(n5300), .C(n9762), .Y(n9827) );
  AOI21X1 U8480 ( .A(n6049), .B(n5800), .C(n10024), .Y(n9765) );
  AOI22X1 U8481 ( .A(n8968), .B(n4895), .C(n3565), .D(n6092), .Y(n9779) );
  AOI22X1 U8482 ( .A(n3886), .B(n5828), .C(n3244), .D(n5827), .Y(n9778) );
  AOI21X1 U8483 ( .A(n21), .B(n9614), .C(n10178), .Y(n9766) );
  NAND3X1 U8484 ( .A(n6060), .B(n6247), .C(n7491), .Y(n10372) );
  OAI21X1 U8485 ( .A(n157), .B(n5445), .C(n4859), .Y(n9776) );
  AOI22X1 U8486 ( .A(n6054), .B(n6077), .C(n6354), .D(n6081), .Y(n9768) );
  AOI22X1 U8487 ( .A(n6354), .B(n5769), .C(n9614), .D(n6356), .Y(n9771) );
  AOI22X1 U8488 ( .A(n5757), .B(n9770), .C(n5754), .D(n5131), .Y(n9773) );
  OAI21X1 U8489 ( .A(n161), .B(n5655), .C(n1890), .Y(n9775) );
  AOI22X1 U8490 ( .A(n6342), .B(n6077), .C(n6081), .D(n6026), .Y(n9781) );
  AOI22X1 U8491 ( .A(n6080), .B(n59), .C(n6083), .D(n6032), .Y(n9780) );
  AOI22X1 U8492 ( .A(n6026), .B(n5769), .C(n59), .D(n9614), .Y(n9782) );
  AOI22X1 U8493 ( .A(n6072), .B(n5237), .C(n10030), .D(n5232), .Y(n9790) );
  NAND3X1 U8494 ( .A(n4748), .B(n4789), .C(n3680), .Y(n9787) );
  AOI22X1 U8495 ( .A(n6039), .B(n2781), .C(n3368), .D(n5212), .Y(n9789) );
  OAI21X1 U8496 ( .A(n4759), .B(n5032), .C(n9791), .Y(n9794) );
  AOI22X1 U8497 ( .A(n6060), .B(n9794), .C(n6038), .D(n9793), .Y(n9800) );
  OAI21X1 U8498 ( .A(n6032), .B(n6091), .C(n6089), .Y(n9796) );
  AOI22X1 U8499 ( .A(n5885), .B(n6066), .C(n6247), .D(n9796), .Y(n9798) );
  NOR3X1 U8500 ( .A(n4069), .B(n4278), .C(n4534), .Y(n9819) );
  AOI22X1 U8501 ( .A(n2281), .B(n6104), .C(n2602), .D(n6102), .Y(n9810) );
  AOI22X1 U8502 ( .A(n2923), .B(n6086), .C(n427), .D(n5839), .Y(n9809) );
  AOI22X1 U8503 ( .A(n748), .B(n6137), .C(n6351), .D(n9969), .Y(n9807) );
  MUX2X1 U8504 ( .B(n6091), .A(n6068), .S(n6247), .Y(n9802) );
  NOR3X1 U8505 ( .A(n5728), .B(n9731), .C(n9802), .Y(n9804) );
  MUX2X1 U8506 ( .B(n10522), .A(n9804), .S(n6032), .Y(n9805) );
  AOI21X1 U8507 ( .A(n1085), .B(n5826), .C(n9805), .Y(n9806) );
  NAND3X1 U8508 ( .A(n5372), .B(n5611), .C(n9808), .Y(n9817) );
  AOI22X1 U8509 ( .A(n5961), .B(n10502), .C(n371), .D(n5778), .Y(n9812) );
  AOI22X1 U8510 ( .A(n603), .B(n6135), .C(n692), .D(n5790), .Y(n9811) );
  AOI22X1 U8511 ( .A(n1744), .B(n5777), .C(n1005), .D(n6129), .Y(n9815) );
  AOI22X1 U8512 ( .A(n1519), .B(n5779), .C(n924), .D(n5824), .Y(n9813) );
  NOR3X1 U8513 ( .A(n4073), .B(n4279), .C(n4538), .Y(n9818) );
  AOI22X1 U8514 ( .A(n2993), .B(n6141), .C(n1824), .D(n5783), .Y(n9825) );
  AOI22X1 U8515 ( .A(n1599), .B(n6147), .C(n5276), .D(n10480), .Y(n9824) );
  AOI22X1 U8516 ( .A(n2827), .B(n6110), .C(n2506), .D(n5781), .Y(n9822) );
  NAND3X1 U8517 ( .A(n2658), .B(n3039), .C(n9823), .Y(n9826) );
  AOI22X1 U8518 ( .A(n3791), .B(n6108), .C(n3470), .D(n6106), .Y(n9832) );
  AOI22X1 U8519 ( .A(n1343), .B(n5772), .C(n829), .D(n6145), .Y(n9829) );
  NAND3X1 U8520 ( .A(n2659), .B(n3312), .C(n9830), .Y(n9881) );
  AOI22X1 U8521 ( .A(n5754), .B(n5255), .C(n9774), .D(n5207), .Y(n9837) );
  AOI22X1 U8522 ( .A(n9767), .B(n5125), .C(n8968), .D(n5149), .Y(n9836) );
  AOI22X1 U8523 ( .A(n3566), .B(n5830), .C(n3887), .D(n5828), .Y(n9834) );
  AOI22X1 U8524 ( .A(n3245), .B(n5827), .C(n1745), .D(n5777), .Y(n9833) );
  AOI22X1 U8525 ( .A(n6032), .B(n6077), .C(n6081), .D(n6029), .Y(n9838) );
  AOI21X1 U8526 ( .A(n9614), .B(n6026), .C(n9841), .Y(n9842) );
  AOI22X1 U8527 ( .A(n5628), .B(n5062), .C(n10030), .D(n5134), .Y(n9849) );
  OAI21X1 U8528 ( .A(n9846), .B(n6246), .C(n5696), .Y(n10026) );
  AOI22X1 U8529 ( .A(n5746), .B(n10026), .C(n5212), .D(n4965), .Y(n9848) );
  OAI21X1 U8530 ( .A(n10375), .B(n9784), .C(n6345), .Y(n9850) );
  NAND3X1 U8531 ( .A(n2749), .B(n4859), .C(n9850), .Y(n9904) );
  OAI21X1 U8532 ( .A(n5885), .B(n6091), .C(n6089), .Y(n9854) );
  AOI22X1 U8533 ( .A(n6249), .B(n9854), .C(n4959), .D(n6073), .Y(n9855) );
  NOR3X1 U8534 ( .A(n4074), .B(n4280), .C(n4542), .Y(n9873) );
  AOI22X1 U8535 ( .A(n1006), .B(n5786), .C(n1263), .D(n5785), .Y(n9862) );
  AOI22X1 U8536 ( .A(n1520), .B(n5779), .C(n925), .D(n6133), .Y(n9861) );
  AOI22X1 U8537 ( .A(n5964), .B(n10502), .C(n372), .D(n5778), .Y(n9859) );
  AOI22X1 U8538 ( .A(n604), .B(n5823), .C(n693), .D(n5790), .Y(n9858) );
  NAND3X1 U8539 ( .A(n5472), .B(n5555), .C(n9860), .Y(n9871) );
  MUX2X1 U8540 ( .B(n6090), .A(n6067), .S(n6249), .Y(n9863) );
  MUX2X1 U8541 ( .B(n6088), .A(n5299), .S(n5885), .Y(n9867) );
  AOI22X1 U8542 ( .A(n749), .B(n5825), .C(n6053), .D(n9969), .Y(n9865) );
  AOI22X1 U8543 ( .A(n2282), .B(n5838), .C(n2603), .D(n5831), .Y(n9869) );
  AOI22X1 U8544 ( .A(n2924), .B(n6086), .C(n428), .D(n6131), .Y(n9868) );
  NOR3X1 U8545 ( .A(n4079), .B(n4208), .C(n4616), .Y(n9872) );
  AOI22X1 U8546 ( .A(n2994), .B(n6141), .C(n1825), .D(n5783), .Y(n9879) );
  AOI22X1 U8547 ( .A(n1600), .B(n6147), .C(n27), .D(n10480), .Y(n9878) );
  AOI22X1 U8548 ( .A(n2828), .B(n6110), .C(n2507), .D(n5781), .Y(n9876) );
  NAND3X1 U8549 ( .A(n2660), .B(n3040), .C(n9877), .Y(n9880) );
  AOI22X1 U8550 ( .A(n3792), .B(n6108), .C(n3471), .D(n6106), .Y(n9886) );
  AOI22X1 U8551 ( .A(n1344), .B(n6139), .C(n830), .D(n5771), .Y(n9883) );
  NAND3X1 U8552 ( .A(n2661), .B(n3313), .C(n9884), .Y(n9947) );
  AOI22X1 U8553 ( .A(n9500), .B(n6026), .C(n5966), .D(n10502), .Y(n9888) );
  AOI22X1 U8554 ( .A(n373), .B(n6117), .C(n605), .D(n5823), .Y(n9887) );
  AOI22X1 U8555 ( .A(n1746), .B(n6121), .C(n1007), .D(n6129), .Y(n9891) );
  AOI22X1 U8556 ( .A(n1521), .B(n5779), .C(n926), .D(n5824), .Y(n9889) );
  NAND3X1 U8557 ( .A(n2662), .B(n5484), .C(n3608), .Y(n9892) );
  MUX2X1 U8558 ( .B(n6090), .A(n6067), .S(n6251), .Y(n9894) );
  MUX2X1 U8559 ( .B(n6088), .A(n5338), .S(n6034), .Y(n9898) );
  AOI22X1 U8560 ( .A(n750), .B(n5825), .C(n6354), .D(n9969), .Y(n9896) );
  NAND3X1 U8561 ( .A(n9898), .B(n5391), .C(n5357), .Y(n9903) );
  AOI22X1 U8562 ( .A(n694), .B(n5790), .C(n2283), .D(n6104), .Y(n9901) );
  AOI22X1 U8563 ( .A(n2925), .B(n6086), .C(n429), .D(n6131), .Y(n9899) );
  NAND3X1 U8564 ( .A(n2663), .B(n3314), .C(n3609), .Y(n9902) );
  OAI21X1 U8565 ( .A(n6034), .B(n6091), .C(n6089), .Y(n9905) );
  AOI21X1 U8566 ( .A(n6251), .B(n9905), .C(n4721), .Y(n9927) );
  AOI22X1 U8567 ( .A(n5885), .B(n6077), .C(n6081), .D(n6032), .Y(n9907) );
  AOI22X1 U8568 ( .A(n6080), .B(n6029), .C(n6083), .D(n6034), .Y(n9906) );
  MUX2X1 U8569 ( .B(n10179), .A(n9909), .S(n5890), .Y(n10418) );
  AOI21X1 U8570 ( .A(n6034), .B(n9577), .C(n5811), .Y(n9910) );
  MUX2X1 U8571 ( .B(n4906), .A(n5706), .S(n6245), .Y(n9914) );
  AOI22X1 U8572 ( .A(n10418), .B(n9916), .C(n10425), .D(n4946), .Y(n9926) );
  AOI22X1 U8573 ( .A(n9920), .B(n9917), .C(n9919), .D(n9918), .Y(n9924) );
  AOI22X1 U8574 ( .A(n9922), .B(n5822), .C(n9921), .D(n7147), .Y(n9923) );
  AOI22X1 U8575 ( .A(n8968), .B(n5077), .C(n3567), .D(n5830), .Y(n9929) );
  AOI22X1 U8576 ( .A(n3888), .B(n6096), .C(n3246), .D(n5827), .Y(n9928) );
  AOI22X1 U8577 ( .A(n10034), .B(n10438), .C(n9767), .D(n5128), .Y(n9935) );
  AOI22X1 U8578 ( .A(n5833), .B(n10431), .C(n6791), .D(n4947), .Y(n9933) );
  NOR3X1 U8579 ( .A(n4080), .B(n4281), .C(n4545), .Y(n9937) );
  NAND3X1 U8580 ( .A(n2750), .B(n3315), .C(n9937), .Y(n9940) );
  AOI22X1 U8581 ( .A(n2966), .B(n6141), .C(n1826), .D(n6149), .Y(n9945) );
  AOI22X1 U8582 ( .A(n1601), .B(n6147), .C(n6000), .D(n6112), .Y(n9944) );
  AOI22X1 U8583 ( .A(n2829), .B(n6110), .C(n2508), .D(n6115), .Y(n9942) );
  NAND3X1 U8584 ( .A(n2664), .B(n3041), .C(n9943), .Y(n9946) );
  AOI22X1 U8585 ( .A(n3793), .B(n6108), .C(n3472), .D(n5774), .Y(n9952) );
  AOI22X1 U8586 ( .A(n1345), .B(n5772), .C(n831), .D(n5771), .Y(n9949) );
  NAND3X1 U8587 ( .A(n2665), .B(n3316), .C(n9950), .Y(n10011) );
  AOI22X1 U8588 ( .A(n1522), .B(n5779), .C(n927), .D(n5824), .Y(n9955) );
  AOI22X1 U8589 ( .A(n6296), .B(n10502), .C(n374), .D(n5778), .Y(n9953) );
  NAND3X1 U8590 ( .A(n2666), .B(n3317), .C(n3610), .Y(n9960) );
  AOI22X1 U8591 ( .A(n3889), .B(n5828), .C(n3247), .D(n5827), .Y(n9958) );
  AOI22X1 U8592 ( .A(n1008), .B(n5786), .C(n1265), .D(n5785), .Y(n9956) );
  NAND3X1 U8593 ( .A(n2667), .B(n5609), .C(n3611), .Y(n9959) );
  AOI22X1 U8594 ( .A(n606), .B(n5823), .C(n695), .D(n5790), .Y(n9963) );
  AOI22X1 U8595 ( .A(n2605), .B(n5831), .C(n2926), .D(n5829), .Y(n9961) );
  MUX2X1 U8596 ( .B(n6090), .A(n6067), .S(n6253), .Y(n9964) );
  MUX2X1 U8597 ( .B(n6088), .A(n5673), .S(n6037), .Y(n9967) );
  AOI22X1 U8598 ( .A(n430), .B(n5839), .C(n751), .D(n5825), .Y(n9968) );
  OAI21X1 U8599 ( .A(n6358), .B(n6095), .C(n5527), .Y(n9970) );
  NOR3X1 U8600 ( .A(n4085), .B(n4282), .C(n9970), .Y(n10002) );
  AOI22X1 U8601 ( .A(n9767), .B(n5197), .C(n9930), .D(n4998), .Y(n9975) );
  AOI22X1 U8602 ( .A(n8968), .B(n5584), .C(n3568), .D(n6092), .Y(n9973) );
  NAND3X1 U8603 ( .A(n2668), .B(n3318), .C(n3612), .Y(n9984) );
  AOI22X1 U8604 ( .A(n5770), .B(n5865), .C(n9917), .D(n9977), .Y(n9982) );
  AOI22X1 U8605 ( .A(n5649), .B(n5822), .C(n7147), .D(n9978), .Y(n9980) );
  NAND3X1 U8606 ( .A(n2669), .B(n3319), .C(n3613), .Y(n9983) );
  AOI22X1 U8607 ( .A(n6079), .B(n6032), .C(n6083), .D(n6037), .Y(n9985) );
  AOI22X1 U8608 ( .A(n10026), .B(n5203), .C(n5628), .D(n5137), .Y(n9995) );
  AOI21X1 U8609 ( .A(n5277), .B(n9577), .C(n9988), .Y(n9989) );
  AOI22X1 U8610 ( .A(n9992), .B(n10034), .C(n8954), .D(n10506), .Y(n9993) );
  NAND3X1 U8611 ( .A(n10487), .B(n6247), .C(n10486), .Y(n9999) );
  OAI21X1 U8612 ( .A(n6037), .B(n6091), .C(n6089), .Y(n9997) );
  AOI22X1 U8613 ( .A(n6253), .B(n9997), .C(n10504), .D(n10574), .Y(n9998) );
  NOR3X1 U8614 ( .A(n10000), .B(n4212), .C(n4549), .Y(n10001) );
  NAND3X1 U8615 ( .A(n2751), .B(n10002), .C(n10001), .Y(n10004) );
  AOI22X1 U8616 ( .A(n2967), .B(n6141), .C(n1827), .D(n6149), .Y(n10009) );
  AOI22X1 U8617 ( .A(n1602), .B(n6147), .C(n5283), .D(n6112), .Y(n10008) );
  AOI22X1 U8618 ( .A(n2830), .B(n6110), .C(n2509), .D(n6115), .Y(n10006) );
  NAND3X1 U8619 ( .A(n2670), .B(n5388), .C(n10007), .Y(n10010) );
  AOI22X1 U8620 ( .A(n3794), .B(n6108), .C(n3473), .D(n5774), .Y(n10016) );
  AOI22X1 U8621 ( .A(n1346), .B(n6139), .C(n832), .D(n5771), .Y(n10013) );
  NAND3X1 U8622 ( .A(n2671), .B(n3320), .C(n10014), .Y(n10062) );
  AOI22X1 U8623 ( .A(n9767), .B(n5131), .C(n9930), .D(n4822), .Y(n10022) );
  AOI22X1 U8624 ( .A(n6791), .B(n4895), .C(n8968), .D(n5022), .Y(n10021) );
  AOI22X1 U8625 ( .A(n3569), .B(n5830), .C(n3890), .D(n5828), .Y(n10019) );
  AOI22X1 U8626 ( .A(n3248), .B(n5827), .C(n1748), .D(n6121), .Y(n10018) );
  AOI22X1 U8627 ( .A(n6037), .B(n6077), .C(n6081), .D(n6034), .Y(n10023) );
  AOI22X1 U8628 ( .A(n10026), .B(n5232), .C(n6072), .D(n5171), .Y(n10032) );
  AOI21X1 U8629 ( .A(n6037), .B(n9639), .C(n9770), .Y(n10027) );
  AOI22X1 U8630 ( .A(n10030), .B(n5092), .C(n9770), .D(n9918), .Y(n10031) );
  OAI21X1 U8631 ( .A(n4760), .B(n5032), .C(n10033), .Y(n10035) );
  OAI21X1 U8632 ( .A(n6039), .B(n6091), .C(n6089), .Y(n10036) );
  AOI22X1 U8633 ( .A(n6255), .B(n10036), .C(n10574), .D(n5237), .Y(n10037) );
  NOR3X1 U8634 ( .A(n4089), .B(n4283), .C(n4553), .Y(n10054) );
  AOI22X1 U8635 ( .A(n1009), .B(n5786), .C(n1266), .D(n5785), .Y(n10044) );
  AOI22X1 U8636 ( .A(n1523), .B(n5779), .C(n928), .D(n5824), .Y(n10043) );
  AOI22X1 U8637 ( .A(n9500), .B(n6032), .C(n5970), .D(n10502), .Y(n10041) );
  AOI22X1 U8638 ( .A(n375), .B(n6117), .C(n607), .D(n5823), .Y(n10040) );
  MUX2X1 U8639 ( .B(n6090), .A(n6067), .S(n6255), .Y(n10045) );
  MUX2X1 U8640 ( .B(n6088), .A(n2941), .S(n6039), .Y(n10049) );
  AOI22X1 U8641 ( .A(n431), .B(n5839), .C(n752), .D(n5825), .Y(n10047) );
  AOI22X1 U8642 ( .A(n696), .B(n5790), .C(n2285), .D(n6104), .Y(n10051) );
  AOI22X1 U8643 ( .A(n2606), .B(n5831), .C(n2927), .D(n5829), .Y(n10050) );
  NOR3X1 U8644 ( .A(n4094), .B(n4216), .C(n4617), .Y(n10053) );
  AOI22X1 U8645 ( .A(n2995), .B(n6141), .C(n1828), .D(n5783), .Y(n10060) );
  AOI22X1 U8646 ( .A(n1603), .B(n6147), .C(n6003), .D(n10480), .Y(n10059) );
  AOI22X1 U8647 ( .A(n2831), .B(n6110), .C(n2510), .D(n6115), .Y(n10057) );
  NAND3X1 U8648 ( .A(n131), .B(n3042), .C(n10058), .Y(n10061) );
  AOI22X1 U8649 ( .A(n3795), .B(n6108), .C(n3474), .D(n6106), .Y(n10067) );
  AOI22X1 U8650 ( .A(n1347), .B(n5772), .C(n833), .D(n5771), .Y(n10064) );
  NAND3X1 U8651 ( .A(n5536), .B(n5674), .C(n10065), .Y(n10125) );
  AOI21X1 U8652 ( .A(n6079), .B(n6034), .C(n10068), .Y(n10069) );
  AOI22X1 U8653 ( .A(n59), .B(n10072), .C(n6625), .D(n5000), .Y(n10081) );
  AOI21X1 U8654 ( .A(n6345), .B(n9639), .C(n10073), .Y(n10074) );
  AOI22X1 U8655 ( .A(n10500), .B(n5062), .C(n9689), .D(n4930), .Y(n10080) );
  AOI22X1 U8656 ( .A(n3570), .B(n5830), .C(n3891), .D(n6096), .Y(n10078) );
  AOI22X1 U8657 ( .A(n3249), .B(n5827), .C(n1749), .D(n5777), .Y(n10077) );
  AOI22X1 U8658 ( .A(n5746), .B(n5797), .C(n9767), .D(n5255), .Y(n10084) );
  AOI22X1 U8659 ( .A(n10082), .B(n5134), .C(n9930), .D(n5125), .Y(n10083) );
  OAI21X1 U8660 ( .A(n6042), .B(n6091), .C(n6089), .Y(n10086) );
  OAI21X1 U8661 ( .A(n6359), .B(n5729), .C(n5399), .Y(n10225) );
  AOI21X1 U8662 ( .A(n6257), .B(n10086), .C(n10225), .Y(n10097) );
  OAI21X1 U8663 ( .A(n6352), .B(n5723), .C(n5597), .Y(n10089) );
  AOI21X1 U8664 ( .A(n6046), .B(n10154), .C(n10089), .Y(n10092) );
  AOI22X1 U8665 ( .A(n5793), .B(n6356), .C(n6061), .D(n10216), .Y(n10091) );
  AOI22X1 U8666 ( .A(n6354), .B(n10154), .C(n6054), .D(n10355), .Y(n10090) );
  MUX2X1 U8667 ( .B(n2772), .A(n10386), .S(n6261), .Y(n10094) );
  AOI22X1 U8668 ( .A(n5149), .B(n6073), .C(n10094), .D(n5733), .Y(n10095) );
  NOR3X1 U8669 ( .A(n4099), .B(n4284), .C(n4556), .Y(n10117) );
  AOI22X1 U8670 ( .A(n1010), .B(n6129), .C(n1267), .D(n5785), .Y(n10103) );
  AOI22X1 U8671 ( .A(n1524), .B(n5779), .C(n929), .D(n6133), .Y(n10102) );
  AOI22X1 U8672 ( .A(n6055), .B(n9500), .C(n5973), .D(n10502), .Y(n10100) );
  AOI22X1 U8673 ( .A(n360), .B(n5778), .C(n608), .D(n6135), .Y(n10099) );
  NAND3X1 U8674 ( .A(n5533), .B(n5625), .C(n10101), .Y(n10115) );
  NAND3X1 U8675 ( .A(n10355), .B(n51), .C(n5589), .Y(n10105) );
  MUX2X1 U8676 ( .B(n6091), .A(n6068), .S(n6257), .Y(n10106) );
  AOI21X1 U8677 ( .A(n10208), .B(n10355), .C(n10106), .Y(n10107) );
  NAND3X1 U8678 ( .A(n10556), .B(n6085), .C(n3648), .Y(n10108) );
  MUX2X1 U8679 ( .B(n6088), .A(n2805), .S(n6043), .Y(n10111) );
  AOI22X1 U8680 ( .A(n432), .B(n6131), .C(n753), .D(n5825), .Y(n10109) );
  AOI22X1 U8681 ( .A(n681), .B(n5790), .C(n2286), .D(n6104), .Y(n10113) );
  AOI22X1 U8682 ( .A(n2607), .B(n5831), .C(n2928), .D(n5829), .Y(n10112) );
  NOR3X1 U8683 ( .A(n4104), .B(n4220), .C(n4618), .Y(n10116) );
  AOI22X1 U8684 ( .A(n2996), .B(n6141), .C(n1829), .D(n6149), .Y(n10123) );
  AOI22X1 U8685 ( .A(n1604), .B(n6147), .C(n6328), .D(n6112), .Y(n10122) );
  AOI22X1 U8686 ( .A(n2832), .B(n6110), .C(n2511), .D(n6115), .Y(n10120) );
  NAND3X1 U8687 ( .A(n2672), .B(n5434), .C(n10121), .Y(n10124) );
  AOI22X1 U8688 ( .A(n3796), .B(n6108), .C(n3475), .D(n6106), .Y(n10130) );
  AOI22X1 U8689 ( .A(n1348), .B(n6139), .C(n834), .D(n5771), .Y(n10127) );
  NAND3X1 U8690 ( .A(n2673), .B(n3321), .C(n10128), .Y(n10200) );
  AOI22X1 U8691 ( .A(n930), .B(n5824), .C(n6354), .D(n9500), .Y(n10133) );
  AOI22X1 U8692 ( .A(n361), .B(n6117), .C(n609), .D(n6135), .Y(n10131) );
  NAND3X1 U8693 ( .A(n2674), .B(n3322), .C(n3614), .Y(n10138) );
  AOI22X1 U8694 ( .A(n3250), .B(n5827), .C(n1750), .D(n5777), .Y(n10136) );
  AOI22X1 U8695 ( .A(n1268), .B(n6125), .C(n1525), .D(n6123), .Y(n10134) );
  NAND3X1 U8696 ( .A(n2675), .B(n5545), .C(n5492), .Y(n10137) );
  MUX2X1 U8697 ( .B(n6090), .A(n6067), .S(n6259), .Y(n10139) );
  MUX2X1 U8698 ( .B(n5832), .A(n5477), .S(n5734), .Y(n10143) );
  AOI22X1 U8699 ( .A(n754), .B(n5825), .C(n6094), .D(n6026), .Y(n10141) );
  NAND3X1 U8700 ( .A(n10143), .B(n5694), .C(n5553), .Y(n10148) );
  AOI22X1 U8701 ( .A(n682), .B(n5790), .C(n2287), .D(n6104), .Y(n10146) );
  AOI22X1 U8702 ( .A(n2929), .B(n5829), .C(n433), .D(n6131), .Y(n10144) );
  NAND3X1 U8703 ( .A(n2676), .B(n3323), .C(n3615), .Y(n10147) );
  AOI21X1 U8704 ( .A(n5793), .B(n6351), .C(n10297), .Y(n10150) );
  OAI21X1 U8705 ( .A(n5723), .B(n6353), .C(n1914), .Y(n10165) );
  NAND3X1 U8706 ( .A(n6043), .B(n5819), .C(n10154), .Y(n10151) );
  OAI21X1 U8707 ( .A(n10104), .B(n4807), .C(n1915), .Y(n10152) );
  AOI21X1 U8708 ( .A(n10291), .B(n10165), .C(n10152), .Y(n10160) );
  AOI21X1 U8709 ( .A(n10355), .B(n6355), .C(n2377), .Y(n10157) );
  OAI21X1 U8710 ( .A(n6356), .B(n4806), .C(n4845), .Y(n10155) );
  NAND3X1 U8711 ( .A(n4845), .B(n5723), .C(n3681), .Y(n10158) );
  AOI22X1 U8712 ( .A(n10439), .B(n10290), .C(n10437), .D(n10291), .Y(n10159)
         );
  MUX2X1 U8713 ( .B(n2773), .A(n2785), .S(n6261), .Y(n10161) );
  NOR3X1 U8714 ( .A(n4127), .B(n10161), .C(n10225), .Y(n10174) );
  OAI21X1 U8715 ( .A(n6046), .B(n6091), .C(n6089), .Y(n10163) );
  AOI22X1 U8716 ( .A(n6259), .B(n10163), .C(n5077), .D(n6073), .Y(n10173) );
  OAI21X1 U8717 ( .A(n10164), .B(n10165), .C(n10208), .Y(n10166) );
  OAI21X1 U8718 ( .A(n10168), .B(n5703), .C(n10166), .Y(n10169) );
  AOI21X1 U8719 ( .A(n5836), .B(n5791), .C(n10169), .Y(n10171) );
  AOI22X1 U8720 ( .A(n6721), .B(n10441), .C(n10082), .D(n4906), .Y(n10170) );
  NAND3X1 U8721 ( .A(n10174), .B(n3043), .C(n10172), .Y(n10189) );
  AOI21X1 U8722 ( .A(n6039), .B(n5769), .C(n10175), .Y(n10176) );
  AOI22X1 U8723 ( .A(n10500), .B(n4766), .C(n9689), .D(n5003), .Y(n10181) );
  AOI22X1 U8724 ( .A(n3571), .B(n5830), .C(n3892), .D(n5828), .Y(n10180) );
  AOI22X1 U8725 ( .A(n9930), .B(n5128), .C(n5834), .D(n10431), .Y(n10187) );
  AOI21X1 U8726 ( .A(n6081), .B(n6345), .C(n5713), .Y(n10184) );
  OAI21X1 U8727 ( .A(n6344), .B(n6062), .C(n1916), .Y(n10432) );
  AOI22X1 U8728 ( .A(n6625), .B(n10432), .C(n10375), .D(n10440), .Y(n10185) );
  NOR3X1 U8729 ( .A(n4105), .B(n4289), .C(n4560), .Y(n10190) );
  NAND3X1 U8730 ( .A(n2752), .B(n3324), .C(n10190), .Y(n10193) );
  AOI22X1 U8731 ( .A(n2968), .B(n6141), .C(n1830), .D(n5783), .Y(n10198) );
  AOI22X1 U8732 ( .A(n1605), .B(n6147), .C(n6330), .D(n6112), .Y(n10197) );
  AOI22X1 U8733 ( .A(n2833), .B(n6110), .C(n2512), .D(n6115), .Y(n10195) );
  NAND3X1 U8734 ( .A(n2677), .B(n3044), .C(n10196), .Y(n10199) );
  AOI22X1 U8735 ( .A(n3797), .B(n6108), .C(n3476), .D(n5774), .Y(n10205) );
  AOI22X1 U8736 ( .A(n1349), .B(n6139), .C(n835), .D(n6145), .Y(n10202) );
  NAND3X1 U8737 ( .A(n2678), .B(n3325), .C(n10203), .Y(n10274) );
  AOI22X1 U8738 ( .A(n6054), .B(n5793), .C(n6354), .D(n10216), .Y(n10207) );
  AOI22X1 U8739 ( .A(n6351), .B(n10154), .C(n10355), .D(n21), .Y(n10206) );
  MUX2X1 U8740 ( .B(n6061), .A(n6356), .S(n10355), .Y(n10209) );
  MUX2X1 U8741 ( .B(n6356), .A(n6061), .S(n6257), .Y(n10210) );
  AOI22X1 U8742 ( .A(n5710), .B(n10291), .C(n5818), .D(n6), .Y(n10211) );
  NAND3X1 U8743 ( .A(n2753), .B(n6089), .C(n3616), .Y(n10213) );
  AOI22X1 U8744 ( .A(n2997), .B(n5106), .C(n6261), .D(n3376), .Y(n10221) );
  AOI22X1 U8745 ( .A(n6257), .B(n6348), .C(n6259), .D(n6040), .Y(n10215) );
  AOI22X1 U8746 ( .A(n154), .B(n10356), .C(n10218), .D(n6248), .Y(n10219) );
  OAI21X1 U8747 ( .A(n10224), .B(n8171), .C(n1940), .Y(n10229) );
  NAND3X1 U8748 ( .A(n7491), .B(n5794), .C(n5197), .Y(n10228) );
  NOR3X1 U8749 ( .A(n4106), .B(n10229), .C(n4564), .Y(n10266) );
  AOI22X1 U8750 ( .A(n9689), .B(n4933), .C(n3572), .D(n6092), .Y(n10236) );
  AOI22X1 U8751 ( .A(n3893), .B(n6096), .C(n3251), .D(n5827), .Y(n10235) );
  AOI22X1 U8752 ( .A(n10082), .B(n5050), .C(n7172), .D(n10504), .Y(n10243) );
  AOI22X1 U8753 ( .A(n5886), .B(n6348), .C(shift_amount[3]), .D(n6040), .Y(
        n10237) );
  AOI22X1 U8754 ( .A(n6625), .B(n4767), .C(n10500), .D(n5137), .Y(n10241) );
  NAND3X1 U8755 ( .A(n2679), .B(n3326), .C(n3617), .Y(n10244) );
  MUX2X1 U8756 ( .B(n6090), .A(n6067), .S(n6261), .Y(n10246) );
  MUX2X1 U8757 ( .B(n6088), .A(n5605), .S(n6049), .Y(n10250) );
  AOI22X1 U8758 ( .A(n755), .B(n6137), .C(n6094), .D(n6029), .Y(n10248) );
  NAND3X1 U8759 ( .A(n10250), .B(n3328), .C(n3618), .Y(n10255) );
  AOI22X1 U8760 ( .A(n683), .B(n5790), .C(n2288), .D(n6104), .Y(n10253) );
  AOI22X1 U8761 ( .A(n2930), .B(n5829), .C(n434), .D(n6131), .Y(n10251) );
  NAND3X1 U8762 ( .A(n2680), .B(n3330), .C(n3619), .Y(n10254) );
  AOI22X1 U8763 ( .A(n9500), .B(n6356), .C(n5977), .D(n10502), .Y(n10257) );
  AOI22X1 U8764 ( .A(n362), .B(n5778), .C(n610), .D(n5823), .Y(n10256) );
  AOI22X1 U8765 ( .A(n1751), .B(n5777), .C(n1012), .D(n6129), .Y(n10260) );
  AOI22X1 U8766 ( .A(n1526), .B(n5779), .C(n931), .D(n6133), .Y(n10258) );
  NAND3X1 U8767 ( .A(n2681), .B(n5546), .C(n5693), .Y(n10261) );
  NOR3X1 U8768 ( .A(n10263), .B(n4290), .C(n4567), .Y(n10264) );
  NAND3X1 U8769 ( .A(n10266), .B(n3327), .C(n10264), .Y(n10267) );
  AOI22X1 U8770 ( .A(n2969), .B(n6141), .C(n1831), .D(n5783), .Y(n10272) );
  AOI22X1 U8771 ( .A(n1606), .B(n6147), .C(n6332), .D(n6112), .Y(n10271) );
  AOI22X1 U8772 ( .A(n2834), .B(n5780), .C(n2513), .D(n5781), .Y(n10269) );
  NAND3X1 U8773 ( .A(n2682), .B(n5498), .C(n10270), .Y(n10273) );
  AOI22X1 U8774 ( .A(n3798), .B(n6108), .C(n3477), .D(n6106), .Y(n10279) );
  AOI22X1 U8775 ( .A(n1350), .B(n6139), .C(n836), .D(n5771), .Y(n10276) );
  NAND3X1 U8776 ( .A(n2683), .B(n3331), .C(n10277), .Y(n10341) );
  AOI22X1 U8777 ( .A(n10082), .B(n5092), .C(n9930), .D(n5131), .Y(n10289) );
  AOI22X1 U8778 ( .A(n7172), .B(n5237), .C(n10500), .D(n5171), .Y(n10288) );
  AOI22X1 U8779 ( .A(n9689), .B(n4936), .C(n3573), .D(n6092), .Y(n10286) );
  AOI22X1 U8780 ( .A(n3894), .B(n5828), .C(n3252), .D(n5827), .Y(n10285) );
  OAI21X1 U8781 ( .A(n5513), .B(n5656), .C(n5588), .Y(n10295) );
  NAND3X1 U8782 ( .A(n2754), .B(n4790), .C(n5756), .Y(n10294) );
  AOI22X1 U8783 ( .A(n5765), .B(n10295), .C(n6061), .D(n3378), .Y(n10299) );
  AOI22X1 U8784 ( .A(n5793), .B(n5734), .C(n10216), .D(n6043), .Y(n10296) );
  AOI22X1 U8785 ( .A(n5797), .B(n5232), .C(n10356), .D(n4863), .Y(n10298) );
  OAI21X1 U8786 ( .A(n6351), .B(n6091), .C(n6089), .Y(n10301) );
  AOI21X1 U8787 ( .A(n6263), .B(n10301), .C(n10300), .Y(n10313) );
  NAND3X1 U8788 ( .A(n4746), .B(n10305), .C(n4973), .Y(n10575) );
  AOI22X1 U8789 ( .A(n6354), .B(n5793), .C(n10216), .D(n6356), .Y(n10307) );
  NAND3X1 U8790 ( .A(n2755), .B(n4874), .C(n3620), .Y(n10310) );
  AOI22X1 U8791 ( .A(n6072), .B(n4876), .C(n3370), .D(n5106), .Y(n10311) );
  NOR3X1 U8792 ( .A(n4110), .B(n4291), .C(n4568), .Y(n10333) );
  AOI22X1 U8793 ( .A(n2289), .B(n5838), .C(n2610), .D(n6102), .Y(n10323) );
  AOI22X1 U8794 ( .A(n2931), .B(n5829), .C(n435), .D(n6131), .Y(n10322) );
  AOI22X1 U8795 ( .A(n756), .B(n6137), .C(n9969), .D(n6032), .Y(n10320) );
  MUX2X1 U8796 ( .B(n6091), .A(n6068), .S(n6263), .Y(n10316) );
  MUX2X1 U8797 ( .B(n10522), .A(n5672), .S(n6052), .Y(n10318) );
  AOI21X1 U8798 ( .A(n1093), .B(n6127), .C(n10318), .Y(n10319) );
  NAND3X1 U8799 ( .A(n5415), .B(n5550), .C(n10321), .Y(n10331) );
  AOI22X1 U8800 ( .A(n5980), .B(n10502), .C(n363), .D(n5778), .Y(n10325) );
  AOI22X1 U8801 ( .A(n611), .B(n5823), .C(n684), .D(n5790), .Y(n10324) );
  AOI22X1 U8802 ( .A(n1752), .B(n5777), .C(n1013), .D(n6129), .Y(n10328) );
  AOI22X1 U8803 ( .A(n1527), .B(n6123), .C(n932), .D(n5824), .Y(n10326) );
  NOR3X1 U8804 ( .A(n4115), .B(n4292), .C(n75), .Y(n10332) );
  AOI22X1 U8805 ( .A(n2998), .B(n6142), .C(n1832), .D(n5783), .Y(n10339) );
  AOI22X1 U8806 ( .A(n1607), .B(n6147), .C(n5269), .D(n6112), .Y(n10338) );
  AOI22X1 U8807 ( .A(n2835), .B(n5780), .C(n2514), .D(n5781), .Y(n10336) );
  NAND3X1 U8808 ( .A(n2685), .B(n3045), .C(n10337), .Y(n10340) );
  AOI22X1 U8809 ( .A(n3799), .B(n6108), .C(n3478), .D(n5774), .Y(n10346) );
  AOI22X1 U8810 ( .A(n1351), .B(n5772), .C(n837), .D(n5771), .Y(n10343) );
  NAND3X1 U8811 ( .A(n2686), .B(n3332), .C(n10344), .Y(n10411) );
  AOI22X1 U8812 ( .A(n933), .B(n5824), .C(n5982), .D(n6098), .Y(n10348) );
  AOI22X1 U8813 ( .A(n364), .B(n5778), .C(n612), .D(n6135), .Y(n10347) );
  AOI22X1 U8814 ( .A(n3253), .B(n5827), .C(n1753), .D(n5777), .Y(n10351) );
  AOI22X1 U8815 ( .A(n1271), .B(n6125), .C(n1528), .D(n6123), .Y(n10349) );
  NAND3X1 U8816 ( .A(n2687), .B(n3333), .C(n3621), .Y(n10352) );
  OAI21X1 U8817 ( .A(n5397), .B(n5513), .C(n5732), .Y(n10518) );
  MUX2X1 U8818 ( .B(n6090), .A(n6067), .S(n3), .Y(n10357) );
  NAND3X1 U8819 ( .A(n10449), .B(n10357), .C(n10447), .Y(n10358) );
  MUX2X1 U8820 ( .B(n6088), .A(n2806), .S(n6054), .Y(n10361) );
  AOI22X1 U8821 ( .A(n757), .B(n6137), .C(n6094), .D(n5885), .Y(n10359) );
  NAND3X1 U8822 ( .A(n10361), .B(n3334), .C(n3622), .Y(n10366) );
  AOI22X1 U8823 ( .A(n685), .B(n5790), .C(n2290), .D(n6104), .Y(n10364) );
  AOI22X1 U8824 ( .A(n2932), .B(n5829), .C(n436), .D(n6131), .Y(n10362) );
  NAND3X1 U8825 ( .A(n2688), .B(n3335), .C(n3623), .Y(n10365) );
  AOI21X1 U8826 ( .A(n10154), .B(n10356), .C(n5749), .Y(n10367) );
  OAI21X1 U8827 ( .A(n10370), .B(n5654), .C(n6060), .Y(n10373) );
  OAI21X1 U8828 ( .A(n6359), .B(n5719), .C(n5526), .Y(n10489) );
  AOI21X1 U8829 ( .A(n6351), .B(n5180), .C(n4722), .Y(n10393) );
  AOI21X1 U8830 ( .A(n5793), .B(n10356), .C(n5751), .Y(n10377) );
  AOI21X1 U8831 ( .A(n10216), .B(n10356), .C(n5750), .Y(n10380) );
  AOI22X1 U8832 ( .A(n6048), .B(n5175), .C(n6347), .D(n5220), .Y(n10392) );
  OAI21X1 U8833 ( .A(n6054), .B(n6091), .C(n6089), .Y(n10384) );
  AOI22X1 U8834 ( .A(n6042), .B(n2782), .C(n3), .D(n10384), .Y(n10390) );
  AOI22X1 U8835 ( .A(n5207), .B(n6073), .C(n5106), .D(n4829), .Y(n10389) );
  AOI22X1 U8836 ( .A(n7172), .B(n5062), .C(n10500), .D(n5000), .Y(n10395) );
  AOI22X1 U8837 ( .A(n3574), .B(n6092), .C(n3895), .D(n6096), .Y(n10394) );
  AOI22X1 U8838 ( .A(n5746), .B(n5804), .C(n5797), .D(n5134), .Y(n10399) );
  AOI22X1 U8839 ( .A(n10082), .B(n4930), .C(n9930), .D(n5255), .Y(n10397) );
  NOR3X1 U8840 ( .A(n4116), .B(n4293), .C(n4573), .Y(n10401) );
  NAND3X1 U8841 ( .A(n2756), .B(n3336), .C(n10401), .Y(n10404) );
  AOI22X1 U8842 ( .A(n2971), .B(n6142), .C(n1833), .D(n5783), .Y(n10409) );
  AOI22X1 U8843 ( .A(n1608), .B(n6147), .C(n5286), .D(n6112), .Y(n10408) );
  AOI22X1 U8844 ( .A(n2836), .B(n6110), .C(n2515), .D(n6115), .Y(n10406) );
  NAND3X1 U8845 ( .A(n132), .B(n3046), .C(n10407), .Y(n10410) );
  AOI22X1 U8846 ( .A(n3800), .B(n6108), .C(n3479), .D(n6106), .Y(n10416) );
  AOI22X1 U8847 ( .A(n1352), .B(n6139), .C(n838), .D(n5771), .Y(n10413) );
  AND2X2 U8848 ( .A(n5461), .B(n5462), .Y(n10414) );
  NAND3X1 U8849 ( .A(n2689), .B(n3338), .C(n10414), .Y(n10478) );
  AOI22X1 U8850 ( .A(n6351), .B(n5175), .C(n6049), .D(n5220), .Y(n10422) );
  OAI21X1 U8851 ( .A(n9500), .B(n10417), .C(n6347), .Y(n10421) );
  OAI21X1 U8852 ( .A(n6354), .B(n6091), .C(n6089), .Y(n10419) );
  AOI22X1 U8853 ( .A(n6267), .B(n10419), .C(n5791), .D(n10418), .Y(n10420) );
  NAND3X1 U8854 ( .A(n2690), .B(n10421), .C(n3624), .Y(n10429) );
  NAND3X1 U8855 ( .A(n6042), .B(n10154), .C(n10498), .Y(n10427) );
  AOI22X1 U8856 ( .A(n10424), .B(n10425), .C(n6054), .D(n5180), .Y(n10426) );
  NAND3X1 U8857 ( .A(n10423), .B(n3058), .C(n3625), .Y(n10428) );
  AOI22X1 U8858 ( .A(n7351), .B(n5713), .C(n10082), .D(n5003), .Y(n10435) );
  AOI22X1 U8859 ( .A(n10500), .B(n10432), .C(n3575), .D(n5830), .Y(n10433) );
  NAND3X1 U8860 ( .A(n2691), .B(n3339), .C(n3626), .Y(n10446) );
  AOI22X1 U8861 ( .A(n5794), .B(n10438), .C(n10437), .D(n10436), .Y(n10444) );
  AOI22X1 U8862 ( .A(n5822), .B(n10441), .C(n7147), .D(n10440), .Y(n10442) );
  NAND3X1 U8863 ( .A(n2692), .B(n3340), .C(n3627), .Y(n10445) );
  MUX2X1 U8864 ( .B(n6090), .A(n6067), .S(n6267), .Y(n10448) );
  NAND3X1 U8865 ( .A(n10449), .B(n10448), .C(n10447), .Y(n10450) );
  MUX2X1 U8866 ( .B(n6088), .A(n2807), .S(n6354), .Y(n10453) );
  AOI22X1 U8867 ( .A(n6137), .B(n758), .C(n9969), .D(n6034), .Y(n10451) );
  AOI22X1 U8868 ( .A(n686), .B(n5790), .C(n2291), .D(n6104), .Y(n10456) );
  AOI22X1 U8869 ( .A(n2933), .B(n5829), .C(n437), .D(n6131), .Y(n10454) );
  NAND3X1 U8870 ( .A(n2693), .B(n3342), .C(n3628), .Y(n10457) );
  AOI22X1 U8871 ( .A(n1529), .B(n6123), .C(n934), .D(n6133), .Y(n10461) );
  AOI22X1 U8872 ( .A(n365), .B(n5778), .C(n613), .D(n6135), .Y(n10459) );
  NAND3X1 U8873 ( .A(n133), .B(n3343), .C(n3630), .Y(n10466) );
  AOI22X1 U8874 ( .A(n3896), .B(n5828), .C(n3254), .D(n5827), .Y(n10464) );
  AOI22X1 U8875 ( .A(n1015), .B(n5786), .C(n1272), .D(n5785), .Y(n10462) );
  NOR3X1 U8876 ( .A(n38), .B(n10467), .C(n146), .Y(n10468) );
  NAND3X1 U8877 ( .A(n2757), .B(n3341), .C(n10468), .Y(n10471) );
  AOI22X1 U8878 ( .A(n6142), .B(n139), .C(n1834), .D(n6149), .Y(n10476) );
  AOI22X1 U8879 ( .A(n1609), .B(n6147), .C(n6018), .D(n10480), .Y(n10475) );
  AOI22X1 U8880 ( .A(n2837), .B(n5780), .C(n2516), .D(n5781), .Y(n10473) );
  NAND3X1 U8881 ( .A(n10474), .B(n3048), .C(n134), .Y(n10477) );
  OR2X2 U8882 ( .A(n119), .B(n106), .Y(result[2]) );
  AOI22X1 U8883 ( .A(n6147), .B(n1610), .C(n5783), .D(n1835), .Y(n10553) );
  AOI22X1 U8884 ( .A(n3480), .B(n6106), .C(n3801), .D(n6108), .Y(n10484) );
  AOI22X1 U8885 ( .A(n2196), .B(n6113), .C(n2517), .D(n6115), .Y(n10483) );
  OAI21X1 U8886 ( .A(n5722), .B(n6338), .C(n5315), .Y(n10481) );
  AOI21X1 U8887 ( .A(n3159), .B(n5776), .C(n10481), .Y(n10482) );
  NAND3X1 U8888 ( .A(n2694), .B(n3049), .C(n3649), .Y(n10485) );
  AOI21X1 U8889 ( .A(n1353), .B(n5772), .C(n2354), .Y(n10550) );
  AOI22X1 U8890 ( .A(n759), .B(n5825), .C(n1016), .D(n6129), .Y(n10546) );
  AOI22X1 U8891 ( .A(n9992), .B(n5794), .C(n5429), .D(n6248), .Y(n10515) );
  OAI21X1 U8892 ( .A(n6356), .B(n6091), .C(n6089), .Y(n10490) );
  AOI21X1 U8893 ( .A(n6269), .B(n10490), .C(n10489), .Y(n10493) );
  NAND3X1 U8894 ( .A(n5738), .B(n3059), .C(n3682), .Y(n10494) );
  AOI21X1 U8895 ( .A(n5797), .B(n5050), .C(n2355), .Y(n10514) );
  AOI22X1 U8896 ( .A(n7351), .B(n153), .C(n10208), .D(n10495), .Y(n10496) );
  OAI21X1 U8897 ( .A(n4761), .B(n4791), .C(n1891), .Y(n10512) );
  AOI22X1 U8898 ( .A(n6094), .B(n6038), .C(n21), .D(n9500), .Y(n10501) );
  OAI21X1 U8899 ( .A(n6099), .B(n6309), .C(n1892), .Y(n10503) );
  AOI21X1 U8900 ( .A(n8485), .B(n10504), .C(n10503), .Y(n10510) );
  AOI22X1 U8901 ( .A(n7172), .B(n5137), .C(n10436), .D(n5710), .Y(n10508) );
  NOR3X1 U8902 ( .A(n10512), .B(n4294), .C(n4578), .Y(n10513) );
  NAND3X1 U8903 ( .A(n2696), .B(n3060), .C(n10513), .Y(n10516) );
  AOI21X1 U8904 ( .A(n3255), .B(n5827), .C(n2356), .Y(n10530) );
  MUX2X1 U8905 ( .B(n6091), .A(n6068), .S(n6269), .Y(n10519) );
  NOR3X1 U8906 ( .A(n4847), .B(n10519), .C(n10518), .Y(n10521) );
  MUX2X1 U8907 ( .B(n10522), .A(n10521), .S(n6356), .Y(n10527) );
  AOI22X1 U8908 ( .A(n5804), .B(n5203), .C(n10082), .D(n4933), .Y(n10525) );
  AOI22X1 U8909 ( .A(n6354), .B(n5180), .C(n6351), .D(n5220), .Y(n10523) );
  NAND3X1 U8910 ( .A(n2697), .B(n3346), .C(n3631), .Y(n10526) );
  NAND3X1 U8911 ( .A(n2711), .B(n3347), .C(n3683), .Y(n10531) );
  AOI21X1 U8912 ( .A(n2613), .B(n5831), .C(n2357), .Y(n10534) );
  AOI22X1 U8913 ( .A(n3897), .B(n6096), .C(n3576), .D(n6092), .Y(n10533) );
  NAND3X1 U8914 ( .A(n2712), .B(n3050), .C(n3684), .Y(n10535) );
  AOI21X1 U8915 ( .A(n366), .B(n5778), .C(n2358), .Y(n10538) );
  NAND3X1 U8916 ( .A(n2713), .B(n3348), .C(n3685), .Y(n10539) );
  AOI21X1 U8917 ( .A(n1530), .B(n6123), .C(n123), .Y(n10542) );
  AOI22X1 U8918 ( .A(n438), .B(n5839), .C(n5785), .D(n1273), .Y(n10540) );
  NAND3X1 U8919 ( .A(n135), .B(n3349), .C(n3632), .Y(n10543) );
  NAND3X1 U8920 ( .A(n2695), .B(n3344), .C(n10544), .Y(n10547) );
  NAND3X1 U8921 ( .A(n136), .B(n2710), .C(n3686), .Y(n10551) );
  AOI21X1 U8922 ( .A(n10292), .B(n5794), .C(n10554), .Y(n10560) );
  MUX2X1 U8923 ( .B(n6090), .A(n6067), .S(n6271), .Y(n10559) );
  NOR3X1 U8924 ( .A(n5265), .B(n4848), .C(n5263), .Y(n10558) );
  NAND3X1 U8925 ( .A(n2714), .B(n10559), .C(n10558), .Y(n10561) );
  MUX2X1 U8926 ( .B(n5832), .A(n2936), .S(n6061), .Y(n10582) );
  AOI22X1 U8927 ( .A(n5804), .B(n5232), .C(n5797), .D(n5092), .Y(n10562) );
  OAI21X1 U8928 ( .A(n168), .B(n6358), .C(n1893), .Y(n10580) );
  OAI21X1 U8929 ( .A(n166), .B(n6355), .C(n1941), .Y(n10579) );
  OAI21X1 U8930 ( .A(n6061), .B(n6091), .C(n6089), .Y(n10568) );
  AOI22X1 U8931 ( .A(n6094), .B(n6039), .C(n3577), .D(n5830), .Y(n10566) );
  AOI21X1 U8932 ( .A(n6271), .B(n10568), .C(n5669), .Y(n10572) );
  AOI22X1 U8933 ( .A(n6351), .B(n9500), .C(n5988), .D(n6098), .Y(n10571) );
  AOI22X1 U8934 ( .A(n8485), .B(n5237), .C(n7172), .D(n5171), .Y(n10570) );
  NAND3X1 U8935 ( .A(n2715), .B(n3051), .C(n3633), .Y(n10573) );
  AOI21X1 U8936 ( .A(n4876), .B(n10574), .C(n2359), .Y(n10578) );
  AOI22X1 U8937 ( .A(n3256), .B(n6100), .C(n10082), .D(n4936), .Y(n10576) );
  NOR3X1 U8938 ( .A(n10580), .B(n10579), .C(n4582), .Y(n10581) );
  NAND3X1 U8939 ( .A(n2758), .B(n10582), .C(n10581), .Y(n10584) );
  AOI21X1 U8940 ( .A(n2614), .B(n5831), .C(n2360), .Y(n10593) );
  AOI22X1 U8941 ( .A(n3802), .B(n5775), .C(n3481), .D(n5774), .Y(n10586) );
  AOI22X1 U8942 ( .A(n5272), .B(n10480), .C(n2839), .D(n5780), .Y(n10588) );
  AOI22X1 U8943 ( .A(n2518), .B(n5781), .C(n2197), .D(n6113), .Y(n10587) );
  NAND3X1 U8944 ( .A(n2716), .B(n3350), .C(n3687), .Y(n10594) );
  AOI21X1 U8945 ( .A(n367), .B(n5778), .C(n2361), .Y(n10597) );
  NAND3X1 U8946 ( .A(n2717), .B(n3351), .C(n3688), .Y(n10598) );
  AOI22X1 U8947 ( .A(n5786), .B(n1017), .C(n6127), .D(n1097), .Y(n10599) );
  NAND3X1 U8948 ( .A(n10601), .B(n141), .C(n144), .Y(n10602) );
  AOI22X1 U8949 ( .A(n6137), .B(n760), .C(n5823), .D(n615), .Y(n10603) );
  AOI22X1 U8950 ( .A(n6141), .B(n10605), .C(n1354), .D(n6139), .Y(n10607) );
  AOI22X1 U8951 ( .A(n1836), .B(n5783), .C(n1611), .D(n6147), .Y(n10609) );
endmodule


module gold_processor ( clk, reset, pc, instruction, memAddr, memEn, memWrEn, 
        dataIn, dataOut );
  output [0:31] pc;
  input [0:31] instruction;
  output [0:31] memAddr;
  input [0:63] dataIn;
  output [0:63] dataOut;
  input clk, reset;
  output memEn, memWrEn;
  wire   n3315, n3316, n3317, WB_reg_write_load, ID_flush_ff, WB_reg_write,
         WB_is_load, WB_is_mul32, PREVIOUS_STALL, PREVIOUS_2_STALL,
         EX_reg_write, EX_is_load, EX_is_mul32, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n291, n299, n1178, n1180, n1181, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1312, n1313, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2573, n2575, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314;
  wire   [0:4] ID_rf_rd1_addr;
  wire   [0:4] WB_dest_reg;
  wire   [0:63] WB_data;
  wire   [0:63] ID_oprB;
  wire   [0:2] WB_PPP;
  wire   [0:63] EX_alu_A;
  wire   [0:63] EX_alu_B;
  wire   [0:5] EX_alu_func;
  wire   [0:4] EX_shift_amt;
  wire   [0:1] EX_WW;
  wire   [0:63] EX_alu_result;
  wire   [0:63] WB_mult32_result;
  wire   [0:15] ID_instruction;
  wire   [0:63] EX_oprA;
  wire   [0:63] EX_oprB;
  wire   [0:63] WB_alu_result;
  wire   [0:4] EX_regA;
  wire   [0:4] EX_regB;
  wire   [0:2] EX_PPP;
  wire   [0:4] EX_dest_reg;
  assign memAddr[15] = 1'b0;
  assign memAddr[14] = 1'b0;
  assign memAddr[13] = 1'b0;
  assign memAddr[12] = 1'b0;
  assign memAddr[11] = 1'b0;
  assign memAddr[10] = 1'b0;
  assign memAddr[9] = 1'b0;
  assign memAddr[8] = 1'b0;
  assign memAddr[7] = 1'b0;
  assign memAddr[6] = 1'b0;
  assign memAddr[5] = 1'b0;
  assign memAddr[4] = 1'b0;
  assign memAddr[3] = 1'b0;
  assign memAddr[2] = 1'b0;
  assign memAddr[1] = 1'b0;
  assign memAddr[0] = 1'b0;

  DFFPOSX1 WB_is_mul32_reg ( .D(n2448), .CLK(clk), .Q(WB_is_mul32) );
  DFFPOSX1 WB_alu_result_reg_63_ ( .D(n224), .CLK(clk), .Q(WB_alu_result[63])
         );
  DFFPOSX1 WB_alu_result_reg_62_ ( .D(n225), .CLK(clk), .Q(WB_alu_result[62])
         );
  DFFPOSX1 WB_alu_result_reg_61_ ( .D(n226), .CLK(clk), .Q(WB_alu_result[61])
         );
  DFFPOSX1 WB_alu_result_reg_60_ ( .D(n227), .CLK(clk), .Q(WB_alu_result[60])
         );
  DFFPOSX1 WB_alu_result_reg_59_ ( .D(n228), .CLK(clk), .Q(WB_alu_result[59])
         );
  DFFPOSX1 WB_alu_result_reg_58_ ( .D(n229), .CLK(clk), .Q(WB_alu_result[58])
         );
  DFFPOSX1 WB_alu_result_reg_57_ ( .D(n230), .CLK(clk), .Q(WB_alu_result[57])
         );
  DFFPOSX1 WB_alu_result_reg_56_ ( .D(n231), .CLK(clk), .Q(WB_alu_result[56])
         );
  DFFPOSX1 WB_alu_result_reg_55_ ( .D(n232), .CLK(clk), .Q(WB_alu_result[55])
         );
  DFFPOSX1 WB_alu_result_reg_54_ ( .D(n233), .CLK(clk), .Q(WB_alu_result[54])
         );
  DFFPOSX1 WB_alu_result_reg_53_ ( .D(n234), .CLK(clk), .Q(WB_alu_result[53])
         );
  DFFPOSX1 WB_alu_result_reg_52_ ( .D(n235), .CLK(clk), .Q(WB_alu_result[52])
         );
  DFFPOSX1 WB_alu_result_reg_51_ ( .D(n236), .CLK(clk), .Q(WB_alu_result[51])
         );
  DFFPOSX1 WB_alu_result_reg_50_ ( .D(n237), .CLK(clk), .Q(WB_alu_result[50])
         );
  DFFPOSX1 WB_alu_result_reg_49_ ( .D(n238), .CLK(clk), .Q(WB_alu_result[49])
         );
  DFFPOSX1 WB_alu_result_reg_48_ ( .D(n239), .CLK(clk), .Q(WB_alu_result[48])
         );
  DFFPOSX1 WB_alu_result_reg_47_ ( .D(n240), .CLK(clk), .Q(WB_alu_result[47])
         );
  DFFPOSX1 WB_alu_result_reg_46_ ( .D(n241), .CLK(clk), .Q(WB_alu_result[46])
         );
  DFFPOSX1 WB_alu_result_reg_45_ ( .D(n242), .CLK(clk), .Q(WB_alu_result[45])
         );
  DFFPOSX1 WB_alu_result_reg_44_ ( .D(n243), .CLK(clk), .Q(WB_alu_result[44])
         );
  DFFPOSX1 WB_alu_result_reg_43_ ( .D(n244), .CLK(clk), .Q(WB_alu_result[43])
         );
  DFFPOSX1 WB_alu_result_reg_42_ ( .D(n245), .CLK(clk), .Q(WB_alu_result[42])
         );
  DFFPOSX1 WB_alu_result_reg_41_ ( .D(n246), .CLK(clk), .Q(WB_alu_result[41])
         );
  DFFPOSX1 WB_alu_result_reg_40_ ( .D(n247), .CLK(clk), .Q(WB_alu_result[40])
         );
  DFFPOSX1 WB_alu_result_reg_39_ ( .D(n248), .CLK(clk), .Q(WB_alu_result[39])
         );
  DFFPOSX1 WB_alu_result_reg_38_ ( .D(n249), .CLK(clk), .Q(WB_alu_result[38])
         );
  DFFPOSX1 WB_alu_result_reg_37_ ( .D(n250), .CLK(clk), .Q(WB_alu_result[37])
         );
  DFFPOSX1 WB_alu_result_reg_36_ ( .D(n251), .CLK(clk), .Q(WB_alu_result[36])
         );
  DFFPOSX1 WB_alu_result_reg_35_ ( .D(n252), .CLK(clk), .Q(WB_alu_result[35])
         );
  DFFPOSX1 WB_alu_result_reg_34_ ( .D(n253), .CLK(clk), .Q(WB_alu_result[34])
         );
  DFFPOSX1 WB_alu_result_reg_33_ ( .D(n254), .CLK(clk), .Q(WB_alu_result[33])
         );
  DFFPOSX1 WB_alu_result_reg_32_ ( .D(n255), .CLK(clk), .Q(WB_alu_result[32])
         );
  DFFPOSX1 WB_alu_result_reg_31_ ( .D(n256), .CLK(clk), .Q(WB_alu_result[31])
         );
  DFFPOSX1 WB_alu_result_reg_30_ ( .D(n257), .CLK(clk), .Q(WB_alu_result[30])
         );
  DFFPOSX1 WB_alu_result_reg_29_ ( .D(n258), .CLK(clk), .Q(WB_alu_result[29])
         );
  DFFPOSX1 WB_alu_result_reg_28_ ( .D(n259), .CLK(clk), .Q(WB_alu_result[28])
         );
  DFFPOSX1 WB_alu_result_reg_27_ ( .D(n260), .CLK(clk), .Q(WB_alu_result[27])
         );
  DFFPOSX1 WB_alu_result_reg_26_ ( .D(n261), .CLK(clk), .Q(WB_alu_result[26])
         );
  DFFPOSX1 WB_alu_result_reg_25_ ( .D(n262), .CLK(clk), .Q(WB_alu_result[25])
         );
  DFFPOSX1 WB_alu_result_reg_24_ ( .D(n263), .CLK(clk), .Q(WB_alu_result[24])
         );
  DFFPOSX1 WB_alu_result_reg_23_ ( .D(n264), .CLK(clk), .Q(WB_alu_result[23])
         );
  DFFPOSX1 WB_alu_result_reg_22_ ( .D(n265), .CLK(clk), .Q(WB_alu_result[22])
         );
  DFFPOSX1 WB_alu_result_reg_21_ ( .D(n266), .CLK(clk), .Q(WB_alu_result[21])
         );
  DFFPOSX1 WB_alu_result_reg_20_ ( .D(n267), .CLK(clk), .Q(WB_alu_result[20])
         );
  DFFPOSX1 WB_alu_result_reg_19_ ( .D(n268), .CLK(clk), .Q(WB_alu_result[19])
         );
  DFFPOSX1 WB_alu_result_reg_18_ ( .D(n269), .CLK(clk), .Q(WB_alu_result[18])
         );
  DFFPOSX1 WB_alu_result_reg_17_ ( .D(n270), .CLK(clk), .Q(WB_alu_result[17])
         );
  DFFPOSX1 WB_alu_result_reg_16_ ( .D(n271), .CLK(clk), .Q(WB_alu_result[16])
         );
  DFFPOSX1 WB_alu_result_reg_15_ ( .D(n272), .CLK(clk), .Q(WB_alu_result[15])
         );
  DFFPOSX1 WB_alu_result_reg_14_ ( .D(n273), .CLK(clk), .Q(WB_alu_result[14])
         );
  DFFPOSX1 WB_alu_result_reg_13_ ( .D(n274), .CLK(clk), .Q(WB_alu_result[13])
         );
  DFFPOSX1 WB_alu_result_reg_12_ ( .D(n275), .CLK(clk), .Q(WB_alu_result[12])
         );
  DFFPOSX1 WB_alu_result_reg_11_ ( .D(n276), .CLK(clk), .Q(WB_alu_result[11])
         );
  DFFPOSX1 WB_alu_result_reg_10_ ( .D(n277), .CLK(clk), .Q(WB_alu_result[10])
         );
  DFFPOSX1 WB_alu_result_reg_9_ ( .D(n278), .CLK(clk), .Q(WB_alu_result[9]) );
  DFFPOSX1 WB_alu_result_reg_8_ ( .D(n279), .CLK(clk), .Q(WB_alu_result[8]) );
  DFFPOSX1 WB_alu_result_reg_7_ ( .D(n280), .CLK(clk), .Q(WB_alu_result[7]) );
  DFFPOSX1 WB_alu_result_reg_6_ ( .D(n281), .CLK(clk), .Q(WB_alu_result[6]) );
  DFFPOSX1 WB_alu_result_reg_5_ ( .D(n282), .CLK(clk), .Q(WB_alu_result[5]) );
  DFFPOSX1 WB_alu_result_reg_4_ ( .D(n283), .CLK(clk), .Q(WB_alu_result[4]) );
  DFFPOSX1 WB_alu_result_reg_3_ ( .D(n284), .CLK(clk), .Q(WB_alu_result[3]) );
  DFFPOSX1 WB_alu_result_reg_2_ ( .D(n285), .CLK(clk), .Q(WB_alu_result[2]) );
  DFFPOSX1 WB_alu_result_reg_1_ ( .D(n286), .CLK(clk), .Q(WB_alu_result[1]) );
  DFFPOSX1 WB_alu_result_reg_0_ ( .D(n287), .CLK(clk), .Q(WB_alu_result[0]) );
  DFFPOSX1 ID_flush_ff_reg ( .D(n1997), .CLK(clk), .Q(ID_flush_ff) );
  DFFPOSX1 ID_instruction_reg_0_ ( .D(n1996), .CLK(clk), .Q(ID_instruction[0])
         );
  DFFPOSX1 ID_instruction_reg_1_ ( .D(n2321), .CLK(clk), .Q(ID_instruction[1])
         );
  DFFPOSX1 ID_instruction_reg_3_ ( .D(n2358), .CLK(clk), .Q(ID_instruction[3])
         );
  DFFPOSX1 EX_reg_write_reg ( .D(n1913), .CLK(clk), .Q(EX_reg_write) );
  DFFPOSX1 WB_reg_write_reg ( .D(n2449), .CLK(clk), .Q(WB_reg_write) );
  DFFPOSX1 EX_oprB_reg_61_ ( .D(n1912), .CLK(clk), .Q(EX_oprB[61]) );
  DFFPOSX1 EX_oprB_reg_60_ ( .D(n1911), .CLK(clk), .Q(EX_oprB[60]) );
  DFFPOSX1 EX_oprB_reg_59_ ( .D(n1910), .CLK(clk), .Q(EX_oprB[59]) );
  DFFPOSX1 EX_oprB_reg_58_ ( .D(n1909), .CLK(clk), .Q(EX_oprB[58]) );
  DFFPOSX1 EX_oprB_reg_57_ ( .D(n1908), .CLK(clk), .Q(EX_oprB[57]) );
  DFFPOSX1 EX_oprB_reg_56_ ( .D(n1907), .CLK(clk), .Q(EX_oprB[56]) );
  DFFPOSX1 EX_oprB_reg_55_ ( .D(n1906), .CLK(clk), .Q(EX_oprB[55]) );
  DFFPOSX1 EX_oprB_reg_54_ ( .D(n1905), .CLK(clk), .Q(EX_oprB[54]) );
  DFFPOSX1 EX_oprB_reg_53_ ( .D(n1904), .CLK(clk), .Q(EX_oprB[53]) );
  DFFPOSX1 EX_oprB_reg_52_ ( .D(n1903), .CLK(clk), .Q(EX_oprB[52]) );
  DFFPOSX1 EX_oprB_reg_51_ ( .D(n1902), .CLK(clk), .Q(EX_oprB[51]) );
  DFFPOSX1 EX_oprB_reg_50_ ( .D(n1901), .CLK(clk), .Q(EX_oprB[50]) );
  DFFPOSX1 EX_oprB_reg_49_ ( .D(n1900), .CLK(clk), .Q(EX_oprB[49]) );
  DFFPOSX1 EX_oprB_reg_48_ ( .D(n1899), .CLK(clk), .Q(EX_oprB[48]) );
  DFFPOSX1 EX_oprB_reg_47_ ( .D(n1898), .CLK(clk), .Q(EX_oprB[47]) );
  DFFPOSX1 EX_oprB_reg_46_ ( .D(n1897), .CLK(clk), .Q(EX_oprB[46]) );
  DFFPOSX1 EX_oprB_reg_45_ ( .D(n1896), .CLK(clk), .Q(EX_oprB[45]) );
  DFFPOSX1 EX_oprB_reg_44_ ( .D(n1895), .CLK(clk), .Q(EX_oprB[44]) );
  DFFPOSX1 EX_oprB_reg_43_ ( .D(n1894), .CLK(clk), .Q(EX_oprB[43]) );
  DFFPOSX1 EX_oprB_reg_42_ ( .D(n1893), .CLK(clk), .Q(EX_oprB[42]) );
  DFFPOSX1 EX_oprB_reg_41_ ( .D(n1892), .CLK(clk), .Q(EX_oprB[41]) );
  DFFPOSX1 EX_oprB_reg_40_ ( .D(n1891), .CLK(clk), .Q(EX_oprB[40]) );
  DFFPOSX1 EX_oprB_reg_39_ ( .D(n1890), .CLK(clk), .Q(EX_oprB[39]) );
  DFFPOSX1 EX_oprB_reg_38_ ( .D(n1889), .CLK(clk), .Q(EX_oprB[38]) );
  DFFPOSX1 EX_oprB_reg_37_ ( .D(n1888), .CLK(clk), .Q(EX_oprB[37]) );
  DFFPOSX1 EX_oprB_reg_36_ ( .D(n1887), .CLK(clk), .Q(EX_oprB[36]) );
  DFFPOSX1 EX_oprB_reg_35_ ( .D(n1886), .CLK(clk), .Q(EX_oprB[35]) );
  DFFPOSX1 EX_oprB_reg_34_ ( .D(n1885), .CLK(clk), .Q(EX_oprB[34]) );
  DFFPOSX1 EX_oprB_reg_33_ ( .D(n1884), .CLK(clk), .Q(EX_oprB[33]) );
  DFFPOSX1 EX_oprB_reg_32_ ( .D(n1883), .CLK(clk), .Q(EX_oprB[32]) );
  DFFPOSX1 EX_oprB_reg_31_ ( .D(n1882), .CLK(clk), .Q(EX_oprB[31]) );
  DFFPOSX1 EX_oprB_reg_30_ ( .D(n1881), .CLK(clk), .Q(EX_oprB[30]) );
  DFFPOSX1 EX_oprB_reg_29_ ( .D(n1880), .CLK(clk), .Q(EX_oprB[29]) );
  DFFPOSX1 EX_oprB_reg_28_ ( .D(n1879), .CLK(clk), .Q(EX_oprB[28]) );
  DFFPOSX1 EX_oprB_reg_27_ ( .D(n1878), .CLK(clk), .Q(EX_oprB[27]) );
  DFFPOSX1 EX_oprB_reg_26_ ( .D(n1877), .CLK(clk), .Q(EX_oprB[26]) );
  DFFPOSX1 EX_oprB_reg_25_ ( .D(n1876), .CLK(clk), .Q(EX_oprB[25]) );
  DFFPOSX1 EX_oprB_reg_24_ ( .D(n1875), .CLK(clk), .Q(EX_oprB[24]) );
  DFFPOSX1 EX_oprB_reg_23_ ( .D(n1874), .CLK(clk), .Q(EX_oprB[23]) );
  DFFPOSX1 EX_oprB_reg_22_ ( .D(n1873), .CLK(clk), .Q(EX_oprB[22]) );
  DFFPOSX1 EX_oprB_reg_21_ ( .D(n1872), .CLK(clk), .Q(EX_oprB[21]) );
  DFFPOSX1 EX_oprB_reg_20_ ( .D(n1871), .CLK(clk), .Q(EX_oprB[20]) );
  DFFPOSX1 EX_oprB_reg_19_ ( .D(n1870), .CLK(clk), .Q(EX_oprB[19]) );
  DFFPOSX1 EX_oprB_reg_18_ ( .D(n1869), .CLK(clk), .Q(EX_oprB[18]) );
  DFFPOSX1 EX_oprB_reg_17_ ( .D(n1868), .CLK(clk), .Q(EX_oprB[17]) );
  DFFPOSX1 EX_oprB_reg_16_ ( .D(n1867), .CLK(clk), .Q(EX_oprB[16]) );
  DFFPOSX1 EX_oprB_reg_15_ ( .D(n1866), .CLK(clk), .Q(EX_oprB[15]) );
  DFFPOSX1 EX_oprB_reg_14_ ( .D(n1865), .CLK(clk), .Q(EX_oprB[14]) );
  DFFPOSX1 EX_oprB_reg_13_ ( .D(n1864), .CLK(clk), .Q(EX_oprB[13]) );
  DFFPOSX1 EX_oprB_reg_12_ ( .D(n1863), .CLK(clk), .Q(EX_oprB[12]) );
  DFFPOSX1 EX_oprB_reg_11_ ( .D(n1862), .CLK(clk), .Q(EX_oprB[11]) );
  DFFPOSX1 EX_oprB_reg_10_ ( .D(n1861), .CLK(clk), .Q(EX_oprB[10]) );
  DFFPOSX1 EX_oprB_reg_9_ ( .D(n1860), .CLK(clk), .Q(EX_oprB[9]) );
  DFFPOSX1 EX_oprB_reg_8_ ( .D(n1859), .CLK(clk), .Q(EX_oprB[8]) );
  DFFPOSX1 EX_oprB_reg_7_ ( .D(n1858), .CLK(clk), .Q(EX_oprB[7]) );
  DFFPOSX1 EX_oprB_reg_6_ ( .D(n1857), .CLK(clk), .Q(EX_oprB[6]) );
  DFFPOSX1 EX_oprB_reg_5_ ( .D(n1856), .CLK(clk), .Q(EX_oprB[5]) );
  DFFPOSX1 EX_oprB_reg_4_ ( .D(n1855), .CLK(clk), .Q(EX_oprB[4]) );
  DFFPOSX1 EX_oprB_reg_3_ ( .D(n1854), .CLK(clk), .Q(EX_oprB[3]) );
  DFFPOSX1 EX_oprB_reg_2_ ( .D(n1853), .CLK(clk), .Q(EX_oprB[2]) );
  DFFPOSX1 EX_oprB_reg_1_ ( .D(n1852), .CLK(clk), .Q(EX_oprB[1]) );
  DFFPOSX1 EX_oprB_reg_0_ ( .D(n1851), .CLK(clk), .Q(EX_oprB[0]) );
  DFFPOSX1 ID_instruction_reg_31_ ( .D(n1850), .CLK(clk), .Q(memAddr[31]) );
  DFFPOSX1 ID_instruction_reg_30_ ( .D(n1849), .CLK(clk), .Q(memAddr[30]) );
  DFFPOSX1 ID_instruction_reg_29_ ( .D(n1848), .CLK(clk), .Q(memAddr[29]) );
  DFFPOSX1 ID_instruction_reg_28_ ( .D(n1847), .CLK(clk), .Q(memAddr[28]) );
  DFFPOSX1 ID_instruction_reg_27_ ( .D(n1846), .CLK(clk), .Q(memAddr[27]) );
  DFFPOSX1 ID_instruction_reg_26_ ( .D(n1845), .CLK(clk), .Q(memAddr[26]) );
  DFFPOSX1 ID_instruction_reg_25_ ( .D(n1838), .CLK(clk), .Q(memAddr[25]) );
  DFFPOSX1 ID_instruction_reg_24_ ( .D(n1837), .CLK(clk), .Q(memAddr[24]) );
  DFFPOSX1 ID_instruction_reg_23_ ( .D(n1834), .CLK(clk), .Q(memAddr[23]) );
  DFFPOSX1 ID_instruction_reg_22_ ( .D(n1833), .CLK(clk), .Q(memAddr[22]) );
  DFFPOSX1 ID_instruction_reg_21_ ( .D(n1832), .CLK(clk), .Q(memAddr[21]) );
  DFFPOSX1 ID_instruction_reg_20_ ( .D(n1828), .CLK(clk), .Q(n3317) );
  DFFPOSX1 EX_regB_reg_4_ ( .D(n1827), .CLK(clk), .Q(EX_regB[4]) );
  DFFPOSX1 ID_instruction_reg_19_ ( .D(n1826), .CLK(clk), .Q(n3316) );
  DFFPOSX1 EX_regB_reg_3_ ( .D(n1825), .CLK(clk), .Q(EX_regB[3]) );
  DFFPOSX1 ID_instruction_reg_18_ ( .D(n1824), .CLK(clk), .Q(n3315) );
  DFFPOSX1 EX_regB_reg_2_ ( .D(n1823), .CLK(clk), .Q(EX_regB[2]) );
  DFFPOSX1 ID_instruction_reg_17_ ( .D(n1822), .CLK(clk), .Q(memAddr[17]) );
  DFFPOSX1 EX_regB_reg_1_ ( .D(n1821), .CLK(clk), .Q(EX_regB[1]) );
  DFFPOSX1 ID_instruction_reg_16_ ( .D(n1820), .CLK(clk), .Q(memAddr[16]) );
  DFFPOSX1 EX_regB_reg_0_ ( .D(n1819), .CLK(clk), .Q(EX_regB[0]) );
  DFFPOSX1 ID_instruction_reg_15_ ( .D(n1813), .CLK(clk), .Q(
        ID_instruction[15]) );
  DFFPOSX1 EX_regA_reg_4_ ( .D(n1812), .CLK(clk), .Q(EX_regA[4]) );
  DFFPOSX1 ID_instruction_reg_14_ ( .D(n1811), .CLK(clk), .Q(
        ID_instruction[14]) );
  DFFPOSX1 EX_regA_reg_3_ ( .D(n1810), .CLK(clk), .Q(EX_regA[3]) );
  DFFPOSX1 ID_instruction_reg_13_ ( .D(n1809), .CLK(clk), .Q(
        ID_instruction[13]) );
  DFFPOSX1 EX_regA_reg_2_ ( .D(n1808), .CLK(clk), .Q(EX_regA[2]) );
  DFFPOSX1 ID_instruction_reg_12_ ( .D(n1807), .CLK(clk), .Q(
        ID_instruction[12]) );
  DFFPOSX1 EX_regA_reg_1_ ( .D(n1806), .CLK(clk), .Q(EX_regA[1]) );
  DFFPOSX1 ID_instruction_reg_11_ ( .D(n1805), .CLK(clk), .Q(
        ID_instruction[11]) );
  DFFPOSX1 EX_regA_reg_0_ ( .D(n1804), .CLK(clk), .Q(EX_regA[0]) );
  DFFPOSX1 ID_instruction_reg_10_ ( .D(n1803), .CLK(clk), .Q(
        ID_instruction[10]) );
  DFFPOSX1 ID_instruction_reg_9_ ( .D(n1802), .CLK(clk), .Q(ID_instruction[9])
         );
  DFFPOSX1 ID_instruction_reg_8_ ( .D(n1801), .CLK(clk), .Q(ID_instruction[8])
         );
  DFFPOSX1 ID_instruction_reg_7_ ( .D(n1800), .CLK(clk), .Q(ID_instruction[7])
         );
  DFFPOSX1 ID_instruction_reg_6_ ( .D(n1799), .CLK(clk), .Q(ID_instruction[6])
         );
  DFFPOSX1 ID_instruction_reg_5_ ( .D(n1793), .CLK(clk), .Q(ID_instruction[5])
         );
  DFFPOSX1 ID_instruction_reg_4_ ( .D(n1792), .CLK(clk), .Q(ID_instruction[4])
         );
  DFFPOSX1 EX_oprB_reg_63_ ( .D(n1785), .CLK(clk), .Q(EX_oprB[63]) );
  DFFPOSX1 EX_oprB_reg_62_ ( .D(n1784), .CLK(clk), .Q(EX_oprB[62]) );
  DFFPOSX1 EX_oprA_reg_1_ ( .D(n1721), .CLK(clk), .Q(EX_oprA[1]) );
  DFFPOSX1 EX_oprA_reg_2_ ( .D(n1722), .CLK(clk), .Q(EX_oprA[2]) );
  DFFPOSX1 EX_oprA_reg_3_ ( .D(n1723), .CLK(clk), .Q(EX_oprA[3]) );
  DFFPOSX1 EX_oprA_reg_4_ ( .D(n1724), .CLK(clk), .Q(EX_oprA[4]) );
  DFFPOSX1 EX_oprA_reg_5_ ( .D(n1725), .CLK(clk), .Q(EX_oprA[5]) );
  DFFPOSX1 EX_oprA_reg_6_ ( .D(n1726), .CLK(clk), .Q(EX_oprA[6]) );
  DFFPOSX1 EX_oprA_reg_7_ ( .D(n1727), .CLK(clk), .Q(EX_oprA[7]) );
  DFFPOSX1 EX_oprA_reg_8_ ( .D(n1728), .CLK(clk), .Q(EX_oprA[8]) );
  DFFPOSX1 EX_oprA_reg_9_ ( .D(n1729), .CLK(clk), .Q(EX_oprA[9]) );
  DFFPOSX1 EX_oprA_reg_10_ ( .D(n1730), .CLK(clk), .Q(EX_oprA[10]) );
  DFFPOSX1 EX_oprA_reg_11_ ( .D(n1731), .CLK(clk), .Q(EX_oprA[11]) );
  DFFPOSX1 EX_oprA_reg_12_ ( .D(n1732), .CLK(clk), .Q(EX_oprA[12]) );
  DFFPOSX1 EX_oprA_reg_13_ ( .D(n1733), .CLK(clk), .Q(EX_oprA[13]) );
  DFFPOSX1 EX_oprA_reg_14_ ( .D(n1734), .CLK(clk), .Q(EX_oprA[14]) );
  DFFPOSX1 EX_oprA_reg_15_ ( .D(n1735), .CLK(clk), .Q(EX_oprA[15]) );
  DFFPOSX1 EX_oprA_reg_16_ ( .D(n1736), .CLK(clk), .Q(EX_oprA[16]) );
  DFFPOSX1 EX_oprA_reg_17_ ( .D(n1737), .CLK(clk), .Q(EX_oprA[17]) );
  DFFPOSX1 EX_oprA_reg_18_ ( .D(n1738), .CLK(clk), .Q(EX_oprA[18]) );
  DFFPOSX1 EX_oprA_reg_19_ ( .D(n1739), .CLK(clk), .Q(EX_oprA[19]) );
  DFFPOSX1 EX_oprA_reg_20_ ( .D(n1740), .CLK(clk), .Q(EX_oprA[20]) );
  DFFPOSX1 EX_oprA_reg_21_ ( .D(n1741), .CLK(clk), .Q(EX_oprA[21]) );
  DFFPOSX1 EX_oprA_reg_22_ ( .D(n1742), .CLK(clk), .Q(EX_oprA[22]) );
  DFFPOSX1 EX_oprA_reg_23_ ( .D(n1743), .CLK(clk), .Q(EX_oprA[23]) );
  DFFPOSX1 EX_oprA_reg_24_ ( .D(n1744), .CLK(clk), .Q(EX_oprA[24]) );
  DFFPOSX1 EX_oprA_reg_25_ ( .D(n1745), .CLK(clk), .Q(EX_oprA[25]) );
  DFFPOSX1 EX_oprA_reg_26_ ( .D(n1746), .CLK(clk), .Q(EX_oprA[26]) );
  DFFPOSX1 EX_oprA_reg_27_ ( .D(n1747), .CLK(clk), .Q(EX_oprA[27]) );
  DFFPOSX1 EX_oprA_reg_28_ ( .D(n1748), .CLK(clk), .Q(EX_oprA[28]) );
  DFFPOSX1 EX_oprA_reg_29_ ( .D(n1749), .CLK(clk), .Q(EX_oprA[29]) );
  DFFPOSX1 EX_oprA_reg_30_ ( .D(n1750), .CLK(clk), .Q(EX_oprA[30]) );
  DFFPOSX1 EX_oprA_reg_31_ ( .D(n1751), .CLK(clk), .Q(EX_oprA[31]) );
  DFFPOSX1 EX_oprA_reg_32_ ( .D(n1752), .CLK(clk), .Q(EX_oprA[32]) );
  DFFPOSX1 EX_oprA_reg_33_ ( .D(n1753), .CLK(clk), .Q(EX_oprA[33]) );
  DFFPOSX1 EX_oprA_reg_34_ ( .D(n1754), .CLK(clk), .Q(EX_oprA[34]) );
  DFFPOSX1 EX_oprA_reg_35_ ( .D(n1755), .CLK(clk), .Q(EX_oprA[35]) );
  DFFPOSX1 EX_oprA_reg_36_ ( .D(n1756), .CLK(clk), .Q(EX_oprA[36]) );
  DFFPOSX1 EX_oprA_reg_37_ ( .D(n1757), .CLK(clk), .Q(EX_oprA[37]) );
  DFFPOSX1 EX_oprA_reg_38_ ( .D(n1758), .CLK(clk), .Q(EX_oprA[38]) );
  DFFPOSX1 EX_oprA_reg_39_ ( .D(n1759), .CLK(clk), .Q(EX_oprA[39]) );
  DFFPOSX1 EX_oprA_reg_40_ ( .D(n1760), .CLK(clk), .Q(EX_oprA[40]) );
  DFFPOSX1 EX_oprA_reg_41_ ( .D(n1761), .CLK(clk), .Q(EX_oprA[41]) );
  DFFPOSX1 EX_oprA_reg_42_ ( .D(n1762), .CLK(clk), .Q(EX_oprA[42]) );
  DFFPOSX1 EX_oprA_reg_43_ ( .D(n1763), .CLK(clk), .Q(EX_oprA[43]) );
  DFFPOSX1 EX_oprA_reg_44_ ( .D(n1764), .CLK(clk), .Q(EX_oprA[44]) );
  DFFPOSX1 EX_oprA_reg_45_ ( .D(n1765), .CLK(clk), .Q(EX_oprA[45]) );
  DFFPOSX1 EX_oprA_reg_46_ ( .D(n1766), .CLK(clk), .Q(EX_oprA[46]) );
  DFFPOSX1 EX_oprA_reg_47_ ( .D(n1767), .CLK(clk), .Q(EX_oprA[47]) );
  DFFPOSX1 EX_oprA_reg_48_ ( .D(n1768), .CLK(clk), .Q(EX_oprA[48]) );
  DFFPOSX1 EX_oprA_reg_49_ ( .D(n1769), .CLK(clk), .Q(EX_oprA[49]) );
  DFFPOSX1 EX_oprA_reg_50_ ( .D(n1770), .CLK(clk), .Q(EX_oprA[50]) );
  DFFPOSX1 EX_oprA_reg_51_ ( .D(n1771), .CLK(clk), .Q(EX_oprA[51]) );
  DFFPOSX1 EX_oprA_reg_52_ ( .D(n1772), .CLK(clk), .Q(EX_oprA[52]) );
  DFFPOSX1 EX_oprA_reg_53_ ( .D(n1773), .CLK(clk), .Q(EX_oprA[53]) );
  DFFPOSX1 EX_oprA_reg_54_ ( .D(n1774), .CLK(clk), .Q(EX_oprA[54]) );
  DFFPOSX1 EX_oprA_reg_55_ ( .D(n1775), .CLK(clk), .Q(EX_oprA[55]) );
  DFFPOSX1 EX_oprA_reg_56_ ( .D(n1776), .CLK(clk), .Q(EX_oprA[56]) );
  DFFPOSX1 EX_oprA_reg_57_ ( .D(n1777), .CLK(clk), .Q(EX_oprA[57]) );
  DFFPOSX1 EX_oprA_reg_58_ ( .D(n1778), .CLK(clk), .Q(EX_oprA[58]) );
  DFFPOSX1 EX_oprA_reg_59_ ( .D(n1779), .CLK(clk), .Q(EX_oprA[59]) );
  DFFPOSX1 EX_oprA_reg_60_ ( .D(n1780), .CLK(clk), .Q(EX_oprA[60]) );
  DFFPOSX1 EX_oprA_reg_61_ ( .D(n1781), .CLK(clk), .Q(EX_oprA[61]) );
  DFFPOSX1 EX_oprA_reg_62_ ( .D(n1782), .CLK(clk), .Q(EX_oprA[62]) );
  DFFPOSX1 EX_oprA_reg_63_ ( .D(n1783), .CLK(clk), .Q(EX_oprA[63]) );
  DFFPOSX1 ID_instruction_reg_2_ ( .D(n1995), .CLK(clk), .Q(ID_instruction[2])
         );
  DFFPOSX1 EX_is_mul32_reg ( .D(n1787), .CLK(clk), .Q(EX_is_mul32) );
  DFFPOSX1 EX_is_load_reg ( .D(n1786), .CLK(clk), .Q(EX_is_load) );
  DFFPOSX1 WB_is_load_reg ( .D(n2447), .CLK(clk), .Q(WB_is_load) );
  DFFPOSX1 EX_dest_reg_reg_0_ ( .D(n1794), .CLK(clk), .Q(EX_dest_reg[0]) );
  DFFPOSX1 WB_dest_reg_reg_0_ ( .D(n2450), .CLK(clk), .Q(WB_dest_reg[0]) );
  DFFPOSX1 EX_dest_reg_reg_1_ ( .D(n1795), .CLK(clk), .Q(EX_dest_reg[1]) );
  DFFPOSX1 WB_dest_reg_reg_1_ ( .D(n2451), .CLK(clk), .Q(WB_dest_reg[1]) );
  DFFPOSX1 EX_dest_reg_reg_2_ ( .D(n1796), .CLK(clk), .Q(EX_dest_reg[2]) );
  DFFPOSX1 WB_dest_reg_reg_2_ ( .D(n220), .CLK(clk), .Q(WB_dest_reg[2]) );
  DFFPOSX1 EX_dest_reg_reg_3_ ( .D(n1797), .CLK(clk), .Q(EX_dest_reg[3]) );
  DFFPOSX1 WB_dest_reg_reg_3_ ( .D(n219), .CLK(clk), .Q(WB_dest_reg[3]) );
  DFFPOSX1 EX_dest_reg_reg_4_ ( .D(n1798), .CLK(clk), .Q(EX_dest_reg[4]) );
  DFFPOSX1 WB_dest_reg_reg_4_ ( .D(n218), .CLK(clk), .Q(WB_dest_reg[4]) );
  DFFPOSX1 EX_shift_amt_reg_0_ ( .D(n1814), .CLK(clk), .Q(EX_shift_amt[0]) );
  DFFPOSX1 EX_shift_amt_reg_1_ ( .D(n1815), .CLK(clk), .Q(EX_shift_amt[1]) );
  DFFPOSX1 EX_shift_amt_reg_2_ ( .D(n1816), .CLK(clk), .Q(EX_shift_amt[2]) );
  DFFPOSX1 EX_shift_amt_reg_3_ ( .D(n1817), .CLK(clk), .Q(EX_shift_amt[3]) );
  DFFPOSX1 EX_shift_amt_reg_4_ ( .D(n1818), .CLK(clk), .Q(EX_shift_amt[4]) );
  DFFPOSX1 EX_PPP_reg_0_ ( .D(n1829), .CLK(clk), .Q(EX_PPP[0]) );
  DFFPOSX1 WB_PPP_reg_0_ ( .D(n217), .CLK(clk), .Q(WB_PPP[0]) );
  DFFPOSX1 EX_PPP_reg_1_ ( .D(n1830), .CLK(clk), .Q(EX_PPP[1]) );
  DFFPOSX1 WB_PPP_reg_1_ ( .D(n216), .CLK(clk), .Q(WB_PPP[1]) );
  DFFPOSX1 EX_PPP_reg_2_ ( .D(n1831), .CLK(clk), .Q(EX_PPP[2]) );
  DFFPOSX1 WB_PPP_reg_2_ ( .D(n215), .CLK(clk), .Q(WB_PPP[2]) );
  DFFPOSX1 EX_WW_reg_0_ ( .D(n1835), .CLK(clk), .Q(EX_WW[0]) );
  DFFPOSX1 EX_WW_reg_1_ ( .D(n1836), .CLK(clk), .Q(EX_WW[1]) );
  DFFPOSX1 EX_alu_func_reg_0_ ( .D(n1839), .CLK(clk), .Q(EX_alu_func[0]) );
  DFFPOSX1 EX_alu_func_reg_1_ ( .D(n1840), .CLK(clk), .Q(EX_alu_func[1]) );
  DFFPOSX1 EX_alu_func_reg_2_ ( .D(n1841), .CLK(clk), .Q(EX_alu_func[2]) );
  DFFPOSX1 EX_alu_func_reg_3_ ( .D(n1842), .CLK(clk), .Q(EX_alu_func[3]) );
  DFFPOSX1 EX_alu_func_reg_4_ ( .D(n1843), .CLK(clk), .Q(EX_alu_func[4]) );
  DFFPOSX1 EX_alu_func_reg_5_ ( .D(n1844), .CLK(clk), .Q(EX_alu_func[5]) );
  DFFPOSX1 PREVIOUS_STALL_reg ( .D(n2506), .CLK(clk), .Q(PREVIOUS_STALL) );
  DFFPOSX1 PREVIOUS_2_STALL_reg ( .D(n2452), .CLK(clk), .Q(PREVIOUS_2_STALL)
         );
  DFFPOSX1 EX_oprA_reg_0_ ( .D(n1720), .CLK(clk), .Q(EX_oprA[0]) );
  OAI21X1 U467 ( .A(n1920), .B(n3312), .C(n2041), .Y(n1786) );
  NAND3X1 U468 ( .A(n2500), .B(n3275), .C(n3284), .Y(n1178) );
  OAI21X1 U469 ( .A(n3311), .B(n2554), .C(n2040), .Y(n1787) );
  NAND3X1 U470 ( .A(n2500), .B(n3276), .C(n1183), .Y(n1181) );
  NOR3X1 U471 ( .A(n2473), .B(memAddr[25]), .C(n2441), .Y(n1183) );
  NAND3X1 U472 ( .A(n1920), .B(n2553), .C(n3281), .Y(n1788) );
  NAND3X1 U475 ( .A(n2073), .B(n2553), .C(n2088), .Y(n1790) );
  OAI21X1 U480 ( .A(n3309), .B(n1920), .C(n2210), .Y(n1792) );
  OAI21X1 U482 ( .A(n3277), .B(n2554), .C(n2196), .Y(n1793) );
  OAI21X1 U484 ( .A(n3308), .B(n2559), .C(n2229), .Y(n1794) );
  OAI21X1 U486 ( .A(n3307), .B(n2559), .C(n2348), .Y(n1795) );
  OAI21X1 U488 ( .A(n3306), .B(n2556), .C(n2249), .Y(n1796) );
  OAI21X1 U490 ( .A(n3305), .B(n2559), .C(n2312), .Y(n1797) );
  OAI21X1 U492 ( .A(n3304), .B(n2559), .C(n2392), .Y(n1798) );
  OAI21X1 U494 ( .A(n3308), .B(n1920), .C(n2455), .Y(n1799) );
  OAI21X1 U496 ( .A(n3307), .B(n2554), .C(n2416), .Y(n1800) );
  OAI21X1 U498 ( .A(n3306), .B(n1920), .C(n2386), .Y(n1801) );
  OAI21X1 U500 ( .A(n3305), .B(n2554), .C(n2343), .Y(n1802) );
  OAI21X1 U502 ( .A(n3304), .B(n1920), .C(n2285), .Y(n1803) );
  OAI21X1 U504 ( .A(n3303), .B(n2485), .C(n2385), .Y(n1804) );
  OAI21X1 U506 ( .A(n3303), .B(n2554), .C(n2307), .Y(n1805) );
  OAI21X1 U508 ( .A(n3302), .B(n2485), .C(n2342), .Y(n1806) );
  OAI21X1 U510 ( .A(n3302), .B(n1920), .C(n2262), .Y(n1807) );
  OAI21X1 U512 ( .A(n3301), .B(n2485), .C(n2341), .Y(n1808) );
  OAI21X1 U514 ( .A(n3301), .B(n2554), .C(n2243), .Y(n1809) );
  OAI21X1 U516 ( .A(n3300), .B(n2485), .C(n2384), .Y(n1810) );
  OAI21X1 U518 ( .A(n3300), .B(n1920), .C(n2224), .Y(n1811) );
  OAI21X1 U520 ( .A(n3299), .B(n2485), .C(n2340), .Y(n1812) );
  OAI21X1 U522 ( .A(n3299), .B(n2554), .C(n2454), .Y(n1813) );
  OAI21X1 U524 ( .A(n2579), .B(n2559), .C(n2146), .Y(n1814) );
  OAI21X1 U526 ( .A(n2578), .B(n2556), .C(n2159), .Y(n1815) );
  OAI21X1 U528 ( .A(n2577), .B(n2555), .C(n2172), .Y(n1816) );
  OAI21X1 U530 ( .A(n2575), .B(n2559), .C(n2187), .Y(n1817) );
  OAI21X1 U532 ( .A(n2573), .B(n2555), .C(n2421), .Y(n1818) );
  OAI21X1 U534 ( .A(n2579), .B(n2485), .C(n2339), .Y(n1819) );
  OAI21X1 U536 ( .A(n2579), .B(n1920), .C(n2209), .Y(n1820) );
  OAI21X1 U538 ( .A(n2578), .B(n2485), .C(n2383), .Y(n1821) );
  OAI21X1 U540 ( .A(n2578), .B(n2554), .C(n2195), .Y(n1822) );
  OAI21X1 U542 ( .A(n2577), .B(n2485), .C(n2338), .Y(n1823) );
  OAI21X1 U544 ( .A(n2577), .B(n1920), .C(n2182), .Y(n1824) );
  OAI21X1 U546 ( .A(n2575), .B(n2485), .C(n2337), .Y(n1825) );
  OAI21X1 U548 ( .A(n2575), .B(n2554), .C(n2167), .Y(n1826) );
  OAI21X1 U550 ( .A(n2573), .B(n2485), .C(n2336), .Y(n1827) );
  OAI21X1 U552 ( .A(n2573), .B(n1920), .C(n2154), .Y(n1828) );
  OAI21X1 U554 ( .A(n3298), .B(n2555), .C(n2201), .Y(n1829) );
  OAI21X1 U556 ( .A(n2555), .B(n3297), .C(n2215), .Y(n1830) );
  OAI21X1 U558 ( .A(n2556), .B(n3296), .C(n2230), .Y(n1831) );
  OAI21X1 U560 ( .A(n3298), .B(n2554), .C(n2141), .Y(n1832) );
  OAI21X1 U562 ( .A(n2554), .B(n3297), .C(n2415), .Y(n1833) );
  OAI21X1 U564 ( .A(n2554), .B(n3296), .C(n2382), .Y(n1834) );
  OAI21X1 U566 ( .A(n3295), .B(n2556), .C(n2250), .Y(n1835) );
  OAI21X1 U568 ( .A(n3294), .B(n2555), .C(n2268), .Y(n1836) );
  OAI21X1 U570 ( .A(n3295), .B(n2554), .C(n2335), .Y(n1837) );
  OAI21X1 U572 ( .A(n3294), .B(n1920), .C(n2306), .Y(n1838) );
  OAI21X1 U574 ( .A(n2555), .B(n3293), .C(n2290), .Y(n1839) );
  OAI21X1 U576 ( .A(n2559), .B(n3280), .C(n2313), .Y(n1840) );
  OAI21X1 U578 ( .A(n3292), .B(n2555), .C(n2349), .Y(n1841) );
  OAI21X1 U580 ( .A(n3291), .B(n2556), .C(n2393), .Y(n1842) );
  OAI21X1 U582 ( .A(n2556), .B(n3289), .C(n2422), .Y(n1843) );
  OAI21X1 U584 ( .A(n3288), .B(n2559), .C(n2461), .Y(n1844) );
  OAI21X1 U586 ( .A(n1920), .B(n3293), .C(n2261), .Y(n1845) );
  OAI21X1 U588 ( .A(n2554), .B(n3280), .C(n2284), .Y(n1846) );
  OAI21X1 U590 ( .A(n3292), .B(n2554), .C(n2242), .Y(n1847) );
  OAI21X1 U592 ( .A(n3291), .B(n1920), .C(n2223), .Y(n1848) );
  OAI21X1 U594 ( .A(n1920), .B(n3289), .C(n2208), .Y(n1849) );
  OAI21X1 U596 ( .A(n3288), .B(n1920), .C(n2136), .Y(n1850) );
  OAI21X1 U722 ( .A(n1920), .B(n2488), .C(n2241), .Y(n1913) );
  OAI21X1 U777 ( .A(n3282), .B(n2472), .C(n2325), .Y(memEn) );
  OAI21X1 U780 ( .A(n3311), .B(n1361), .C(n2297), .Y(n1360) );
  NAND3X1 U781 ( .A(n2298), .B(n1364), .C(n1365), .Y(n1362) );
  NOR3X1 U782 ( .A(n1366), .B(n1367), .C(n1368), .Y(n1365) );
  XOR2X1 U783 ( .A(ID_instruction[6]), .B(EX_dest_reg[0]), .Y(n1368) );
  XOR2X1 U784 ( .A(ID_instruction[10]), .B(EX_dest_reg[4]), .Y(n1367) );
  XOR2X1 U785 ( .A(ID_instruction[9]), .B(EX_dest_reg[3]), .Y(n1366) );
  XOR2X1 U786 ( .A(n3306), .B(EX_dest_reg[2]), .Y(n1364) );
  AOI21X1 U787 ( .A(n1369), .B(n1370), .C(n1371), .Y(n1363) );
  XOR2X1 U788 ( .A(ID_instruction[7]), .B(EX_dest_reg[1]), .Y(n1371) );
  OAI21X1 U789 ( .A(n3273), .B(n3274), .C(n3275), .Y(n1370) );
  OAI21X1 U792 ( .A(EX_is_load), .B(EX_reg_write), .C(n3272), .Y(n1369) );
  OAI21X1 U793 ( .A(n1375), .B(n1376), .C(n1313), .Y(n1361) );
  NOR3X1 U794 ( .A(n2429), .B(n1378), .C(n1379), .Y(n1376) );
  XOR2X1 U795 ( .A(ID_instruction[11]), .B(EX_dest_reg[0]), .Y(n1379) );
  XOR2X1 U796 ( .A(ID_instruction[14]), .B(EX_dest_reg[3]), .Y(n1378) );
  NAND3X1 U797 ( .A(n1380), .B(n1381), .C(n1382), .Y(n1377) );
  XOR2X1 U798 ( .A(n3299), .B(EX_dest_reg[4]), .Y(n1382) );
  XOR2X1 U799 ( .A(n3302), .B(EX_dest_reg[1]), .Y(n1381) );
  XOR2X1 U800 ( .A(n3301), .B(EX_dest_reg[2]), .Y(n1380) );
  NOR3X1 U801 ( .A(n2465), .B(n1384), .C(n1385), .Y(n1375) );
  XOR2X1 U802 ( .A(memAddr[16]), .B(EX_dest_reg[0]), .Y(n1385) );
  XOR2X1 U803 ( .A(memAddr[19]), .B(EX_dest_reg[3]), .Y(n1384) );
  NAND3X1 U804 ( .A(n1386), .B(n1387), .C(n1388), .Y(n1383) );
  XOR2X1 U805 ( .A(n2573), .B(EX_dest_reg[4]), .Y(n1388) );
  XOR2X1 U806 ( .A(n2578), .B(EX_dest_reg[1]), .Y(n1387) );
  XOR2X1 U807 ( .A(n2577), .B(EX_dest_reg[2]), .Y(n1386) );
  NAND3X1 U808 ( .A(n3313), .B(n3314), .C(n1389), .Y(n1359) );
  NOR3X1 U809 ( .A(EX_dest_reg[2]), .B(EX_dest_reg[4]), .C(EX_dest_reg[3]), 
        .Y(n1389) );
  NAND3X1 U811 ( .A(n3309), .B(n3277), .C(n2517), .Y(n1180) );
  NOR3X1 U812 ( .A(n2361), .B(ID_instruction[15]), .C(ID_instruction[14]), .Y(
        n1393) );
  NAND3X1 U813 ( .A(n3310), .B(n3287), .C(n3286), .Y(n1394) );
  NOR3X1 U814 ( .A(n2323), .B(ID_instruction[11]), .C(n3285), .Y(n1392) );
  OAI21X1 U816 ( .A(n1313), .B(n3304), .C(n2319), .Y(ID_rf_rd1_addr[4]) );
  OAI21X1 U818 ( .A(n1313), .B(n3305), .C(n2428), .Y(ID_rf_rd1_addr[3]) );
  OAI21X1 U820 ( .A(n1313), .B(n3306), .C(n2355), .Y(ID_rf_rd1_addr[2]) );
  OAI21X1 U822 ( .A(n1313), .B(n3307), .C(n2399), .Y(ID_rf_rd1_addr[1]) );
  OAI21X1 U824 ( .A(n1313), .B(n3308), .C(n2296), .Y(ID_rf_rd1_addr[0]) );
  NAND3X1 U828 ( .A(ID_instruction[2]), .B(ID_instruction[0]), .C(
        ID_instruction[4]), .Y(n1402) );
  NAND3X1 U829 ( .A(n3287), .B(n3277), .C(n3286), .Y(n1401) );
  AOI22X1 U833 ( .A(n1407), .B(n3289), .C(memAddr[25]), .D(n3290), .Y(n1406)
         );
  NAND3X1 U834 ( .A(memAddr[28]), .B(n3291), .C(memAddr[24]), .Y(n1185) );
  OAI21X1 U835 ( .A(n3291), .B(n1408), .C(n2039), .Y(n1407) );
  NAND3X1 U836 ( .A(n3291), .B(n3288), .C(n3292), .Y(n1409) );
  OAI21X1 U837 ( .A(n3292), .B(n3288), .C(n2038), .Y(n1408) );
  NAND3X1 U838 ( .A(n2579), .B(n2578), .C(n1411), .Y(n1410) );
  NOR3X1 U839 ( .A(memAddr[18]), .B(memAddr[20]), .C(memAddr[19]), .Y(n1411)
         );
  AOI21X1 U840 ( .A(n3296), .B(n3297), .C(n3298), .Y(n1404) );
  program_counter PC ( .clk(clk), .reset(reset), .stall(n3283), .pc_load(n3270), .data_in(memAddr[16:31]), .data_out(pc) );
  register_file reg_file ( .clk(clk), .reset(reset), .write_en(
        WB_reg_write_load), .read1_addr(ID_rf_rd1_addr), .read2_addr(
        memAddr[16:20]), .write_addr(WB_dest_reg), .Din({WB_data[0], n2477, 
        n2374, n2443, n2220, n2280, n2411, WB_data[7:14], n1927, WB_data[16], 
        n2303, WB_data[18], n2177, WB_data[20], n1938, n2378, n1928, 
        WB_data[24:31], n2331, n2205, n2238, n2162, n2191, n2258, n2519, n2518, 
        WB_data[40:63]}), .Dout1(dataOut), .Dout2(ID_oprB), .PPP({WB_PPP[0:1], 
        n2486}) );
  alu ALU ( .clk(clk), .oprA({n2334, EX_alu_A[1:10], n2570, EX_alu_A[12:14], 
        n2568, EX_alu_A[16:41], n2469, EX_alu_A[43:47], n2567, EX_alu_A[49:63]}), .oprB({EX_alu_B[0:24], n2685, EX_alu_B[26:30], n2407, EX_alu_B[32:63]}), 
        .shift_amount(EX_shift_amt), .op(EX_alu_func), .ww(EX_WW), .result(
        EX_alu_result), .mult32_result(WB_mult32_result) );
  BUFX2 U1341 ( .A(WB_mult32_result[7]), .Y(n1915) );
  INVX2 U1342 ( .A(WB_mult32_result[14]), .Y(n2901) );
  AND2X2 U1343 ( .A(n2494), .B(WB_is_mul32), .Y(n1918) );
  INVX2 U1344 ( .A(n2544), .Y(n2540) );
  BUFX4 U1345 ( .A(n2869), .Y(n2490) );
  AND2X2 U1346 ( .A(EX_alu_result[0]), .B(n2553), .Y(n287) );
  AND2X2 U1347 ( .A(EX_alu_result[1]), .B(n2553), .Y(n286) );
  AND2X2 U1348 ( .A(n2684), .B(WB_data[24]), .Y(n2686) );
  INVX8 U1349 ( .A(n2804), .Y(n2133) );
  INVX1 U1350 ( .A(n2535), .Y(n1916) );
  INVX2 U1351 ( .A(n1916), .Y(n1917) );
  AND2X2 U1352 ( .A(n2413), .B(n2412), .Y(WB_data[6]) );
  INVX1 U1353 ( .A(n2403), .Y(n2756) );
  AND2X1 U1354 ( .A(n2504), .B(WB_data[16]), .Y(n2706) );
  AND2X1 U1355 ( .A(n2504), .B(n2374), .Y(n2732) );
  BUFX2 U1356 ( .A(n2923), .Y(n2494) );
  AND2X1 U1357 ( .A(EX_oprB[28]), .B(n2484), .Y(n2668) );
  AND2X1 U1358 ( .A(n2505), .B(n2162), .Y(n2644) );
  INVX1 U1359 ( .A(n2545), .Y(n2134) );
  AND2X1 U1360 ( .A(n2684), .B(WB_data[13]), .Y(n2709) );
  AND2X1 U1361 ( .A(n2512), .B(n2414), .Y(n2508) );
  AND2X1 U1362 ( .A(n2504), .B(WB_data[7]), .Y(n2717) );
  AND2X1 U1363 ( .A(n2684), .B(WB_data[8]), .Y(n2714) );
  AND2X1 U1364 ( .A(n2684), .B(WB_data[9]), .Y(n2713) );
  AND2X1 U1365 ( .A(n2504), .B(n2378), .Y(n2693) );
  OR2X1 U1366 ( .A(n2566), .B(n2482), .Y(n2892) );
  AND2X1 U1367 ( .A(n1918), .B(WB_mult32_result[20]), .Y(n1934) );
  AND2X1 U1368 ( .A(EX_oprA[20]), .B(n2537), .Y(n1935) );
  OR2X1 U1369 ( .A(n2566), .B(n2789), .Y(n2790) );
  OR2X1 U1370 ( .A(n2566), .B(n2776), .Y(n2778) );
  AND2X1 U1371 ( .A(n2505), .B(n2518), .Y(n2632) );
  AND2X1 U1372 ( .A(n2503), .B(WB_data[40]), .Y(n2628) );
  AND2X1 U1373 ( .A(n2503), .B(WB_data[41]), .Y(n2627) );
  AND2X1 U1374 ( .A(n2503), .B(WB_data[47]), .Y(n2621) );
  AND2X1 U1375 ( .A(n2505), .B(WB_data[49]), .Y(n2618) );
  INVX1 U1376 ( .A(WB_PPP[0]), .Y(n2592) );
  INVX1 U1377 ( .A(WB_PPP[1]), .Y(n2591) );
  AND2X1 U1378 ( .A(n2505), .B(WB_data[50]), .Y(n2617) );
  AND2X1 U1379 ( .A(n2505), .B(WB_data[51]), .Y(n2616) );
  AND2X1 U1380 ( .A(n2505), .B(WB_data[55]), .Y(n2611) );
  OR2X1 U1381 ( .A(n2566), .B(n2801), .Y(n2802) );
  INVX1 U1382 ( .A(n2602), .Y(n2600) );
  AND2X1 U1383 ( .A(n2495), .B(n2566), .Y(n2515) );
  INVX1 U1384 ( .A(n2868), .Y(n2866) );
  INVX1 U1385 ( .A(n2509), .Y(n2536) );
  INVX1 U1386 ( .A(n2510), .Y(n2537) );
  AND2X1 U1387 ( .A(n2329), .B(n2924), .Y(n2926) );
  AND2X1 U1388 ( .A(n2963), .B(n2481), .Y(n2870) );
  AND2X1 U1389 ( .A(n2504), .B(n1928), .Y(n2690) );
  INVX1 U1390 ( .A(n2509), .Y(n2535) );
  OR2X1 U1391 ( .A(n2566), .B(n2797), .Y(n2798) );
  AND2X1 U1392 ( .A(n2505), .B(n2238), .Y(n2647) );
  AND2X1 U1393 ( .A(n2463), .B(n2135), .Y(n2522) );
  AND2X1 U1394 ( .A(n2127), .B(n2612), .Y(n2782) );
  INVX1 U1395 ( .A(n2367), .Y(n2750) );
  INVX1 U1396 ( .A(n2515), .Y(n2552) );
  INVX2 U1397 ( .A(n2552), .Y(n2547) );
  BUFX2 U1398 ( .A(WB_PPP[2]), .Y(n2486) );
  AND2X1 U1399 ( .A(n2977), .B(n2976), .Y(n2982) );
  AND2X1 U1400 ( .A(n2684), .B(n2683), .Y(n1936) );
  INVX2 U1401 ( .A(n2502), .Y(n2922) );
  OR2X1 U1402 ( .A(n2474), .B(n2656), .Y(n2655) );
  AND2X1 U1403 ( .A(n2514), .B(n2446), .Y(n2679) );
  AND2X1 U1404 ( .A(n2505), .B(n2331), .Y(n2653) );
  AND2X1 U1405 ( .A(n1956), .B(n1957), .Y(EX_alu_A[48]) );
  INVX2 U1406 ( .A(n2133), .Y(n2135) );
  INVX1 U1407 ( .A(n2491), .Y(n2493) );
  INVX1 U1408 ( .A(n2278), .Y(n2748) );
  INVX2 U1409 ( .A(n2544), .Y(n2542) );
  AND2X1 U1410 ( .A(n2151), .B(n2150), .Y(WB_data[39]) );
  AND2X1 U1411 ( .A(n2332), .B(n2333), .Y(WB_data[32]) );
  INVX1 U1412 ( .A(WB_mult32_result[24]), .Y(n2876) );
  INVX1 U1413 ( .A(WB_mult32_result[18]), .Y(n2887) );
  AND2X1 U1414 ( .A(n2304), .B(n2305), .Y(WB_data[17]) );
  INVX1 U1415 ( .A(WB_mult32_result[15]), .Y(n2526) );
  INVX1 U1416 ( .A(WB_mult32_result[13]), .Y(n2521) );
  INVX1 U1417 ( .A(WB_mult32_result[12]), .Y(n2528) );
  INVX1 U1418 ( .A(WB_mult32_result[11]), .Y(n2530) );
  INVX1 U1419 ( .A(WB_mult32_result[10]), .Y(n2914) );
  INVX1 U1420 ( .A(WB_mult32_result[8]), .Y(n2921) );
  AND2X1 U1421 ( .A(n2282), .B(n2283), .Y(WB_data[5]) );
  AND2X1 U1422 ( .A(n2375), .B(n2376), .Y(WB_data[2]) );
  AND2X1 U1423 ( .A(WB_mult32_result[1]), .B(n2561), .Y(n2733) );
  BUFX2 U1424 ( .A(n2149), .Y(n2518) );
  INVX1 U1425 ( .A(WB_data[36]), .Y(n2191) );
  AND2X1 U1426 ( .A(n2164), .B(n2163), .Y(WB_data[35]) );
  AND2X1 U1427 ( .A(n2206), .B(n2207), .Y(WB_data[33]) );
  INVX1 U1428 ( .A(WB_mult32_result[30]), .Y(n2953) );
  INVX1 U1429 ( .A(WB_data[5]), .Y(n2280) );
  INVX1 U1430 ( .A(WB_data[3]), .Y(n2443) );
  INVX1 U1431 ( .A(WB_mult32_result[0]), .Y(n2736) );
  OR2X1 U1432 ( .A(n2363), .B(n2473), .Y(n1405) );
  OR2X1 U1433 ( .A(n2071), .B(n2072), .Y(n3013) );
  AND2X1 U1434 ( .A(n3008), .B(n3275), .Y(n3270) );
  AND2X1 U1435 ( .A(EX_regA[0]), .B(n2485), .Y(n1203) );
  AND2X1 U1436 ( .A(EX_regA[1]), .B(n2485), .Y(n1205) );
  AND2X1 U1437 ( .A(EX_regA[2]), .B(n2485), .Y(n1207) );
  AND2X1 U1438 ( .A(EX_regA[3]), .B(n2485), .Y(n1209) );
  AND2X1 U1439 ( .A(EX_regA[4]), .B(n2485), .Y(n1211) );
  AND2X1 U1440 ( .A(EX_regB[0]), .B(n2485), .Y(n1218) );
  AND2X1 U1441 ( .A(EX_regB[1]), .B(n2485), .Y(n1220) );
  AND2X1 U1442 ( .A(EX_regB[2]), .B(n2485), .Y(n1222) );
  AND2X1 U1443 ( .A(EX_regB[3]), .B(n2485), .Y(n1224) );
  AND2X1 U1444 ( .A(EX_regB[4]), .B(n2485), .Y(n1226) );
  AND2X1 U1445 ( .A(n2359), .B(n2553), .Y(n1791) );
  AND2X1 U1446 ( .A(n2322), .B(n2553), .Y(n1789) );
  INVX1 U1447 ( .A(WB_mult32_result[28]), .Y(n2527) );
  INVX2 U1448 ( .A(n2128), .Y(n2684) );
  INVX2 U1449 ( .A(memAddr[17]), .Y(n2578) );
  INVX4 U1450 ( .A(n2501), .Y(n2843) );
  INVX1 U1451 ( .A(n2506), .Y(n1919) );
  INVX1 U1452 ( .A(n2506), .Y(n1920) );
  AND2X2 U1453 ( .A(n3283), .B(n2553), .Y(n2506) );
  INVX1 U1454 ( .A(n2487), .Y(n2741) );
  INVX1 U1455 ( .A(WB_mult32_result[29]), .Y(n2955) );
  INVX1 U1456 ( .A(n2679), .Y(n2484) );
  INVX1 U1457 ( .A(n2516), .Y(n2545) );
  INVX1 U1458 ( .A(n2544), .Y(n2539) );
  AND2X1 U1459 ( .A(n2370), .B(n2553), .Y(n1202) );
  OR2X1 U1460 ( .A(n2682), .B(n1936), .Y(n2685) );
  AND2X1 U1461 ( .A(WB_data[15]), .B(n2684), .Y(n2707) );
  BUFX2 U1462 ( .A(n2526), .Y(n1921) );
  OR2X2 U1463 ( .A(n1934), .B(n1935), .Y(n2884) );
  INVX1 U1464 ( .A(n2884), .Y(n1922) );
  AND2X1 U1465 ( .A(n2446), .B(n2132), .Y(n1933) );
  INVX1 U1466 ( .A(n2527), .Y(n1923) );
  INVX8 U1467 ( .A(n2552), .Y(n2546) );
  AND2X1 U1468 ( .A(n2511), .B(n2111), .Y(n1991) );
  INVX2 U1469 ( .A(n2544), .Y(n2496) );
  INVX1 U1470 ( .A(n2544), .Y(n2497) );
  INVX1 U1471 ( .A(WB_mult32_result[16]), .Y(n2705) );
  INVX2 U1472 ( .A(n2516), .Y(n2544) );
  INVX2 U1473 ( .A(WB_data[34]), .Y(n2238) );
  OAI21X1 U1474 ( .A(WB_reg_write), .B(WB_is_load), .C(n2581), .Y(n1924) );
  INVX4 U1475 ( .A(n2571), .Y(n2570) );
  INVX8 U1476 ( .A(n2533), .Y(n2534) );
  INVX1 U1477 ( .A(WB_mult32_result[25]), .Y(n2963) );
  INVX1 U1478 ( .A(WB_mult32_result[20]), .Y(n2883) );
  INVX1 U1479 ( .A(n2531), .Y(n1925) );
  AND2X2 U1480 ( .A(n2503), .B(WB_data[57]), .Y(n2608) );
  INVX1 U1481 ( .A(n2955), .Y(n1926) );
  INVX4 U1482 ( .A(WB_data[37]), .Y(n2258) );
  OAI21X1 U1483 ( .A(n2563), .B(n1921), .C(n2237), .Y(n1927) );
  INVX2 U1484 ( .A(n1953), .Y(n1929) );
  AND2X2 U1485 ( .A(n2501), .B(WB_mult32_result[42]), .Y(n2520) );
  OR2X2 U1486 ( .A(n2687), .B(n2113), .Y(n1928) );
  INVX2 U1487 ( .A(WB_mult32_result[31]), .Y(n2529) );
  INVX4 U1488 ( .A(n2498), .Y(n2499) );
  INVX1 U1489 ( .A(n2959), .Y(n1930) );
  AND2X2 U1490 ( .A(n2505), .B(n2191), .Y(n2641) );
  AND2X2 U1491 ( .A(n2504), .B(n2477), .Y(n2735) );
  INVX1 U1492 ( .A(WB_data[1]), .Y(n2477) );
  INVX1 U1493 ( .A(n2219), .Y(n1931) );
  INVX2 U1494 ( .A(n2492), .Y(n2629) );
  INVX1 U1495 ( .A(WB_mult32_result[26]), .Y(n1932) );
  INVX1 U1496 ( .A(WB_mult32_result[26]), .Y(n2961) );
  INVX8 U1497 ( .A(WB_is_mul32), .Y(n2566) );
  AND2X2 U1498 ( .A(n2512), .B(n1933), .Y(n2531) );
  AND2X2 U1499 ( .A(n2589), .B(n2588), .Y(n2511) );
  AND2X1 U1500 ( .A(WB_mult32_result[23]), .B(n2561), .Y(n2687) );
  INVX1 U1501 ( .A(EX_reg_write), .Y(n2488) );
  AND2X2 U1502 ( .A(n2107), .B(n2562), .Y(n2501) );
  AND2X1 U1503 ( .A(WB_mult32_result[2]), .B(n2562), .Y(n2730) );
  AND2X1 U1504 ( .A(EX_alu_result[32]), .B(n2553), .Y(n255) );
  INVX8 U1505 ( .A(n2569), .Y(n2568) );
  INVX1 U1506 ( .A(n2961), .Y(n1937) );
  AND2X2 U1507 ( .A(n2562), .B(n1937), .Y(n2677) );
  AND2X2 U1508 ( .A(n2684), .B(WB_data[10]), .Y(n2712) );
  OR2X2 U1509 ( .A(n2694), .B(n2115), .Y(n1938) );
  AND2X1 U1510 ( .A(EX_alu_result[33]), .B(n2553), .Y(n254) );
  INVX2 U1511 ( .A(WB_mult32_result[27]), .Y(n2959) );
  INVX1 U1512 ( .A(n2778), .Y(n1939) );
  INVX1 U1513 ( .A(n2790), .Y(n1940) );
  INVX1 U1514 ( .A(n2798), .Y(n1941) );
  INVX1 U1515 ( .A(n2617), .Y(n1942) );
  INVX1 U1516 ( .A(n2618), .Y(n1943) );
  AND2X2 U1517 ( .A(n2505), .B(WB_data[48]), .Y(n2620) );
  INVX1 U1518 ( .A(n2620), .Y(n1944) );
  AND2X2 U1519 ( .A(n2503), .B(WB_data[43]), .Y(n2625) );
  INVX1 U1520 ( .A(n2625), .Y(n1945) );
  INVX1 U1521 ( .A(n2628), .Y(n1946) );
  INVX1 U1522 ( .A(n2653), .Y(n1947) );
  INVX1 U1523 ( .A(n2686), .Y(n1948) );
  AND2X2 U1524 ( .A(n2504), .B(WB_data[20]), .Y(n2697) );
  INVX1 U1525 ( .A(n2697), .Y(n1949) );
  INVX1 U1526 ( .A(n2706), .Y(n1950) );
  AND2X2 U1527 ( .A(n2684), .B(WB_data[14]), .Y(n2708) );
  INVX1 U1528 ( .A(n2708), .Y(n1951) );
  INVX1 U1529 ( .A(n2709), .Y(n1952) );
  AND2X2 U1530 ( .A(n2489), .B(n2105), .Y(n2766) );
  INVX1 U1531 ( .A(n2766), .Y(n1953) );
  AND2X2 U1532 ( .A(n1990), .B(n1998), .Y(n2804) );
  INVX1 U1533 ( .A(n2782), .Y(n1954) );
  OR2X2 U1534 ( .A(n2887), .B(n2566), .Y(n2888) );
  INVX1 U1535 ( .A(n2888), .Y(n1955) );
  BUFX2 U1536 ( .A(n2809), .Y(n1956) );
  BUFX2 U1537 ( .A(n2808), .Y(n1957) );
  BUFX2 U1538 ( .A(n2751), .Y(n1958) );
  BUFX2 U1539 ( .A(n2754), .Y(n1959) );
  BUFX2 U1540 ( .A(n2760), .Y(n1960) );
  BUFX2 U1541 ( .A(n2764), .Y(n1961) );
  BUFX2 U1542 ( .A(n2791), .Y(n1962) );
  BUFX2 U1543 ( .A(n2813), .Y(n1963) );
  BUFX2 U1544 ( .A(n2822), .Y(n1964) );
  BUFX2 U1545 ( .A(n2826), .Y(n1965) );
  BUFX2 U1546 ( .A(n2829), .Y(n1966) );
  BUFX2 U1547 ( .A(n2837), .Y(n1967) );
  BUFX2 U1548 ( .A(n2841), .Y(n1968) );
  BUFX2 U1549 ( .A(n2859), .Y(n1969) );
  BUFX2 U1550 ( .A(n2889), .Y(n1970) );
  INVX1 U1551 ( .A(n2611), .Y(n1971) );
  INVX1 U1552 ( .A(n2616), .Y(n1972) );
  INVX1 U1553 ( .A(n2627), .Y(n1973) );
  INVX1 U1554 ( .A(n2693), .Y(n1974) );
  AND2X2 U1555 ( .A(n2504), .B(n1938), .Y(n2696) );
  INVX1 U1556 ( .A(n2696), .Y(n1975) );
  AND2X2 U1557 ( .A(n2504), .B(n2177), .Y(n2700) );
  INVX1 U1558 ( .A(n2700), .Y(n1976) );
  AND2X2 U1559 ( .A(n2504), .B(n2303), .Y(n2704) );
  INVX1 U1560 ( .A(n2704), .Y(n1977) );
  INVX1 U1561 ( .A(n2707), .Y(n1978) );
  AND2X2 U1562 ( .A(n2684), .B(WB_data[11]), .Y(n2711) );
  INVX1 U1563 ( .A(n2711), .Y(n1979) );
  AND2X2 U1564 ( .A(n2504), .B(n2411), .Y(n2720) );
  INVX1 U1565 ( .A(n2720), .Y(n1980) );
  AND2X2 U1566 ( .A(n2504), .B(n2281), .Y(n2723) );
  INVX1 U1567 ( .A(n2723), .Y(n1981) );
  AND2X2 U1568 ( .A(n2504), .B(n2219), .Y(n2726) );
  INVX1 U1569 ( .A(n2726), .Y(n1982) );
  AND2X2 U1570 ( .A(n2504), .B(n2443), .Y(n2729) );
  INVX1 U1571 ( .A(n2729), .Y(n1983) );
  INVX1 U1572 ( .A(n2732), .Y(n1984) );
  AND2X2 U1573 ( .A(n2504), .B(WB_data[0]), .Y(n2737) );
  INVX1 U1574 ( .A(n2737), .Y(n1985) );
  AND2X1 U1575 ( .A(WB_mult32_result[21]), .B(n2561), .Y(n2694) );
  BUFX2 U1576 ( .A(n2744), .Y(n1986) );
  BUFX2 U1577 ( .A(n2783), .Y(n1987) );
  INVX1 U1578 ( .A(n2870), .Y(n1988) );
  OR2X2 U1579 ( .A(n1986), .B(n2070), .Y(n2879) );
  INVX1 U1580 ( .A(n2879), .Y(n1989) );
  INVX1 U1581 ( .A(n2879), .Y(n1990) );
  AND2X2 U1582 ( .A(n2684), .B(WB_data[12]), .Y(n2710) );
  INVX8 U1583 ( .A(n2531), .Y(n2532) );
  INVX1 U1584 ( .A(n2522), .Y(n1992) );
  BUFX2 U1585 ( .A(n2788), .Y(n1993) );
  BUFX2 U1586 ( .A(n2938), .Y(n1994) );
  BUFX2 U1587 ( .A(n1790), .Y(n1995) );
  BUFX2 U1588 ( .A(n1788), .Y(n1996) );
  OR2X1 U1589 ( .A(n2555), .B(n2106), .Y(n1914) );
  INVX1 U1590 ( .A(n1914), .Y(n1997) );
  BUFX2 U1591 ( .A(n2775), .Y(n1998) );
  INVX1 U1592 ( .A(n2937), .Y(n1999) );
  INVX1 U1593 ( .A(n1999), .Y(n2000) );
  INVX1 U1594 ( .A(n2594), .Y(n2001) );
  INVX1 U1595 ( .A(n2001), .Y(n2002) );
  BUFX2 U1596 ( .A(n2597), .Y(n2003) );
  INVX1 U1597 ( .A(n2599), .Y(n2004) );
  INVX1 U1598 ( .A(n2004), .Y(n2005) );
  INVX1 U1599 ( .A(n2601), .Y(n2006) );
  INVX1 U1600 ( .A(n2006), .Y(n2007) );
  BUFX2 U1601 ( .A(n2603), .Y(n2008) );
  BUFX2 U1602 ( .A(n2604), .Y(n2009) );
  INVX1 U1603 ( .A(n2749), .Y(n2010) );
  INVX1 U1604 ( .A(n2010), .Y(n2011) );
  BUFX2 U1605 ( .A(n2773), .Y(n2012) );
  BUFX2 U1606 ( .A(n2779), .Y(n2013) );
  BUFX2 U1607 ( .A(n2799), .Y(n2014) );
  INVX1 U1608 ( .A(n2803), .Y(n2015) );
  INVX1 U1609 ( .A(n2015), .Y(n2016) );
  INVX1 U1610 ( .A(n2818), .Y(n2017) );
  INVX1 U1611 ( .A(n2017), .Y(n2018) );
  BUFX2 U1612 ( .A(n2857), .Y(n2019) );
  INVX1 U1613 ( .A(n2861), .Y(n2020) );
  INVX1 U1614 ( .A(n2020), .Y(n2021) );
  BUFX2 U1615 ( .A(n2863), .Y(n2022) );
  BUFX2 U1616 ( .A(n2864), .Y(n2023) );
  BUFX2 U1617 ( .A(n2867), .Y(n2024) );
  INVX1 U1618 ( .A(n2875), .Y(n2025) );
  INVX1 U1619 ( .A(n2025), .Y(n2026) );
  BUFX2 U1620 ( .A(n2897), .Y(n2027) );
  INVX1 U1621 ( .A(n2900), .Y(n2028) );
  INVX1 U1622 ( .A(n2028), .Y(n2029) );
  BUFX2 U1623 ( .A(n2904), .Y(n2030) );
  BUFX2 U1624 ( .A(n2907), .Y(n2031) );
  BUFX2 U1625 ( .A(n2910), .Y(n2032) );
  BUFX2 U1626 ( .A(n2913), .Y(n2033) );
  BUFX2 U1627 ( .A(n2917), .Y(n2034) );
  BUFX2 U1628 ( .A(n2920), .Y(n2035) );
  BUFX2 U1629 ( .A(n2673), .Y(n2036) );
  BUFX2 U1630 ( .A(n2680), .Y(n2037) );
  BUFX2 U1631 ( .A(n1410), .Y(n2038) );
  BUFX2 U1632 ( .A(n1409), .Y(n2039) );
  BUFX2 U1633 ( .A(n1181), .Y(n2040) );
  BUFX2 U1634 ( .A(n1178), .Y(n2041) );
  INVX1 U1635 ( .A(n2608), .Y(n2042) );
  AND2X1 U1636 ( .A(n2503), .B(WB_data[56]), .Y(n2609) );
  INVX1 U1637 ( .A(n2609), .Y(n2043) );
  AND2X1 U1638 ( .A(n2505), .B(WB_data[54]), .Y(n2613) );
  INVX1 U1639 ( .A(n2613), .Y(n2044) );
  AND2X1 U1640 ( .A(n2505), .B(WB_data[53]), .Y(n2614) );
  INVX1 U1641 ( .A(n2614), .Y(n2045) );
  AND2X1 U1642 ( .A(n2505), .B(WB_data[52]), .Y(n2615) );
  INVX1 U1643 ( .A(n2615), .Y(n2046) );
  INVX1 U1644 ( .A(n2621), .Y(n2047) );
  AND2X1 U1645 ( .A(n2503), .B(WB_data[46]), .Y(n2622) );
  INVX1 U1646 ( .A(n2622), .Y(n2048) );
  AND2X1 U1647 ( .A(n2503), .B(WB_data[45]), .Y(n2623) );
  INVX1 U1648 ( .A(n2623), .Y(n2049) );
  AND2X1 U1649 ( .A(n2503), .B(WB_data[44]), .Y(n2624) );
  INVX1 U1650 ( .A(n2624), .Y(n2050) );
  AND2X2 U1651 ( .A(n2503), .B(WB_data[42]), .Y(n2626) );
  INVX1 U1652 ( .A(n2626), .Y(n2051) );
  INVX1 U1653 ( .A(n2632), .Y(n2052) );
  AND2X1 U1654 ( .A(n2505), .B(n2519), .Y(n2635) );
  INVX1 U1655 ( .A(n2635), .Y(n2053) );
  AND2X1 U1656 ( .A(n2505), .B(n2258), .Y(n2638) );
  INVX1 U1657 ( .A(n2638), .Y(n2054) );
  INVX1 U1658 ( .A(n2641), .Y(n2055) );
  INVX1 U1659 ( .A(n2644), .Y(n2056) );
  INVX1 U1660 ( .A(n2647), .Y(n2057) );
  AND2X2 U1661 ( .A(n2505), .B(n2205), .Y(n2650) );
  INVX1 U1662 ( .A(n2650), .Y(n2058) );
  AND2X1 U1663 ( .A(EX_oprB[29]), .B(n2484), .Y(n2663) );
  INVX1 U1664 ( .A(n2663), .Y(n2059) );
  AND2X1 U1665 ( .A(EX_oprB[26]), .B(n2484), .Y(n2675) );
  INVX1 U1666 ( .A(n2675), .Y(n2060) );
  INVX1 U1667 ( .A(n2690), .Y(n2061) );
  AND2X1 U1668 ( .A(n2504), .B(WB_data[18]), .Y(n2701) );
  INVX1 U1669 ( .A(n2701), .Y(n2062) );
  INVX1 U1670 ( .A(n2710), .Y(n2063) );
  INVX1 U1671 ( .A(n2712), .Y(n2064) );
  INVX1 U1672 ( .A(n2713), .Y(n2065) );
  INVX1 U1673 ( .A(n2714), .Y(n2066) );
  INVX1 U1674 ( .A(n2717), .Y(n2067) );
  INVX1 U1675 ( .A(n2735), .Y(n2068) );
  INVX1 U1676 ( .A(n2745), .Y(n2069) );
  INVX1 U1677 ( .A(n2069), .Y(n2070) );
  BUFX2 U1678 ( .A(n1402), .Y(n2071) );
  BUFX2 U1679 ( .A(n1401), .Y(n2072) );
  AND2X1 U1680 ( .A(n2506), .B(ID_instruction[2]), .Y(n1187) );
  INVX1 U1681 ( .A(n1187), .Y(n2073) );
  BUFX2 U1682 ( .A(n3279), .Y(n2074) );
  INVX1 U1683 ( .A(n2802), .Y(n2075) );
  INVX1 U1684 ( .A(n2795), .Y(n2076) );
  INVX1 U1685 ( .A(n2076), .Y(n2077) );
  BUFX2 U1686 ( .A(n2769), .Y(n2078) );
  BUFX2 U1687 ( .A(n2871), .Y(n2079) );
  BUFX2 U1688 ( .A(n2927), .Y(n2080) );
  AND2X1 U1689 ( .A(n2475), .B(n2606), .Y(n2768) );
  INVX1 U1690 ( .A(n2768), .Y(n2081) );
  INVX1 U1691 ( .A(n2926), .Y(n2082) );
  OR2X1 U1692 ( .A(dataOut[39]), .B(dataOut[38]), .Y(n2966) );
  INVX1 U1693 ( .A(n2966), .Y(n2083) );
  OR2X1 U1694 ( .A(dataOut[47]), .B(dataOut[46]), .Y(n2970) );
  INVX1 U1695 ( .A(n2970), .Y(n2084) );
  OR2X1 U1696 ( .A(dataOut[55]), .B(dataOut[54]), .Y(n2978) );
  INVX1 U1697 ( .A(n2978), .Y(n2085) );
  OR2X1 U1698 ( .A(dataOut[51]), .B(dataOut[50]), .Y(n2979) );
  INVX1 U1699 ( .A(n2979), .Y(n2086) );
  OR2X1 U1700 ( .A(dataOut[31]), .B(dataOut[30]), .Y(n2988) );
  INVX1 U1701 ( .A(n2988), .Y(n2087) );
  AND2X1 U1702 ( .A(instruction[2]), .B(n1920), .Y(n1188) );
  INVX1 U1703 ( .A(n1188), .Y(n2088) );
  BUFX2 U1704 ( .A(n2969), .Y(n2089) );
  BUFX2 U1705 ( .A(n2973), .Y(n2090) );
  BUFX2 U1706 ( .A(n3006), .Y(n2091) );
  BUFX2 U1707 ( .A(n2991), .Y(n2092) );
  BUFX2 U1708 ( .A(n2981), .Y(n2093) );
  BUFX2 U1709 ( .A(n3005), .Y(n2094) );
  BUFX2 U1710 ( .A(n1404), .Y(n2095) );
  AND2X1 U1711 ( .A(n3076), .B(n3074), .Y(n2968) );
  INVX1 U1712 ( .A(n2968), .Y(n2096) );
  AND2X1 U1713 ( .A(n3060), .B(n3058), .Y(n2972) );
  INVX1 U1714 ( .A(n2972), .Y(n2097) );
  AND2X1 U1715 ( .A(n3092), .B(n3090), .Y(n2990) );
  INVX1 U1716 ( .A(n2990), .Y(n2098) );
  BUFX2 U1717 ( .A(n2980), .Y(n2099) );
  BUFX2 U1718 ( .A(n3004), .Y(n2100) );
  AND2X1 U1719 ( .A(n3080), .B(n3078), .Y(n2967) );
  INVX1 U1720 ( .A(n2967), .Y(n2101) );
  AND2X1 U1721 ( .A(n3064), .B(n3062), .Y(n2971) );
  INVX1 U1722 ( .A(n2971), .Y(n2102) );
  AND2X1 U1723 ( .A(n3096), .B(n3094), .Y(n2989) );
  INVX1 U1724 ( .A(n2989), .Y(n2103) );
  INVX1 U1725 ( .A(n2746), .Y(n2104) );
  INVX1 U1726 ( .A(n2104), .Y(n2105) );
  INVX1 U1727 ( .A(n3270), .Y(n2106) );
  INVX1 U1728 ( .A(n1953), .Y(n2107) );
  INVX1 U1729 ( .A(n2109), .Y(n2108) );
  AND2X2 U1730 ( .A(n2489), .B(n2111), .Y(n2869) );
  INVX1 U1731 ( .A(n2869), .Y(n2109) );
  INVX1 U1732 ( .A(n2853), .Y(n2110) );
  INVX1 U1733 ( .A(n2110), .Y(n2111) );
  BUFX2 U1734 ( .A(n2878), .Y(n2112) );
  INVX1 U1735 ( .A(n2114), .Y(n2113) );
  BUFX2 U1736 ( .A(n2688), .Y(n2114) );
  INVX1 U1737 ( .A(n2116), .Y(n2115) );
  BUFX2 U1738 ( .A(n2695), .Y(n2116) );
  AND2X2 U1739 ( .A(n2511), .B(n1998), .Y(n2505) );
  INVX1 U1740 ( .A(n2780), .Y(n2117) );
  INVX1 U1741 ( .A(n2117), .Y(n2118) );
  INVX1 U1742 ( .A(n2792), .Y(n2119) );
  INVX1 U1743 ( .A(n2119), .Y(n2120) );
  INVX1 U1744 ( .A(n2800), .Y(n2121) );
  INVX1 U1745 ( .A(n2121), .Y(n2122) );
  INVX1 U1746 ( .A(n2805), .Y(n2123) );
  INVX1 U1747 ( .A(n2123), .Y(n2124) );
  INVX1 U1748 ( .A(n2126), .Y(n2125) );
  BUFX2 U1749 ( .A(n2958), .Y(n2126) );
  BUFX2 U1750 ( .A(n2781), .Y(n2127) );
  INVX1 U1751 ( .A(n1991), .Y(n2128) );
  INVX1 U1752 ( .A(n1991), .Y(n2129) );
  INVX1 U1753 ( .A(n2689), .Y(n2130) );
  INVX1 U1754 ( .A(n2130), .Y(n2131) );
  BUFX2 U1755 ( .A(n2777), .Y(n2132) );
  AND2X2 U1756 ( .A(n2566), .B(n2580), .Y(n2516) );
  AND2X1 U1757 ( .A(instruction[31]), .B(n2557), .Y(n1249) );
  INVX1 U1758 ( .A(n1249), .Y(n2136) );
  AND2X1 U1759 ( .A(EX_oprA[1]), .B(n2506), .Y(n3141) );
  INVX1 U1760 ( .A(n3141), .Y(n2137) );
  AND2X1 U1761 ( .A(ID_oprB[20]), .B(n2558), .Y(n3187) );
  INVX1 U1762 ( .A(n3187), .Y(n2138) );
  AND2X1 U1763 ( .A(ID_oprB[61]), .B(n2500), .Y(n3268) );
  INVX1 U1764 ( .A(n3268), .Y(n2139) );
  AND2X1 U1765 ( .A(ID_oprB[31]), .B(n2557), .Y(n3208) );
  INVX1 U1766 ( .A(n3208), .Y(n2140) );
  AND2X1 U1767 ( .A(instruction[21]), .B(n2500), .Y(n1231) );
  INVX1 U1768 ( .A(n1231), .Y(n2141) );
  AND2X1 U1769 ( .A(EX_oprA[2]), .B(n2506), .Y(n3139) );
  INVX1 U1770 ( .A(n3139), .Y(n2142) );
  AND2X1 U1771 ( .A(EX_oprA[17]), .B(n2506), .Y(n3109) );
  INVX1 U1772 ( .A(n3109), .Y(n2143) );
  AND2X1 U1773 ( .A(EX_oprA[30]), .B(n2506), .Y(n3083) );
  INVX1 U1774 ( .A(n3083), .Y(n2144) );
  AND2X1 U1775 ( .A(EX_oprA[45]), .B(n2506), .Y(n3053) );
  INVX1 U1776 ( .A(n3053), .Y(n2145) );
  AND2X1 U1777 ( .A(EX_shift_amt[0]), .B(n2506), .Y(n1213) );
  INVX1 U1778 ( .A(n1213), .Y(n2146) );
  AND2X1 U1779 ( .A(ID_oprB[49]), .B(n2557), .Y(n3244) );
  INVX1 U1780 ( .A(n3244), .Y(n2147) );
  AND2X1 U1781 ( .A(ID_oprB[19]), .B(n2558), .Y(n3185) );
  INVX1 U1782 ( .A(n3185), .Y(n2148) );
  INVX1 U1783 ( .A(WB_data[39]), .Y(n2149) );
  AND2X1 U1784 ( .A(n2562), .B(WB_mult32_result[39]), .Y(n2630) );
  INVX1 U1785 ( .A(n2630), .Y(n2150) );
  BUFX2 U1786 ( .A(n2631), .Y(n2151) );
  AND2X1 U1787 ( .A(ID_oprB[60]), .B(n2500), .Y(n3266) );
  INVX1 U1788 ( .A(n3266), .Y(n2152) );
  AND2X1 U1789 ( .A(ID_oprB[30]), .B(n2558), .Y(n3206) );
  INVX1 U1790 ( .A(n3206), .Y(n2153) );
  AND2X1 U1791 ( .A(instruction[20]), .B(n2500), .Y(n1227) );
  INVX1 U1792 ( .A(n1227), .Y(n2154) );
  AND2X1 U1793 ( .A(EX_oprA[3]), .B(n2506), .Y(n3137) );
  INVX1 U1794 ( .A(n3137), .Y(n2155) );
  AND2X1 U1795 ( .A(EX_oprA[18]), .B(n2506), .Y(n3107) );
  INVX1 U1796 ( .A(n3107), .Y(n2156) );
  AND2X1 U1797 ( .A(EX_oprA[31]), .B(n2506), .Y(n3081) );
  INVX1 U1798 ( .A(n3081), .Y(n2157) );
  AND2X1 U1799 ( .A(EX_oprA[46]), .B(n2506), .Y(n3051) );
  INVX1 U1800 ( .A(n3051), .Y(n2158) );
  AND2X1 U1801 ( .A(EX_shift_amt[1]), .B(n2506), .Y(n1214) );
  INVX1 U1802 ( .A(n1214), .Y(n2159) );
  AND2X1 U1803 ( .A(ID_oprB[48]), .B(n2557), .Y(n3242) );
  INVX1 U1804 ( .A(n3242), .Y(n2160) );
  AND2X1 U1805 ( .A(ID_oprB[16]), .B(n2558), .Y(n3179) );
  INVX1 U1806 ( .A(n3179), .Y(n2161) );
  INVX1 U1807 ( .A(WB_data[35]), .Y(n2162) );
  BUFX2 U1808 ( .A(n2643), .Y(n2163) );
  AND2X1 U1809 ( .A(WB_mult32_result[35]), .B(n2562), .Y(n2642) );
  INVX1 U1810 ( .A(n2642), .Y(n2164) );
  AND2X1 U1811 ( .A(ID_oprB[59]), .B(n2500), .Y(n3264) );
  INVX1 U1812 ( .A(n3264), .Y(n2165) );
  AND2X1 U1813 ( .A(ID_oprB[29]), .B(n2557), .Y(n3204) );
  INVX1 U1814 ( .A(n3204), .Y(n2166) );
  AND2X1 U1815 ( .A(instruction[19]), .B(n2500), .Y(n1225) );
  INVX1 U1816 ( .A(n1225), .Y(n2167) );
  AND2X1 U1817 ( .A(EX_oprA[4]), .B(n2506), .Y(n3135) );
  INVX1 U1818 ( .A(n3135), .Y(n2168) );
  AND2X1 U1819 ( .A(EX_oprA[19]), .B(n2506), .Y(n3105) );
  INVX1 U1820 ( .A(n3105), .Y(n2169) );
  AND2X1 U1821 ( .A(EX_oprA[32]), .B(n2506), .Y(n3079) );
  INVX1 U1822 ( .A(n3079), .Y(n2170) );
  AND2X1 U1823 ( .A(EX_oprA[47]), .B(n2506), .Y(n3049) );
  INVX1 U1824 ( .A(n3049), .Y(n2171) );
  AND2X1 U1825 ( .A(EX_shift_amt[2]), .B(n2506), .Y(n1215) );
  INVX1 U1826 ( .A(n1215), .Y(n2172) );
  AND2X1 U1827 ( .A(ID_oprB[47]), .B(n2557), .Y(n3240) );
  INVX1 U1828 ( .A(n3240), .Y(n2173) );
  AND2X1 U1829 ( .A(ID_oprB[15]), .B(n2558), .Y(n3177) );
  INVX1 U1830 ( .A(n3177), .Y(n2174) );
  BUFX2 U1831 ( .A(n2905), .Y(n2175) );
  AND2X2 U1832 ( .A(n2178), .B(n2179), .Y(WB_data[19]) );
  INVX1 U1833 ( .A(WB_data[19]), .Y(n2176) );
  INVX1 U1834 ( .A(WB_data[19]), .Y(n2177) );
  BUFX2 U1835 ( .A(n2699), .Y(n2178) );
  AND2X1 U1836 ( .A(WB_mult32_result[19]), .B(n2562), .Y(n2698) );
  INVX1 U1837 ( .A(n2698), .Y(n2179) );
  AND2X1 U1838 ( .A(ID_oprB[58]), .B(n2500), .Y(n3262) );
  INVX1 U1839 ( .A(n3262), .Y(n2180) );
  AND2X1 U1840 ( .A(ID_oprB[28]), .B(n2558), .Y(n3202) );
  INVX1 U1841 ( .A(n3202), .Y(n2181) );
  AND2X1 U1842 ( .A(instruction[18]), .B(n2500), .Y(n1223) );
  INVX1 U1843 ( .A(n1223), .Y(n2182) );
  AND2X1 U1844 ( .A(EX_oprA[5]), .B(n2506), .Y(n3133) );
  INVX1 U1845 ( .A(n3133), .Y(n2183) );
  AND2X1 U1846 ( .A(EX_oprA[20]), .B(n2506), .Y(n3103) );
  INVX1 U1847 ( .A(n3103), .Y(n2184) );
  AND2X1 U1848 ( .A(EX_oprA[33]), .B(n2506), .Y(n3077) );
  INVX1 U1849 ( .A(n3077), .Y(n2185) );
  AND2X1 U1850 ( .A(EX_oprA[48]), .B(n2506), .Y(n3047) );
  INVX1 U1851 ( .A(n3047), .Y(n2186) );
  AND2X1 U1852 ( .A(EX_shift_amt[3]), .B(n2506), .Y(n1216) );
  INVX1 U1853 ( .A(n1216), .Y(n2187) );
  AND2X1 U1854 ( .A(ID_oprB[42]), .B(n2557), .Y(n3230) );
  INVX1 U1855 ( .A(n3230), .Y(n2188) );
  AND2X1 U1856 ( .A(ID_oprB[14]), .B(n2558), .Y(n3175) );
  INVX1 U1857 ( .A(n3175), .Y(n2189) );
  BUFX2 U1858 ( .A(n2915), .Y(n2190) );
  AND2X2 U1859 ( .A(n2192), .B(n2193), .Y(WB_data[36]) );
  BUFX2 U1860 ( .A(n2640), .Y(n2192) );
  AND2X1 U1861 ( .A(WB_mult32_result[36]), .B(n2562), .Y(n2639) );
  INVX1 U1862 ( .A(n2639), .Y(n2193) );
  AND2X1 U1863 ( .A(ID_oprB[25]), .B(n2557), .Y(n3197) );
  INVX1 U1864 ( .A(n3197), .Y(n2194) );
  AND2X1 U1865 ( .A(instruction[17]), .B(n2500), .Y(n1221) );
  INVX1 U1866 ( .A(n1221), .Y(n2195) );
  AND2X1 U1867 ( .A(instruction[5]), .B(n2500), .Y(n1191) );
  INVX1 U1868 ( .A(n1191), .Y(n2196) );
  AND2X1 U1869 ( .A(EX_oprA[6]), .B(n2506), .Y(n3131) );
  INVX1 U1870 ( .A(n3131), .Y(n2197) );
  AND2X1 U1871 ( .A(EX_oprA[21]), .B(n2506), .Y(n3101) );
  INVX1 U1872 ( .A(n3101), .Y(n2198) );
  AND2X1 U1873 ( .A(EX_oprA[34]), .B(n2506), .Y(n3075) );
  INVX1 U1874 ( .A(n3075), .Y(n2199) );
  AND2X1 U1875 ( .A(EX_oprA[49]), .B(n2506), .Y(n3045) );
  INVX1 U1876 ( .A(n3045), .Y(n2200) );
  AND2X1 U1877 ( .A(EX_PPP[0]), .B(n2506), .Y(n1228) );
  INVX1 U1878 ( .A(n1228), .Y(n2201) );
  AND2X1 U1879 ( .A(ID_oprB[41]), .B(n2557), .Y(n3228) );
  INVX1 U1880 ( .A(n3228), .Y(n2202) );
  AND2X1 U1881 ( .A(ID_oprB[13]), .B(n2558), .Y(n3173) );
  INVX1 U1882 ( .A(n3173), .Y(n2203) );
  BUFX2 U1883 ( .A(n2918), .Y(n2204) );
  INVX1 U1884 ( .A(WB_data[33]), .Y(n2205) );
  BUFX2 U1885 ( .A(n2649), .Y(n2206) );
  AND2X1 U1886 ( .A(WB_mult32_result[33]), .B(n2562), .Y(n2648) );
  INVX1 U1887 ( .A(n2648), .Y(n2207) );
  AND2X1 U1888 ( .A(instruction[30]), .B(n2558), .Y(n1248) );
  INVX1 U1889 ( .A(n1248), .Y(n2208) );
  AND2X1 U1890 ( .A(instruction[16]), .B(n2500), .Y(n1219) );
  INVX1 U1891 ( .A(n1219), .Y(n2209) );
  AND2X1 U1892 ( .A(instruction[4]), .B(n2500), .Y(n1190) );
  INVX1 U1893 ( .A(n1190), .Y(n2210) );
  AND2X1 U1894 ( .A(EX_oprA[8]), .B(n2506), .Y(n3127) );
  INVX1 U1895 ( .A(n3127), .Y(n2211) );
  AND2X1 U1896 ( .A(EX_oprA[22]), .B(n2506), .Y(n3099) );
  INVX1 U1897 ( .A(n3099), .Y(n2212) );
  AND2X1 U1898 ( .A(EX_oprA[35]), .B(n2506), .Y(n3073) );
  INVX1 U1899 ( .A(n3073), .Y(n2213) );
  AND2X1 U1900 ( .A(EX_oprA[50]), .B(n2506), .Y(n3043) );
  INVX1 U1901 ( .A(n3043), .Y(n2214) );
  AND2X1 U1902 ( .A(EX_PPP[1]), .B(n2506), .Y(n1229) );
  INVX1 U1903 ( .A(n1229), .Y(n2215) );
  AND2X1 U1904 ( .A(ID_oprB[46]), .B(n2557), .Y(n3238) );
  INVX1 U1905 ( .A(n3238), .Y(n2216) );
  AND2X1 U1906 ( .A(ID_oprB[35]), .B(n2557), .Y(n3216) );
  INVX1 U1907 ( .A(n3216), .Y(n2217) );
  AND2X1 U1908 ( .A(ID_oprB[12]), .B(n2558), .Y(n3171) );
  INVX1 U1909 ( .A(n3171), .Y(n2218) );
  AND2X2 U1910 ( .A(n2221), .B(n2222), .Y(WB_data[4]) );
  INVX1 U1911 ( .A(WB_data[4]), .Y(n2219) );
  INVX1 U1912 ( .A(n1931), .Y(n2220) );
  BUFX2 U1913 ( .A(n2725), .Y(n2221) );
  AND2X1 U1914 ( .A(WB_mult32_result[4]), .B(n2562), .Y(n2724) );
  INVX1 U1915 ( .A(n2724), .Y(n2222) );
  AND2X1 U1916 ( .A(instruction[29]), .B(n2500), .Y(n1247) );
  INVX1 U1917 ( .A(n1247), .Y(n2223) );
  AND2X1 U1918 ( .A(instruction[14]), .B(n2500), .Y(n1210) );
  INVX1 U1919 ( .A(n1210), .Y(n2224) );
  AND2X1 U1920 ( .A(EX_oprA[9]), .B(n2506), .Y(n3125) );
  INVX1 U1921 ( .A(n3125), .Y(n2225) );
  AND2X1 U1922 ( .A(EX_oprA[23]), .B(n2506), .Y(n3097) );
  INVX1 U1923 ( .A(n3097), .Y(n2226) );
  AND2X1 U1924 ( .A(EX_oprA[36]), .B(n2506), .Y(n3071) );
  INVX1 U1925 ( .A(n3071), .Y(n2227) );
  AND2X1 U1926 ( .A(EX_oprA[51]), .B(n2506), .Y(n3041) );
  INVX1 U1927 ( .A(n3041), .Y(n2228) );
  AND2X1 U1928 ( .A(n2506), .B(EX_dest_reg[0]), .Y(n1192) );
  INVX1 U1929 ( .A(n1192), .Y(n2229) );
  AND2X1 U1930 ( .A(EX_PPP[2]), .B(n2506), .Y(n1230) );
  INVX1 U1931 ( .A(n1230), .Y(n2230) );
  AND2X1 U1932 ( .A(ID_oprB[57]), .B(n2500), .Y(n3260) );
  INVX1 U1933 ( .A(n3260), .Y(n2231) );
  AND2X1 U1934 ( .A(ID_oprB[45]), .B(n2557), .Y(n3236) );
  INVX1 U1935 ( .A(n3236), .Y(n2232) );
  AND2X1 U1936 ( .A(ID_oprB[34]), .B(n2558), .Y(n3214) );
  INVX1 U1937 ( .A(n3214), .Y(n2233) );
  AND2X1 U1938 ( .A(ID_oprB[11]), .B(n2558), .Y(n3169) );
  INVX1 U1939 ( .A(n3169), .Y(n2234) );
  BUFX2 U1940 ( .A(n2839), .Y(n2235) );
  BUFX2 U1941 ( .A(n2831), .Y(n2236) );
  BUFX2 U1942 ( .A(n2895), .Y(n2237) );
  AND2X2 U1943 ( .A(n2239), .B(n2240), .Y(WB_data[34]) );
  BUFX2 U1944 ( .A(n2646), .Y(n2239) );
  AND2X1 U1945 ( .A(WB_mult32_result[34]), .B(n2562), .Y(n2645) );
  INVX1 U1946 ( .A(n2645), .Y(n2240) );
  AND2X1 U1947 ( .A(n1202), .B(n1313), .Y(n1312) );
  INVX1 U1948 ( .A(n1312), .Y(n2241) );
  AND2X1 U1949 ( .A(instruction[28]), .B(n2500), .Y(n1246) );
  INVX1 U1950 ( .A(n1246), .Y(n2242) );
  AND2X1 U1951 ( .A(instruction[13]), .B(n2500), .Y(n1208) );
  INVX1 U1952 ( .A(n1208), .Y(n2243) );
  AND2X1 U1953 ( .A(ID_oprB[63]), .B(n2558), .Y(n3145) );
  INVX1 U1954 ( .A(n3145), .Y(n2244) );
  AND2X1 U1955 ( .A(EX_oprA[10]), .B(n2506), .Y(n3123) );
  INVX1 U1956 ( .A(n3123), .Y(n2245) );
  AND2X1 U1957 ( .A(EX_oprA[24]), .B(n2506), .Y(n3095) );
  INVX1 U1958 ( .A(n3095), .Y(n2246) );
  AND2X1 U1959 ( .A(EX_oprA[37]), .B(n2506), .Y(n3069) );
  INVX1 U1960 ( .A(n3069), .Y(n2247) );
  AND2X1 U1961 ( .A(EX_oprA[54]), .B(n2506), .Y(n3035) );
  INVX1 U1962 ( .A(n3035), .Y(n2248) );
  AND2X1 U1963 ( .A(n2506), .B(EX_dest_reg[2]), .Y(n1194) );
  INVX1 U1964 ( .A(n1194), .Y(n2249) );
  AND2X1 U1965 ( .A(EX_WW[0]), .B(n2506), .Y(n1234) );
  INVX1 U1966 ( .A(n1234), .Y(n2250) );
  AND2X1 U1967 ( .A(ID_oprB[54]), .B(n2500), .Y(n3254) );
  INVX1 U1968 ( .A(n3254), .Y(n2251) );
  AND2X1 U1969 ( .A(ID_oprB[40]), .B(n2557), .Y(n3226) );
  INVX1 U1970 ( .A(n3226), .Y(n2252) );
  AND2X1 U1971 ( .A(ID_oprB[27]), .B(n2558), .Y(n3200) );
  INVX1 U1972 ( .A(n3200), .Y(n2253) );
  AND2X1 U1973 ( .A(ID_oprB[10]), .B(n2558), .Y(n3167) );
  INVX1 U1974 ( .A(n3167), .Y(n2254) );
  BUFX2 U1975 ( .A(n2810), .Y(n2255) );
  BUFX2 U1976 ( .A(n2835), .Y(n2256) );
  BUFX2 U1977 ( .A(n2911), .Y(n2257) );
  AND2X2 U1978 ( .A(n2259), .B(n2260), .Y(WB_data[37]) );
  BUFX2 U1979 ( .A(n2637), .Y(n2259) );
  AND2X1 U1980 ( .A(WB_mult32_result[37]), .B(n2562), .Y(n2636) );
  INVX1 U1981 ( .A(n2636), .Y(n2260) );
  AND2X1 U1982 ( .A(instruction[26]), .B(n2558), .Y(n1244) );
  INVX1 U1983 ( .A(n1244), .Y(n2261) );
  AND2X1 U1984 ( .A(instruction[12]), .B(n2500), .Y(n1206) );
  INVX1 U1985 ( .A(n1206), .Y(n2262) );
  AND2X1 U1986 ( .A(EX_oprA[11]), .B(n2506), .Y(n3121) );
  INVX1 U1987 ( .A(n3121), .Y(n2263) );
  AND2X1 U1988 ( .A(EX_oprA[25]), .B(n2506), .Y(n3093) );
  INVX1 U1989 ( .A(n3093), .Y(n2264) );
  AND2X1 U1990 ( .A(EX_oprA[38]), .B(n2506), .Y(n3067) );
  INVX1 U1991 ( .A(n3067), .Y(n2265) );
  AND2X1 U1992 ( .A(EX_oprA[55]), .B(n2506), .Y(n3033) );
  INVX1 U1993 ( .A(n3033), .Y(n2266) );
  AND2X1 U1994 ( .A(EX_oprA[63]), .B(n2506), .Y(n3017) );
  INVX1 U1995 ( .A(n3017), .Y(n2267) );
  AND2X1 U1996 ( .A(EX_WW[1]), .B(n2506), .Y(n1235) );
  INVX1 U1997 ( .A(n1235), .Y(n2268) );
  AND2X1 U1998 ( .A(ID_oprB[53]), .B(n2500), .Y(n3252) );
  INVX1 U1999 ( .A(n3252), .Y(n2269) );
  AND2X1 U2000 ( .A(ID_oprB[39]), .B(n2557), .Y(n3224) );
  INVX1 U2001 ( .A(n3224), .Y(n2270) );
  AND2X1 U2002 ( .A(ID_oprB[24]), .B(n2557), .Y(n3195) );
  INVX1 U2003 ( .A(n3195), .Y(n2271) );
  AND2X1 U2004 ( .A(ID_oprB[9]), .B(n2558), .Y(n3165) );
  INVX1 U2005 ( .A(n3165), .Y(n2272) );
  AND2X1 U2006 ( .A(ID_oprB[3]), .B(n2557), .Y(n3153) );
  INVX1 U2007 ( .A(n3153), .Y(n2273) );
  BUFX2 U2008 ( .A(n2893), .Y(n2274) );
  INVX1 U2009 ( .A(n2892), .Y(n2275) );
  BUFX2 U2010 ( .A(n2873), .Y(n2276) );
  BUFX2 U2011 ( .A(n2806), .Y(n2277) );
  BUFX2 U2012 ( .A(n2939), .Y(n2278) );
  BUFX2 U2013 ( .A(n2935), .Y(n2279) );
  INVX1 U2014 ( .A(WB_data[5]), .Y(n2281) );
  BUFX2 U2015 ( .A(n2722), .Y(n2282) );
  AND2X1 U2016 ( .A(WB_mult32_result[5]), .B(n2562), .Y(n2721) );
  INVX1 U2017 ( .A(n2721), .Y(n2283) );
  AND2X1 U2018 ( .A(instruction[27]), .B(n2557), .Y(n1245) );
  INVX1 U2019 ( .A(n1245), .Y(n2284) );
  AND2X1 U2020 ( .A(instruction[10]), .B(n2500), .Y(n1201) );
  INVX1 U2021 ( .A(n1201), .Y(n2285) );
  AND2X1 U2022 ( .A(EX_oprA[12]), .B(n2506), .Y(n3119) );
  INVX1 U2023 ( .A(n3119), .Y(n2286) );
  AND2X1 U2024 ( .A(EX_oprA[26]), .B(n2506), .Y(n3091) );
  INVX1 U2025 ( .A(n3091), .Y(n2287) );
  AND2X1 U2026 ( .A(EX_oprA[42]), .B(n2506), .Y(n3059) );
  INVX1 U2027 ( .A(n3059), .Y(n2288) );
  AND2X1 U2028 ( .A(EX_oprA[57]), .B(n2506), .Y(n3029) );
  INVX1 U2029 ( .A(n3029), .Y(n2289) );
  AND2X1 U2030 ( .A(EX_alu_func[0]), .B(n2506), .Y(n1238) );
  INVX1 U2031 ( .A(n1238), .Y(n2290) );
  AND2X1 U2032 ( .A(ID_oprB[52]), .B(n2500), .Y(n3250) );
  INVX1 U2033 ( .A(n3250), .Y(n2291) );
  AND2X1 U2034 ( .A(ID_oprB[38]), .B(n2557), .Y(n3222) );
  INVX1 U2035 ( .A(n3222), .Y(n2292) );
  AND2X1 U2036 ( .A(ID_oprB[23]), .B(n2558), .Y(n3193) );
  INVX1 U2037 ( .A(n3193), .Y(n2293) );
  AND2X1 U2038 ( .A(ID_oprB[8]), .B(n2558), .Y(n3163) );
  INVX1 U2039 ( .A(n3163), .Y(n2294) );
  AND2X1 U2040 ( .A(ID_oprB[2]), .B(n2558), .Y(n3151) );
  INVX1 U2041 ( .A(n3151), .Y(n2295) );
  AND2X1 U2042 ( .A(n1313), .B(ID_instruction[11]), .Y(n1400) );
  INVX1 U2043 ( .A(n1400), .Y(n2296) );
  BUFX2 U2044 ( .A(n1362), .Y(n2297) );
  BUFX2 U2045 ( .A(n1363), .Y(n2298) );
  BUFX2 U2046 ( .A(n2908), .Y(n2299) );
  BUFX2 U2047 ( .A(n2816), .Y(n2300) );
  BUFX2 U2048 ( .A(n2954), .Y(n2301) );
  INVX1 U2049 ( .A(WB_data[17]), .Y(n2302) );
  INVX1 U2050 ( .A(WB_data[17]), .Y(n2303) );
  BUFX2 U2051 ( .A(n2703), .Y(n2304) );
  AND2X1 U2052 ( .A(WB_mult32_result[17]), .B(n2562), .Y(n2702) );
  INVX1 U2053 ( .A(n2702), .Y(n2305) );
  AND2X1 U2054 ( .A(instruction[25]), .B(n2558), .Y(n1237) );
  INVX1 U2055 ( .A(n1237), .Y(n2306) );
  AND2X1 U2056 ( .A(instruction[11]), .B(n2500), .Y(n1204) );
  INVX1 U2057 ( .A(n1204), .Y(n2307) );
  AND2X1 U2058 ( .A(EX_oprA[13]), .B(n2506), .Y(n3117) );
  INVX1 U2059 ( .A(n3117), .Y(n2308) );
  AND2X1 U2060 ( .A(EX_oprA[27]), .B(n2506), .Y(n3089) );
  INVX1 U2061 ( .A(n3089), .Y(n2309) );
  AND2X1 U2062 ( .A(EX_oprA[43]), .B(n2506), .Y(n3057) );
  INVX1 U2063 ( .A(n3057), .Y(n2310) );
  AND2X1 U2064 ( .A(EX_oprA[58]), .B(n2506), .Y(n3027) );
  INVX1 U2065 ( .A(n3027), .Y(n2311) );
  AND2X1 U2066 ( .A(n2506), .B(EX_dest_reg[3]), .Y(n1195) );
  INVX1 U2067 ( .A(n1195), .Y(n2312) );
  AND2X1 U2068 ( .A(EX_alu_func[1]), .B(n2506), .Y(n1239) );
  INVX1 U2069 ( .A(n1239), .Y(n2313) );
  AND2X1 U2070 ( .A(ID_oprB[56]), .B(n2500), .Y(n3258) );
  INVX1 U2071 ( .A(n3258), .Y(n2314) );
  AND2X1 U2072 ( .A(ID_oprB[44]), .B(n2557), .Y(n3234) );
  INVX1 U2073 ( .A(n3234), .Y(n2315) );
  AND2X1 U2074 ( .A(ID_oprB[33]), .B(n2557), .Y(n3212) );
  INVX1 U2075 ( .A(n3212), .Y(n2316) );
  AND2X1 U2076 ( .A(ID_oprB[18]), .B(n2558), .Y(n3183) );
  INVX1 U2077 ( .A(n3183), .Y(n2317) );
  AND2X1 U2078 ( .A(ID_oprB[5]), .B(n2558), .Y(n3157) );
  INVX1 U2079 ( .A(n3157), .Y(n2318) );
  AND2X1 U2080 ( .A(n1313), .B(ID_instruction[15]), .Y(n1396) );
  INVX1 U2081 ( .A(n1396), .Y(n2319) );
  BUFX2 U2082 ( .A(n2757), .Y(n2320) );
  INVX1 U2083 ( .A(n1789), .Y(n2321) );
  AND2X1 U2084 ( .A(instruction[1]), .B(n2554), .Y(n1186) );
  INVX1 U2085 ( .A(n1186), .Y(n2322) );
  AND2X1 U2086 ( .A(n3302), .B(n3301), .Y(n1395) );
  INVX1 U2087 ( .A(n1395), .Y(n2323) );
  AND2X1 U2088 ( .A(n3140), .B(n3138), .Y(n2995) );
  INVX1 U2089 ( .A(n2995), .Y(n2324) );
  AND2X1 U2090 ( .A(n3272), .B(n2370), .Y(memWrEn) );
  INVX1 U2091 ( .A(memWrEn), .Y(n2325) );
  BUFX2 U2092 ( .A(n2827), .Y(n2326) );
  BUFX2 U2093 ( .A(n2902), .Y(n2327) );
  BUFX2 U2094 ( .A(n2949), .Y(n2328) );
  BUFX2 U2095 ( .A(n2925), .Y(n2329) );
  INVX1 U2096 ( .A(WB_data[32]), .Y(n2330) );
  INVX1 U2097 ( .A(WB_data[32]), .Y(n2331) );
  BUFX2 U2098 ( .A(n2652), .Y(n2332) );
  AND2X1 U2099 ( .A(WB_mult32_result[32]), .B(n2562), .Y(n2651) );
  INVX1 U2100 ( .A(n2651), .Y(n2333) );
  AND2X2 U2101 ( .A(n1994), .B(n2000), .Y(EX_alu_A[0]) );
  INVX1 U2102 ( .A(EX_alu_A[0]), .Y(n2334) );
  AND2X1 U2103 ( .A(instruction[24]), .B(n2557), .Y(n1236) );
  INVX1 U2104 ( .A(n1236), .Y(n2335) );
  INVX1 U2105 ( .A(n1226), .Y(n2336) );
  INVX1 U2106 ( .A(n1224), .Y(n2337) );
  INVX1 U2107 ( .A(n1222), .Y(n2338) );
  INVX1 U2108 ( .A(n1218), .Y(n2339) );
  INVX1 U2109 ( .A(n1211), .Y(n2340) );
  INVX1 U2110 ( .A(n1207), .Y(n2341) );
  INVX1 U2111 ( .A(n1205), .Y(n2342) );
  AND2X1 U2112 ( .A(instruction[9]), .B(n2500), .Y(n1200) );
  INVX1 U2113 ( .A(n1200), .Y(n2343) );
  AND2X1 U2114 ( .A(EX_oprA[7]), .B(n2506), .Y(n3129) );
  INVX1 U2115 ( .A(n3129), .Y(n2344) );
  AND2X1 U2116 ( .A(EX_oprA[29]), .B(n2506), .Y(n3085) );
  INVX1 U2117 ( .A(n3085), .Y(n2345) );
  AND2X1 U2118 ( .A(EX_oprA[44]), .B(n2506), .Y(n3055) );
  INVX1 U2119 ( .A(n3055), .Y(n2346) );
  AND2X1 U2120 ( .A(EX_oprA[59]), .B(n2506), .Y(n3025) );
  INVX1 U2121 ( .A(n3025), .Y(n2347) );
  AND2X1 U2122 ( .A(n2506), .B(EX_dest_reg[1]), .Y(n1193) );
  INVX1 U2123 ( .A(n1193), .Y(n2348) );
  AND2X1 U2124 ( .A(EX_alu_func[2]), .B(n2506), .Y(n1240) );
  INVX1 U2125 ( .A(n1240), .Y(n2349) );
  AND2X1 U2126 ( .A(ID_oprB[55]), .B(n2500), .Y(n3256) );
  INVX1 U2127 ( .A(n3256), .Y(n2350) );
  AND2X1 U2128 ( .A(ID_oprB[43]), .B(n2557), .Y(n3232) );
  INVX1 U2129 ( .A(n3232), .Y(n2351) );
  AND2X1 U2130 ( .A(ID_oprB[32]), .B(n2558), .Y(n3210) );
  INVX1 U2131 ( .A(n3210), .Y(n2352) );
  AND2X1 U2132 ( .A(ID_oprB[17]), .B(n2558), .Y(n3181) );
  INVX1 U2133 ( .A(n3181), .Y(n2353) );
  AND2X1 U2134 ( .A(ID_oprB[4]), .B(n2557), .Y(n3155) );
  INVX1 U2135 ( .A(n3155), .Y(n2354) );
  AND2X1 U2136 ( .A(n1313), .B(ID_instruction[13]), .Y(n1398) );
  INVX1 U2137 ( .A(n1398), .Y(n2355) );
  INVX1 U2138 ( .A(n2668), .Y(n2356) );
  AND2X2 U2139 ( .A(EX_oprB[30]), .B(n2484), .Y(n2658) );
  INVX1 U2140 ( .A(n2658), .Y(n2357) );
  INVX1 U2141 ( .A(n1791), .Y(n2358) );
  AND2X1 U2142 ( .A(instruction[3]), .B(n2554), .Y(n1189) );
  INVX1 U2143 ( .A(n1189), .Y(n2359) );
  INVX1 U2144 ( .A(n2655), .Y(n2360) );
  BUFX2 U2145 ( .A(n1394), .Y(n2361) );
  INVX1 U2146 ( .A(n1405), .Y(n2362) );
  BUFX2 U2147 ( .A(n1406), .Y(n2363) );
  AND2X1 U2148 ( .A(n3128), .B(n3126), .Y(n2998) );
  INVX1 U2149 ( .A(n2998), .Y(n2364) );
  AND2X1 U2150 ( .A(n3124), .B(n3122), .Y(n2999) );
  INVX1 U2151 ( .A(n2999), .Y(n2365) );
  BUFX2 U2152 ( .A(n3000), .Y(n2366) );
  BUFX2 U2153 ( .A(n2941), .Y(n2367) );
  BUFX2 U2154 ( .A(n2824), .Y(n2368) );
  BUFX2 U2155 ( .A(n2894), .Y(n2369) );
  BUFX2 U2156 ( .A(n3012), .Y(n2370) );
  BUFX2 U2157 ( .A(n1359), .Y(n2371) );
  BUFX2 U2158 ( .A(n2960), .Y(n2372) );
  INVX1 U2159 ( .A(WB_data[2]), .Y(n2373) );
  INVX1 U2160 ( .A(WB_data[2]), .Y(n2374) );
  BUFX2 U2161 ( .A(n2731), .Y(n2375) );
  INVX1 U2162 ( .A(n2730), .Y(n2376) );
  AND2X2 U2163 ( .A(n2380), .B(n2379), .Y(WB_data[22]) );
  INVX1 U2164 ( .A(WB_data[22]), .Y(n2377) );
  INVX1 U2165 ( .A(WB_data[22]), .Y(n2378) );
  BUFX2 U2166 ( .A(n2692), .Y(n2379) );
  AND2X1 U2167 ( .A(WB_mult32_result[22]), .B(n2562), .Y(n2691) );
  INVX1 U2168 ( .A(n2691), .Y(n2380) );
  INVX1 U2169 ( .A(n2551), .Y(n2549) );
  AND2X2 U2170 ( .A(EX_oprA[53]), .B(n2534), .Y(n2523) );
  INVX1 U2171 ( .A(n2523), .Y(n2381) );
  AND2X1 U2172 ( .A(instruction[23]), .B(n2500), .Y(n1233) );
  INVX1 U2173 ( .A(n1233), .Y(n2382) );
  INVX1 U2174 ( .A(n1220), .Y(n2383) );
  INVX1 U2175 ( .A(n1209), .Y(n2384) );
  INVX1 U2176 ( .A(n1203), .Y(n2385) );
  AND2X1 U2177 ( .A(instruction[8]), .B(n2500), .Y(n1199) );
  INVX1 U2178 ( .A(n1199), .Y(n2386) );
  AND2X1 U2179 ( .A(EX_oprA[14]), .B(n2506), .Y(n3115) );
  INVX1 U2180 ( .A(n3115), .Y(n2387) );
  AND2X1 U2181 ( .A(EX_oprA[28]), .B(n2506), .Y(n3087) );
  INVX1 U2182 ( .A(n3087), .Y(n2388) );
  AND2X1 U2183 ( .A(EX_oprA[39]), .B(n2506), .Y(n3065) );
  INVX1 U2184 ( .A(n3065), .Y(n2389) );
  AND2X1 U2185 ( .A(EX_oprA[52]), .B(n2506), .Y(n3039) );
  INVX1 U2186 ( .A(n3039), .Y(n2390) );
  AND2X1 U2187 ( .A(EX_oprA[60]), .B(n2506), .Y(n3023) );
  INVX1 U2188 ( .A(n3023), .Y(n2391) );
  AND2X1 U2189 ( .A(n2506), .B(EX_dest_reg[4]), .Y(n1196) );
  INVX1 U2190 ( .A(n1196), .Y(n2392) );
  AND2X1 U2191 ( .A(EX_alu_func[3]), .B(n2506), .Y(n1241) );
  INVX1 U2192 ( .A(n1241), .Y(n2393) );
  AND2X1 U2193 ( .A(ID_oprB[51]), .B(n2500), .Y(n3248) );
  INVX1 U2194 ( .A(n3248), .Y(n2394) );
  AND2X1 U2195 ( .A(ID_oprB[37]), .B(n2557), .Y(n3220) );
  INVX1 U2196 ( .A(n3220), .Y(n2395) );
  AND2X1 U2197 ( .A(ID_oprB[22]), .B(n2557), .Y(n3191) );
  INVX1 U2198 ( .A(n3191), .Y(n2396) );
  AND2X1 U2199 ( .A(ID_oprB[7]), .B(n2558), .Y(n3161) );
  INVX1 U2200 ( .A(n3161), .Y(n2397) );
  AND2X1 U2201 ( .A(ID_oprB[1]), .B(n2557), .Y(n3149) );
  INVX1 U2202 ( .A(n3149), .Y(n2398) );
  AND2X1 U2203 ( .A(n1313), .B(ID_instruction[12]), .Y(n1399) );
  INVX1 U2204 ( .A(n1399), .Y(n2399) );
  BUFX2 U2205 ( .A(n299), .Y(n2400) );
  OR2X1 U2206 ( .A(memAddr[26]), .B(memAddr[28]), .Y(n3278) );
  INVX1 U2207 ( .A(n3278), .Y(n2401) );
  BUFX2 U2208 ( .A(n2947), .Y(n2402) );
  BUFX2 U2209 ( .A(n2945), .Y(n2403) );
  BUFX2 U2210 ( .A(n2820), .Y(n2404) );
  BUFX2 U2211 ( .A(n3010), .Y(n2405) );
  BUFX2 U2212 ( .A(n2885), .Y(n2406) );
  BUFX2 U2213 ( .A(n3271), .Y(n2407) );
  BUFX2 U2214 ( .A(n2657), .Y(n2408) );
  BUFX2 U2215 ( .A(n2952), .Y(n2409) );
  INVX1 U2216 ( .A(WB_data[6]), .Y(n2410) );
  INVX1 U2217 ( .A(WB_data[6]), .Y(n2411) );
  BUFX2 U2218 ( .A(n2719), .Y(n2412) );
  AND2X1 U2219 ( .A(WB_mult32_result[6]), .B(n2562), .Y(n2718) );
  INVX1 U2220 ( .A(n2718), .Y(n2413) );
  BUFX2 U2221 ( .A(n2854), .Y(n2414) );
  AND2X1 U2222 ( .A(instruction[22]), .B(n2558), .Y(n1232) );
  INVX1 U2223 ( .A(n1232), .Y(n2415) );
  AND2X1 U2224 ( .A(instruction[7]), .B(n2500), .Y(n1198) );
  INVX1 U2225 ( .A(n1198), .Y(n2416) );
  AND2X1 U2226 ( .A(EX_oprA[15]), .B(n2506), .Y(n3113) );
  INVX1 U2227 ( .A(n3113), .Y(n2417) );
  AND2X1 U2228 ( .A(EX_oprA[40]), .B(n2506), .Y(n3063) );
  INVX1 U2229 ( .A(n3063), .Y(n2418) );
  AND2X1 U2230 ( .A(EX_oprA[53]), .B(n2506), .Y(n3037) );
  INVX1 U2231 ( .A(n3037), .Y(n2419) );
  AND2X1 U2232 ( .A(EX_oprA[62]), .B(n2506), .Y(n3019) );
  INVX1 U2233 ( .A(n3019), .Y(n2420) );
  AND2X1 U2234 ( .A(EX_shift_amt[4]), .B(n2506), .Y(n1217) );
  INVX1 U2235 ( .A(n1217), .Y(n2421) );
  AND2X1 U2236 ( .A(EX_alu_func[4]), .B(n2506), .Y(n1242) );
  INVX1 U2237 ( .A(n1242), .Y(n2422) );
  AND2X1 U2238 ( .A(ID_oprB[50]), .B(n2500), .Y(n3246) );
  INVX1 U2239 ( .A(n3246), .Y(n2423) );
  AND2X1 U2240 ( .A(ID_oprB[36]), .B(n2557), .Y(n3218) );
  INVX1 U2241 ( .A(n3218), .Y(n2424) );
  AND2X1 U2242 ( .A(ID_oprB[21]), .B(n2558), .Y(n3189) );
  INVX1 U2243 ( .A(n3189), .Y(n2425) );
  AND2X1 U2244 ( .A(ID_oprB[6]), .B(n2558), .Y(n3159) );
  INVX1 U2245 ( .A(n3159), .Y(n2426) );
  AND2X1 U2246 ( .A(ID_oprB[0]), .B(n2500), .Y(n3147) );
  INVX1 U2247 ( .A(n3147), .Y(n2427) );
  AND2X1 U2248 ( .A(n1313), .B(ID_instruction[14]), .Y(n1397) );
  INVX1 U2249 ( .A(n1397), .Y(n2428) );
  BUFX2 U2250 ( .A(n1377), .Y(n2429) );
  AND2X1 U2251 ( .A(n3108), .B(n3106), .Y(n2986) );
  INVX1 U2252 ( .A(n2986), .Y(n2430) );
  INVX1 U2253 ( .A(n2982), .Y(n2431) );
  AND2X1 U2254 ( .A(n3028), .B(n3026), .Y(n2974) );
  INVX1 U2255 ( .A(n2974), .Y(n2432) );
  BUFX2 U2256 ( .A(n2943), .Y(n2433) );
  BUFX2 U2257 ( .A(n2898), .Y(n2434) );
  BUFX2 U2258 ( .A(n2771), .Y(n2435) );
  BUFX2 U2259 ( .A(n3011), .Y(n2436) );
  AND2X2 U2260 ( .A(n2438), .B(n2439), .Y(WB_data[38]) );
  INVX1 U2261 ( .A(WB_data[38]), .Y(n2437) );
  BUFX2 U2262 ( .A(n2634), .Y(n2438) );
  AND2X1 U2263 ( .A(WB_mult32_result[38]), .B(n2562), .Y(n2633) );
  INVX1 U2264 ( .A(n2633), .Y(n2439) );
  BUFX2 U2265 ( .A(n2890), .Y(n2440) );
  BUFX2 U2266 ( .A(n1185), .Y(n2441) );
  BUFX2 U2267 ( .A(n2956), .Y(n2442) );
  AND2X2 U2268 ( .A(n2444), .B(n2445), .Y(WB_data[3]) );
  BUFX2 U2269 ( .A(n2728), .Y(n2444) );
  AND2X1 U2270 ( .A(WB_mult32_result[3]), .B(n2562), .Y(n2727) );
  INVX1 U2271 ( .A(n2727), .Y(n2445) );
  BUFX2 U2272 ( .A(n2855), .Y(n2446) );
  AND2X2 U2273 ( .A(n2508), .B(n2446), .Y(n2509) );
  OR2X1 U2274 ( .A(reset), .B(n3312), .Y(n288) );
  INVX1 U2275 ( .A(n288), .Y(n2447) );
  OR2X1 U2276 ( .A(reset), .B(n3311), .Y(n289) );
  INVX1 U2277 ( .A(n289), .Y(n2448) );
  OR2X1 U2278 ( .A(reset), .B(n2488), .Y(n223) );
  INVX1 U2279 ( .A(n223), .Y(n2449) );
  OR2X1 U2280 ( .A(reset), .B(n3313), .Y(n222) );
  INVX1 U2281 ( .A(n222), .Y(n2450) );
  OR2X1 U2282 ( .A(reset), .B(n3314), .Y(n221) );
  INVX1 U2283 ( .A(n221), .Y(n2451) );
  OR2X1 U2284 ( .A(reset), .B(n3016), .Y(n291) );
  INVX1 U2285 ( .A(n291), .Y(n2452) );
  AND2X1 U2286 ( .A(ID_oprB[26]), .B(n2557), .Y(n3198) );
  INVX1 U2287 ( .A(n3198), .Y(n2453) );
  AND2X1 U2288 ( .A(instruction[15]), .B(n2500), .Y(n1212) );
  INVX1 U2289 ( .A(n1212), .Y(n2454) );
  AND2X1 U2290 ( .A(instruction[6]), .B(n2500), .Y(n1197) );
  INVX1 U2291 ( .A(n1197), .Y(n2455) );
  AND2X1 U2292 ( .A(ID_oprB[62]), .B(n2557), .Y(n3143) );
  INVX1 U2293 ( .A(n3143), .Y(n2456) );
  AND2X1 U2294 ( .A(EX_oprA[16]), .B(n2506), .Y(n3111) );
  INVX1 U2295 ( .A(n3111), .Y(n2457) );
  AND2X1 U2296 ( .A(EX_oprA[41]), .B(n2506), .Y(n3061) );
  INVX1 U2297 ( .A(n3061), .Y(n2458) );
  AND2X1 U2298 ( .A(EX_oprA[56]), .B(n2506), .Y(n3031) );
  INVX1 U2299 ( .A(n3031), .Y(n2459) );
  AND2X1 U2300 ( .A(EX_oprA[61]), .B(n2506), .Y(n3021) );
  INVX1 U2301 ( .A(n3021), .Y(n2460) );
  AND2X1 U2302 ( .A(EX_alu_func[5]), .B(n2506), .Y(n1243) );
  INVX1 U2303 ( .A(n1243), .Y(n2461) );
  AND2X1 U2304 ( .A(EX_oprA[0]), .B(n2506), .Y(n3014) );
  INVX1 U2305 ( .A(n3014), .Y(n2462) );
  OR2X1 U2306 ( .A(n2565), .B(n2785), .Y(n2786) );
  INVX1 U2307 ( .A(n2786), .Y(n2463) );
  OR2X1 U2308 ( .A(dataOut[15]), .B(dataOut[14]), .Y(n2997) );
  INVX1 U2309 ( .A(n2997), .Y(n2464) );
  BUFX2 U2310 ( .A(n1383), .Y(n2465) );
  AND2X1 U2311 ( .A(n3100), .B(n3098), .Y(n2987) );
  INVX1 U2312 ( .A(n2987), .Y(n2466) );
  AND2X1 U2313 ( .A(n3020), .B(n3018), .Y(n2975) );
  INVX1 U2314 ( .A(n2975), .Y(n2467) );
  AND2X1 U2315 ( .A(n3132), .B(n3130), .Y(n2996) );
  INVX1 U2316 ( .A(n2996), .Y(n2468) );
  AND2X2 U2317 ( .A(n2471), .B(n2470), .Y(EX_alu_A[42]) );
  INVX1 U2318 ( .A(EX_alu_A[42]), .Y(n2469) );
  BUFX2 U2319 ( .A(n2833), .Y(n2470) );
  INVX1 U2320 ( .A(n2520), .Y(n2471) );
  BUFX2 U2321 ( .A(n1180), .Y(n2472) );
  AND2X1 U2322 ( .A(n3293), .B(n3280), .Y(n1184) );
  INVX1 U2323 ( .A(n1184), .Y(n2473) );
  BUFX2 U2324 ( .A(n2951), .Y(n2474) );
  BUFX2 U2325 ( .A(n2767), .Y(n2475) );
  BUFX2 U2326 ( .A(n2794), .Y(n2476) );
  AND2X2 U2327 ( .A(n2478), .B(n2479), .Y(WB_data[1]) );
  BUFX2 U2328 ( .A(n2734), .Y(n2478) );
  INVX1 U2329 ( .A(n2733), .Y(n2479) );
  AND2X1 U2330 ( .A(n2503), .B(n2562), .Y(n2605) );
  INVX1 U2331 ( .A(n2605), .Y(n2480) );
  BUFX2 U2332 ( .A(n2962), .Y(n2481) );
  AND2X2 U2333 ( .A(n2489), .B(n2112), .Y(n2923) );
  INVX1 U2334 ( .A(n2923), .Y(n2482) );
  BUFX2 U2335 ( .A(n2877), .Y(n2483) );
  AND2X2 U2336 ( .A(n2514), .B(n2483), .Y(n2507) );
  INVX1 U2337 ( .A(n1202), .Y(n2485) );
  NOR3X1 U2338 ( .A(n2488), .B(PREVIOUS_STALL), .C(n2582), .Y(n2487) );
  INVX1 U2339 ( .A(n1924), .Y(WB_reg_write_load) );
  BUFX2 U2340 ( .A(n1990), .Y(n2489) );
  INVX2 U2341 ( .A(EX_alu_A[11]), .Y(n2571) );
  INVX1 U2342 ( .A(n2607), .Y(n2491) );
  INVX1 U2343 ( .A(n2491), .Y(n2492) );
  INVX1 U2344 ( .A(n2580), .Y(n2495) );
  INVX1 U2345 ( .A(WB_is_load), .Y(n2580) );
  INVX2 U2346 ( .A(EX_alu_A[15]), .Y(n2569) );
  INVX1 U2347 ( .A(n2766), .Y(n2498) );
  AND2X2 U2348 ( .A(n2511), .B(n2105), .Y(n2503) );
  INVX4 U2349 ( .A(n2551), .Y(n2548) );
  AND2X2 U2350 ( .A(n1989), .B(n2747), .Y(n2512) );
  AND2X2 U2351 ( .A(n2511), .B(n2747), .Y(n2513) );
  AND2X2 U2352 ( .A(n2513), .B(n2414), .Y(n2514) );
  AND2X2 U2353 ( .A(n2508), .B(n2483), .Y(n2510) );
  INVX1 U2354 ( .A(n2500), .Y(n2556) );
  INVX1 U2355 ( .A(n2500), .Y(n2555) );
  INVX1 U2356 ( .A(n2506), .Y(n2554) );
  INVX1 U2357 ( .A(n2559), .Y(n2558) );
  INVX1 U2358 ( .A(n2559), .Y(n2557) );
  INVX1 U2359 ( .A(n2500), .Y(n2559) );
  AND2X1 U2360 ( .A(EX_alu_result[61]), .B(n2553), .Y(n226) );
  AND2X1 U2361 ( .A(EX_alu_result[63]), .B(n2553), .Y(n224) );
  AND2X1 U2362 ( .A(EX_alu_result[12]), .B(n2553), .Y(n275) );
  AND2X1 U2363 ( .A(EX_alu_result[14]), .B(n2553), .Y(n273) );
  AND2X1 U2364 ( .A(EX_alu_result[38]), .B(n2553), .Y(n249) );
  AND2X1 U2365 ( .A(EX_alu_result[40]), .B(n2553), .Y(n247) );
  AND2X1 U2366 ( .A(EX_alu_result[42]), .B(n2553), .Y(n245) );
  AND2X1 U2367 ( .A(EX_alu_result[44]), .B(n2553), .Y(n243) );
  AND2X1 U2368 ( .A(EX_alu_result[46]), .B(n2553), .Y(n241) );
  AND2X1 U2369 ( .A(EX_alu_result[6]), .B(n2553), .Y(n281) );
  AND2X1 U2370 ( .A(EX_alu_result[8]), .B(n2553), .Y(n279) );
  AND2X1 U2371 ( .A(EX_alu_result[10]), .B(n2553), .Y(n277) );
  AND2X1 U2372 ( .A(EX_alu_result[2]), .B(n2553), .Y(n285) );
  AND2X1 U2373 ( .A(EX_alu_result[3]), .B(n2553), .Y(n284) );
  AND2X1 U2374 ( .A(EX_alu_result[4]), .B(n2553), .Y(n283) );
  AND2X1 U2375 ( .A(EX_alu_result[5]), .B(n2553), .Y(n282) );
  AND2X1 U2376 ( .A(EX_alu_result[7]), .B(n2553), .Y(n280) );
  AND2X1 U2377 ( .A(EX_alu_result[34]), .B(n2553), .Y(n253) );
  AND2X1 U2378 ( .A(EX_alu_result[35]), .B(n2553), .Y(n252) );
  AND2X1 U2379 ( .A(EX_alu_result[36]), .B(n2553), .Y(n251) );
  AND2X1 U2380 ( .A(EX_alu_result[15]), .B(n2553), .Y(n272) );
  AND2X1 U2381 ( .A(EX_alu_result[31]), .B(n2553), .Y(n256) );
  AND2X1 U2382 ( .A(EX_alu_result[37]), .B(n2553), .Y(n250) );
  AND2X1 U2383 ( .A(EX_alu_result[39]), .B(n2553), .Y(n248) );
  AND2X1 U2384 ( .A(EX_alu_result[41]), .B(n2553), .Y(n246) );
  AND2X1 U2385 ( .A(EX_alu_result[43]), .B(n2553), .Y(n244) );
  AND2X1 U2386 ( .A(EX_alu_result[45]), .B(n2553), .Y(n242) );
  AND2X1 U2387 ( .A(EX_alu_result[47]), .B(n2553), .Y(n240) );
  AND2X1 U2388 ( .A(EX_alu_result[48]), .B(n2553), .Y(n239) );
  AND2X1 U2389 ( .A(EX_alu_result[49]), .B(n2553), .Y(n238) );
  AND2X1 U2390 ( .A(EX_alu_result[50]), .B(n2553), .Y(n237) );
  AND2X1 U2391 ( .A(EX_alu_result[51]), .B(n2553), .Y(n236) );
  AND2X1 U2392 ( .A(EX_alu_result[52]), .B(n2553), .Y(n235) );
  AND2X1 U2393 ( .A(EX_alu_result[53]), .B(n2553), .Y(n234) );
  AND2X1 U2394 ( .A(EX_alu_result[54]), .B(n2553), .Y(n233) );
  AND2X1 U2395 ( .A(EX_alu_result[55]), .B(n2553), .Y(n232) );
  AND2X1 U2396 ( .A(EX_alu_result[56]), .B(n2553), .Y(n231) );
  AND2X1 U2397 ( .A(EX_alu_result[57]), .B(n2553), .Y(n230) );
  AND2X1 U2398 ( .A(EX_alu_result[58]), .B(n2553), .Y(n229) );
  AND2X1 U2399 ( .A(EX_alu_result[59]), .B(n2553), .Y(n228) );
  AND2X1 U2400 ( .A(EX_alu_result[60]), .B(n2553), .Y(n227) );
  AND2X1 U2401 ( .A(EX_alu_result[16]), .B(n2553), .Y(n271) );
  AND2X1 U2402 ( .A(EX_alu_result[17]), .B(n2553), .Y(n270) );
  AND2X1 U2403 ( .A(EX_alu_result[18]), .B(n2553), .Y(n269) );
  AND2X1 U2404 ( .A(EX_alu_result[9]), .B(n2553), .Y(n278) );
  AND2X1 U2405 ( .A(EX_alu_result[11]), .B(n2553), .Y(n276) );
  AND2X1 U2406 ( .A(EX_alu_result[13]), .B(n2553), .Y(n274) );
  AND2X1 U2407 ( .A(EX_alu_result[19]), .B(n2553), .Y(n268) );
  AND2X1 U2408 ( .A(EX_alu_result[20]), .B(n2553), .Y(n267) );
  AND2X1 U2409 ( .A(EX_alu_result[21]), .B(n2553), .Y(n266) );
  AND2X1 U2410 ( .A(EX_alu_result[22]), .B(n2553), .Y(n265) );
  AND2X1 U2411 ( .A(EX_alu_result[23]), .B(n2553), .Y(n264) );
  AND2X1 U2412 ( .A(EX_alu_result[24]), .B(n2553), .Y(n263) );
  AND2X1 U2413 ( .A(EX_alu_result[25]), .B(n2553), .Y(n262) );
  AND2X1 U2414 ( .A(EX_alu_result[26]), .B(n2553), .Y(n261) );
  AND2X1 U2415 ( .A(EX_alu_result[27]), .B(n2553), .Y(n260) );
  AND2X1 U2416 ( .A(EX_alu_result[28]), .B(n2553), .Y(n259) );
  INVX1 U2417 ( .A(dataOut[53]), .Y(n3038) );
  INVX1 U2418 ( .A(dataOut[49]), .Y(n3046) );
  INVX1 U2419 ( .A(dataOut[45]), .Y(n3054) );
  INVX1 U2420 ( .A(dataOut[37]), .Y(n3070) );
  INVX1 U2421 ( .A(dataOut[29]), .Y(n3086) );
  INVX1 U2422 ( .A(dataOut[13]), .Y(n3118) );
  INVX1 U2423 ( .A(dataOut[52]), .Y(n3040) );
  INVX1 U2424 ( .A(dataOut[48]), .Y(n3048) );
  INVX1 U2425 ( .A(dataOut[44]), .Y(n3056) );
  INVX1 U2426 ( .A(dataOut[36]), .Y(n3072) );
  INVX1 U2427 ( .A(dataOut[28]), .Y(n3088) );
  INVX1 U2428 ( .A(dataOut[12]), .Y(n3120) );
  INVX1 U2429 ( .A(dataOut[62]), .Y(n3020) );
  INVX1 U2430 ( .A(dataOut[58]), .Y(n3028) );
  INVX1 U2431 ( .A(dataOut[42]), .Y(n3060) );
  INVX1 U2432 ( .A(dataOut[40]), .Y(n3064) );
  INVX1 U2433 ( .A(dataOut[34]), .Y(n3076) );
  INVX1 U2434 ( .A(dataOut[32]), .Y(n3080) );
  INVX1 U2435 ( .A(dataOut[26]), .Y(n3092) );
  INVX1 U2436 ( .A(dataOut[24]), .Y(n3096) );
  INVX1 U2437 ( .A(dataOut[22]), .Y(n3100) );
  INVX1 U2438 ( .A(dataOut[18]), .Y(n3108) );
  INVX1 U2439 ( .A(dataOut[10]), .Y(n3124) );
  INVX1 U2440 ( .A(dataOut[8]), .Y(n3128) );
  INVX1 U2441 ( .A(dataOut[6]), .Y(n3132) );
  INVX1 U2442 ( .A(dataOut[2]), .Y(n3140) );
  INVX1 U2443 ( .A(dataOut[63]), .Y(n3018) );
  INVX1 U2444 ( .A(dataOut[59]), .Y(n3026) );
  INVX1 U2445 ( .A(dataOut[43]), .Y(n3058) );
  INVX1 U2446 ( .A(dataOut[41]), .Y(n3062) );
  INVX1 U2447 ( .A(dataOut[35]), .Y(n3074) );
  INVX1 U2448 ( .A(dataOut[33]), .Y(n3078) );
  INVX1 U2449 ( .A(dataOut[27]), .Y(n3090) );
  INVX1 U2450 ( .A(dataOut[25]), .Y(n3094) );
  INVX1 U2451 ( .A(dataOut[23]), .Y(n3098) );
  INVX1 U2452 ( .A(dataOut[19]), .Y(n3106) );
  INVX1 U2453 ( .A(dataOut[11]), .Y(n3122) );
  INVX1 U2454 ( .A(dataOut[9]), .Y(n3126) );
  INVX1 U2455 ( .A(dataOut[7]), .Y(n3130) );
  INVX1 U2456 ( .A(dataOut[3]), .Y(n3138) );
  AND2X1 U2457 ( .A(n1919), .B(n2553), .Y(n2500) );
  AND2X1 U2458 ( .A(EX_alu_result[29]), .B(n2553), .Y(n258) );
  AND2X1 U2459 ( .A(n3275), .B(n3276), .Y(n1313) );
  INVX1 U2460 ( .A(n2484), .Y(n2715) );
  AND2X1 U2461 ( .A(n2869), .B(n2562), .Y(n2502) );
  AND2X1 U2462 ( .A(n2511), .B(n2112), .Y(n2504) );
  INVX1 U2463 ( .A(n2545), .Y(n2541) );
  INVX1 U2464 ( .A(n2551), .Y(n2550) );
  INVX1 U2465 ( .A(n2560), .Y(n2564) );
  INVX1 U2466 ( .A(WB_is_mul32), .Y(n2563) );
  INVX1 U2467 ( .A(n2560), .Y(n2565) );
  INVX1 U2468 ( .A(n2510), .Y(n2538) );
  INVX1 U2469 ( .A(n2544), .Y(n2543) );
  AND2X1 U2470 ( .A(EX_alu_result[30]), .B(n2553), .Y(n257) );
  AND2X1 U2471 ( .A(EX_alu_result[62]), .B(n2553), .Y(n225) );
  INVX1 U2472 ( .A(reset), .Y(n2553) );
  INVX1 U2473 ( .A(n2678), .Y(EX_alu_B[26]) );
  INVX1 U2474 ( .A(n1915), .Y(n2716) );
  INVX1 U2475 ( .A(n2610), .Y(n2654) );
  INVX1 U2476 ( .A(WB_mult32_result[7]), .Y(n2924) );
  INVX1 U2477 ( .A(n3282), .Y(n3275) );
  INVX1 U2478 ( .A(n2851), .Y(n2533) );
  INVX1 U2479 ( .A(n2481), .Y(n2683) );
  INVX1 U2480 ( .A(n2442), .Y(n2862) );
  INVX1 U2481 ( .A(n2409), .Y(n2858) );
  INVX1 U2482 ( .A(n2372), .Y(n2865) );
  INVX1 U2483 ( .A(n2301), .Y(n2860) );
  INVX1 U2484 ( .A(n2474), .Y(n2856) );
  INVX1 U2485 ( .A(n2433), .Y(n2752) );
  INVX1 U2486 ( .A(n2402), .Y(n2758) );
  INVX1 U2487 ( .A(n2328), .Y(n2762) );
  INVX1 U2488 ( .A(n2255), .Y(n2811) );
  INVX1 U2489 ( .A(n2515), .Y(n2551) );
  INVX1 U2490 ( .A(n2299), .Y(n2909) );
  INVX1 U2491 ( .A(n2327), .Y(n2903) );
  INVX1 U2492 ( .A(n2368), .Y(n2825) );
  INVX1 U2493 ( .A(n2326), .Y(n2828) );
  INVX1 U2494 ( .A(n2175), .Y(n2906) );
  INVX1 U2495 ( .A(n2256), .Y(n2836) );
  INVX1 U2496 ( .A(n2566), .Y(n2561) );
  INVX1 U2497 ( .A(n2566), .Y(n2560) );
  INVX1 U2498 ( .A(n2566), .Y(n2562) );
  INVX1 U2499 ( .A(n2575), .Y(memAddr[19]) );
  INVX1 U2500 ( .A(n2667), .Y(EX_alu_B[29]) );
  INVX1 U2501 ( .A(n2664), .Y(n2666) );
  INVX1 U2502 ( .A(n2672), .Y(EX_alu_B[28]) );
  INVX1 U2503 ( .A(n2669), .Y(n2671) );
  INVX1 U2504 ( .A(n2662), .Y(EX_alu_B[30]) );
  INVX1 U2505 ( .A(n2659), .Y(n2661) );
  INVX1 U2506 ( .A(n2573), .Y(memAddr[20]) );
  INVX1 U2507 ( .A(n2577), .Y(memAddr[18]) );
  INVX1 U2508 ( .A(EX_alu_A[48]), .Y(n2567) );
  INVX1 U2509 ( .A(n3013), .Y(n3276) );
  INVX1 U2510 ( .A(n2405), .Y(n3273) );
  INVX1 U2511 ( .A(n2436), .Y(n3274) );
  INVX1 U2512 ( .A(n2472), .Y(n3284) );
  INVX1 U2513 ( .A(n2370), .Y(n3283) );
  INVX1 U2514 ( .A(n2190), .Y(n2916) );
  INVX1 U2515 ( .A(WB_mult32_result[57]), .Y(n2606) );
  INVX1 U2516 ( .A(WB_mult32_result[48]), .Y(n2619) );
  INVX1 U2517 ( .A(ID_flush_ff), .Y(n2964) );
  INVX1 U2518 ( .A(memAddr[27]), .Y(n3280) );
  INVX1 U2519 ( .A(n2934), .Y(EX_alu_A[1]) );
  INVX1 U2520 ( .A(n2784), .Y(EX_alu_A[54]) );
  INVX1 U2521 ( .A(n2930), .Y(EX_alu_A[5]) );
  INVX1 U2522 ( .A(n2815), .Y(n2812) );
  INVX1 U2523 ( .A(n2277), .Y(n2807) );
  INVX1 U2524 ( .A(n2237), .Y(n2896) );
  INVX1 U2525 ( .A(n2279), .Y(n2936) );
  INVX1 U2526 ( .A(n2236), .Y(n2832) );
  INVX1 U2527 ( .A(EX_oprB[25]), .Y(n2681) );
  INVX1 U2528 ( .A(n2434), .Y(n2899) );
  INVX1 U2529 ( .A(n2300), .Y(n2817) );
  INVX1 U2530 ( .A(n2761), .Y(n2759) );
  INVX1 U2531 ( .A(n2435), .Y(n2772) );
  INVX1 U2532 ( .A(n2765), .Y(n2763) );
  INVX1 U2533 ( .A(n2276), .Y(n2874) );
  INVX1 U2534 ( .A(n2204), .Y(n2919) );
  INVX1 U2535 ( .A(n2598), .Y(n2596) );
  INVX1 U2536 ( .A(n2257), .Y(n2912) );
  INVX1 U2537 ( .A(n2441), .Y(n3290) );
  INVX1 U2538 ( .A(memAddr[29]), .Y(n3291) );
  INVX1 U2539 ( .A(n2850), .Y(EX_alu_A[33]) );
  INVX1 U2540 ( .A(n2844), .Y(EX_alu_A[39]) );
  INVX1 U2541 ( .A(n2881), .Y(EX_alu_A[22]) );
  INVX1 U2542 ( .A(n2891), .Y(EX_alu_A[17]) );
  INVX1 U2543 ( .A(n2872), .Y(EX_alu_A[25]) );
  INVX1 U2544 ( .A(n2755), .Y(n2753) );
  INVX1 U2545 ( .A(n2595), .Y(n2593) );
  INVX1 U2546 ( .A(n2404), .Y(n2821) );
  INVX1 U2547 ( .A(n2770), .Y(EX_alu_A[57]) );
  INVX1 U2548 ( .A(n2235), .Y(n2840) );
  INVX1 U2549 ( .A(memAddr[28]), .Y(n3292) );
  INVX1 U2550 ( .A(n2933), .Y(EX_alu_A[2]) );
  INVX1 U2551 ( .A(ID_instruction[5]), .Y(n3277) );
  INVX1 U2552 ( .A(WB_PPP[2]), .Y(n2590) );
  INVX1 U2553 ( .A(memAddr[31]), .Y(n3288) );
  INVX1 U2554 ( .A(PREVIOUS_2_STALL), .Y(n2581) );
  INVX1 U2555 ( .A(memAddr[30]), .Y(n3289) );
  INVX1 U2556 ( .A(memAddr[26]), .Y(n3293) );
  INVX1 U2557 ( .A(n2846), .Y(EX_alu_A[37]) );
  INVX1 U2558 ( .A(n2845), .Y(EX_alu_A[38]) );
  INVX1 U2559 ( .A(n2852), .Y(EX_alu_A[32]) );
  INVX1 U2560 ( .A(n3315), .Y(n2577) );
  INVX1 U2561 ( .A(n3317), .Y(n2573) );
  INVX1 U2562 ( .A(n2929), .Y(EX_alu_A[6]) );
  INVX1 U2563 ( .A(n2849), .Y(EX_alu_A[34]) );
  INVX1 U2564 ( .A(memAddr[23]), .Y(n3296) );
  INVX1 U2565 ( .A(memAddr[22]), .Y(n3297) );
  INVX1 U2566 ( .A(n2882), .Y(EX_alu_A[21]) );
  INVX1 U2567 ( .A(memAddr[16]), .Y(n2579) );
  INVX1 U2568 ( .A(n2928), .Y(EX_alu_A[7]) );
  INVX1 U2569 ( .A(n2796), .Y(EX_alu_A[51]) );
  INVX1 U2570 ( .A(n2848), .Y(EX_alu_A[35]) );
  INVX1 U2571 ( .A(n3316), .Y(n2575) );
  INVX1 U2572 ( .A(n2847), .Y(EX_alu_A[36]) );
  INVX1 U2573 ( .A(n2880), .Y(EX_alu_A[23]) );
  INVX1 U2574 ( .A(memAddr[21]), .Y(n3298) );
  INVX1 U2575 ( .A(n2932), .Y(EX_alu_A[3]) );
  INVX1 U2576 ( .A(n2886), .Y(EX_alu_A[19]) );
  INVX1 U2577 ( .A(WB_mult32_result[63]), .Y(n2940) );
  INVX1 U2578 ( .A(WB_mult32_result[62]), .Y(n2942) );
  INVX1 U2579 ( .A(WB_mult32_result[61]), .Y(n2944) );
  INVX1 U2580 ( .A(WB_mult32_result[60]), .Y(n2946) );
  INVX1 U2581 ( .A(WB_mult32_result[59]), .Y(n2948) );
  INVX1 U2582 ( .A(WB_mult32_result[58]), .Y(n2950) );
  INVX1 U2583 ( .A(PREVIOUS_STALL), .Y(n3016) );
  INVX1 U2584 ( .A(n2931), .Y(EX_alu_A[4]) );
  INVX1 U2585 ( .A(ID_instruction[1]), .Y(n3286) );
  INVX1 U2586 ( .A(WB_mult32_result[51]), .Y(n2793) );
  INVX1 U2587 ( .A(EX_oprB[53]), .Y(n3253) );
  INVX1 U2588 ( .A(EX_oprB[13]), .Y(n3174) );
  INVX1 U2589 ( .A(EX_oprB[5]), .Y(n3158) );
  INVX1 U2590 ( .A(EX_oprB[27]), .Y(n3201) );
  INVX1 U2591 ( .A(EX_oprB[55]), .Y(n3257) );
  INVX1 U2592 ( .A(EX_oprB[52]), .Y(n3251) );
  INVX1 U2593 ( .A(EX_oprB[24]), .Y(n3196) );
  INVX1 U2594 ( .A(EX_oprB[20]), .Y(n3188) );
  INVX1 U2595 ( .A(EX_oprB[33]), .Y(n3213) );
  INVX1 U2596 ( .A(EX_oprB[39]), .Y(n3225) );
  INVX1 U2597 ( .A(EX_oprB[50]), .Y(n3247) );
  INVX1 U2598 ( .A(EX_oprB[49]), .Y(n3245) );
  INVX1 U2599 ( .A(EX_oprB[4]), .Y(n3156) );
  INVX1 U2600 ( .A(EX_oprB[1]), .Y(n3150) );
  INVX1 U2601 ( .A(EX_oprB[15]), .Y(n3178) );
  INVX1 U2602 ( .A(EX_oprB[21]), .Y(n3190) );
  INVX1 U2603 ( .A(EX_oprB[37]), .Y(n3221) );
  INVX1 U2604 ( .A(EX_oprB[42]), .Y(n3231) );
  INVX1 U2605 ( .A(EX_oprB[41]), .Y(n3229) );
  INVX1 U2606 ( .A(EX_oprB[47]), .Y(n3241) );
  INVX1 U2607 ( .A(EX_oprB[3]), .Y(n3154) );
  INVX1 U2608 ( .A(EX_oprB[6]), .Y(n3160) );
  INVX1 U2609 ( .A(EX_oprB[7]), .Y(n3162) );
  INVX1 U2610 ( .A(EX_oprB[14]), .Y(n3176) );
  INVX1 U2611 ( .A(EX_oprB[23]), .Y(n3194) );
  INVX1 U2612 ( .A(EX_oprB[22]), .Y(n3192) );
  INVX1 U2613 ( .A(EX_oprB[35]), .Y(n3217) );
  INVX1 U2614 ( .A(EX_oprB[38]), .Y(n3223) );
  INVX1 U2615 ( .A(EX_oprB[43]), .Y(n3233) );
  INVX1 U2616 ( .A(EX_oprB[46]), .Y(n3239) );
  INVX1 U2617 ( .A(EX_oprB[8]), .Y(n3164) );
  INVX1 U2618 ( .A(EX_oprB[10]), .Y(n3168) );
  INVX1 U2619 ( .A(EX_oprB[32]), .Y(n3211) );
  INVX1 U2620 ( .A(EX_oprB[40]), .Y(n3227) );
  INVX1 U2621 ( .A(WB_mult32_result[56]), .Y(n2774) );
  INVX1 U2622 ( .A(EX_oprB[56]), .Y(n3259) );
  INVX1 U2623 ( .A(EX_oprB[0]), .Y(n3148) );
  INVX1 U2624 ( .A(EX_oprB[12]), .Y(n3172) );
  INVX1 U2625 ( .A(EX_oprB[16]), .Y(n3180) );
  INVX1 U2626 ( .A(EX_oprB[19]), .Y(n3186) );
  INVX1 U2627 ( .A(EX_oprB[45]), .Y(n3237) );
  INVX1 U2628 ( .A(EX_oprB[48]), .Y(n3243) );
  INVX1 U2629 ( .A(EX_oprB[51]), .Y(n3249) );
  INVX1 U2630 ( .A(EX_oprB[2]), .Y(n3152) );
  INVX1 U2631 ( .A(EX_oprB[9]), .Y(n3166) );
  INVX1 U2632 ( .A(EX_oprB[11]), .Y(n3170) );
  INVX1 U2633 ( .A(EX_oprB[18]), .Y(n3184) );
  INVX1 U2634 ( .A(EX_oprB[34]), .Y(n3215) );
  INVX1 U2635 ( .A(EX_oprB[36]), .Y(n3219) );
  INVX1 U2636 ( .A(EX_oprB[44]), .Y(n3235) );
  INVX1 U2637 ( .A(EX_oprB[17]), .Y(n3182) );
  INVX1 U2638 ( .A(EX_oprB[54]), .Y(n3255) );
  INVX1 U2639 ( .A(EX_oprB[57]), .Y(n3261) );
  INVX1 U2640 ( .A(ID_instruction[3]), .Y(n3287) );
  INVX1 U2641 ( .A(WB_mult32_result[49]), .Y(n2801) );
  INVX1 U2642 ( .A(ID_instruction[2]), .Y(n3310) );
  INVX1 U2643 ( .A(dataOut[61]), .Y(n3022) );
  INVX1 U2644 ( .A(dataOut[60]), .Y(n3024) );
  INVX1 U2645 ( .A(dataOut[57]), .Y(n3030) );
  INVX1 U2646 ( .A(dataOut[55]), .Y(n3034) );
  INVX1 U2647 ( .A(dataOut[54]), .Y(n3036) );
  INVX1 U2648 ( .A(EX_oprB[62]), .Y(n3144) );
  INVX1 U2649 ( .A(EX_oprB[63]), .Y(n3146) );
  INVX1 U2650 ( .A(EX_oprB[26]), .Y(n3199) );
  INVX1 U2651 ( .A(EX_oprB[28]), .Y(n3203) );
  INVX1 U2652 ( .A(EX_oprB[29]), .Y(n3205) );
  INVX1 U2653 ( .A(EX_oprB[30]), .Y(n3207) );
  INVX1 U2654 ( .A(EX_oprB[31]), .Y(n3209) );
  INVX1 U2655 ( .A(EX_oprB[58]), .Y(n3263) );
  INVX1 U2656 ( .A(EX_oprB[59]), .Y(n3265) );
  INVX1 U2657 ( .A(EX_oprB[60]), .Y(n3267) );
  INVX1 U2658 ( .A(EX_oprB[61]), .Y(n3269) );
  INVX1 U2659 ( .A(dataOut[0]), .Y(n3015) );
  INVX1 U2660 ( .A(dataOut[56]), .Y(n3032) );
  INVX1 U2661 ( .A(dataOut[51]), .Y(n3042) );
  INVX1 U2662 ( .A(dataOut[50]), .Y(n3044) );
  INVX1 U2663 ( .A(dataOut[47]), .Y(n3050) );
  INVX1 U2664 ( .A(dataOut[46]), .Y(n3052) );
  INVX1 U2665 ( .A(dataOut[39]), .Y(n3066) );
  INVX1 U2666 ( .A(dataOut[38]), .Y(n3068) );
  INVX1 U2667 ( .A(dataOut[31]), .Y(n3082) );
  INVX1 U2668 ( .A(dataOut[30]), .Y(n3084) );
  INVX1 U2669 ( .A(dataOut[21]), .Y(n3102) );
  INVX1 U2670 ( .A(dataOut[20]), .Y(n3104) );
  INVX1 U2671 ( .A(dataOut[17]), .Y(n3110) );
  INVX1 U2672 ( .A(dataOut[16]), .Y(n3112) );
  INVX1 U2673 ( .A(dataOut[15]), .Y(n3114) );
  INVX1 U2674 ( .A(dataOut[14]), .Y(n3116) );
  INVX1 U2675 ( .A(dataOut[5]), .Y(n3134) );
  INVX1 U2676 ( .A(dataOut[4]), .Y(n3136) );
  INVX1 U2677 ( .A(dataOut[1]), .Y(n3142) );
  INVX1 U2678 ( .A(instruction[0]), .Y(n3281) );
  INVX1 U2679 ( .A(ID_instruction[8]), .Y(n3306) );
  INVX1 U2680 ( .A(ID_instruction[12]), .Y(n3302) );
  INVX1 U2681 ( .A(ID_instruction[13]), .Y(n3301) );
  INVX1 U2682 ( .A(EX_dest_reg[1]), .Y(n3314) );
  INVX1 U2683 ( .A(EX_dest_reg[0]), .Y(n3313) );
  INVX1 U2684 ( .A(ID_instruction[15]), .Y(n3299) );
  AND2X1 U2685 ( .A(n1392), .B(n1393), .Y(n2517) );
  INVX1 U2686 ( .A(ID_instruction[6]), .Y(n3308) );
  INVX1 U2687 ( .A(ID_instruction[7]), .Y(n3307) );
  INVX1 U2688 ( .A(ID_instruction[9]), .Y(n3305) );
  INVX1 U2689 ( .A(ID_instruction[10]), .Y(n3304) );
  INVX1 U2690 ( .A(ID_instruction[4]), .Y(n3309) );
  INVX1 U2691 ( .A(n3009), .Y(n3272) );
  AND2X1 U2692 ( .A(n2517), .B(n3309), .Y(n1391) );
  INVX1 U2693 ( .A(EX_is_mul32), .Y(n3311) );
  INVX1 U2694 ( .A(ID_instruction[0]), .Y(n3285) );
  INVX1 U2695 ( .A(ID_instruction[14]), .Y(n3300) );
  INVX1 U2696 ( .A(ID_instruction[11]), .Y(n3303) );
  INVX1 U2697 ( .A(memAddr[25]), .Y(n3294) );
  INVX1 U2698 ( .A(memAddr[24]), .Y(n3295) );
  AND2X1 U2699 ( .A(n2553), .B(EX_dest_reg[3]), .Y(n219) );
  AND2X1 U2700 ( .A(n2553), .B(EX_dest_reg[4]), .Y(n218) );
  AND2X1 U2701 ( .A(n2553), .B(EX_dest_reg[2]), .Y(n220) );
  INVX1 U2702 ( .A(EX_is_load), .Y(n3312) );
  AND2X1 U2703 ( .A(n2553), .B(EX_PPP[2]), .Y(n215) );
  AND2X1 U2704 ( .A(n2553), .B(EX_PPP[1]), .Y(n216) );
  AND2X1 U2705 ( .A(n2553), .B(EX_PPP[0]), .Y(n217) );
  BUFX2 U2706 ( .A(n2437), .Y(n2519) );
  INVX1 U2707 ( .A(WB_mult32_result[53]), .Y(n2785) );
  AND2X2 U2708 ( .A(n1992), .B(n2381), .Y(n2787) );
  INVX1 U2709 ( .A(WB_mult32_result[54]), .Y(n2612) );
  INVX1 U2710 ( .A(WB_mult32_result[40]), .Y(n2842) );
  INVX1 U2711 ( .A(WB_mult32_result[46]), .Y(n2819) );
  INVX1 U2712 ( .A(WB_mult32_result[9]), .Y(n2524) );
  INVX1 U2713 ( .A(WB_mult32_result[44]), .Y(n2525) );
  INVX1 U2714 ( .A(WB_mult32_result[50]), .Y(n2797) );
  INVX1 U2715 ( .A(n1923), .Y(n2957) );
  INVX1 U2716 ( .A(WB_mult32_result[52]), .Y(n2789) );
  INVX1 U2717 ( .A(WB_mult32_result[55]), .Y(n2776) );
  INVX1 U2718 ( .A(WB_mult32_result[42]), .Y(n2834) );
  INVX1 U2719 ( .A(WB_mult32_result[47]), .Y(n2814) );
  INVX1 U2720 ( .A(WB_mult32_result[41]), .Y(n2838) );
  INVX1 U2721 ( .A(WB_mult32_result[45]), .Y(n2823) );
  INVX1 U2722 ( .A(WB_mult32_result[43]), .Y(n2830) );
  AOI22X1 U2723 ( .A(dataIn[63]), .B(n2548), .C(WB_alu_result[63]), .D(n2541), 
        .Y(n2939) );
  XOR2X1 U2724 ( .A(WB_dest_reg[2]), .B(EX_regB[2]), .Y(n2584) );
  XOR2X1 U2725 ( .A(WB_dest_reg[4]), .B(EX_regB[4]), .Y(n2583) );
  OAI21X1 U2726 ( .A(WB_reg_write), .B(WB_is_load), .C(n2581), .Y(n2582) );
  NOR3X1 U2727 ( .A(n2584), .B(n2583), .C(n2741), .Y(n2589) );
  XOR2X1 U2728 ( .A(WB_dest_reg[0]), .B(EX_regB[0]), .Y(n2587) );
  XOR2X1 U2729 ( .A(WB_dest_reg[3]), .B(EX_regB[3]), .Y(n2586) );
  XOR2X1 U2730 ( .A(WB_dest_reg[1]), .B(EX_regB[1]), .Y(n2585) );
  NOR3X1 U2731 ( .A(n2587), .B(n2586), .C(n2585), .Y(n2588) );
  NAND3X1 U2732 ( .A(WB_PPP[1]), .B(n2590), .C(n2592), .Y(n2854) );
  NAND3X1 U2733 ( .A(WB_PPP[0]), .B(n2590), .C(n2591), .Y(n2877) );
  NAND3X1 U2734 ( .A(n2590), .B(n2592), .C(n2591), .Y(n2689) );
  NAND3X1 U2735 ( .A(n2414), .B(n2483), .C(n2131), .Y(n2746) );
  OAI21X1 U2736 ( .A(n2561), .B(n2748), .C(n2503), .Y(n2595) );
  OAI21X1 U2737 ( .A(WB_PPP[1]), .B(n2486), .C(WB_PPP[0]), .Y(n2747) );
  NAND3X1 U2738 ( .A(WB_PPP[1]), .B(n2486), .C(n2592), .Y(n2855) );
  NAND3X1 U2739 ( .A(n2486), .B(n2592), .C(n2591), .Y(n2777) );
  NAND3X1 U2740 ( .A(n2513), .B(n2446), .C(n2132), .Y(n2607) );
  AOI22X1 U2741 ( .A(EX_oprB[63]), .B(n2493), .C(n2593), .D(n2748), .Y(n2594)
         );
  OAI21X1 U2742 ( .A(n2940), .B(n2595), .C(n2002), .Y(EX_alu_B[63]) );
  AOI22X1 U2743 ( .A(dataIn[62]), .B(n2546), .C(WB_alu_result[62]), .D(n2497), 
        .Y(n2941) );
  OAI21X1 U2744 ( .A(n2561), .B(n2750), .C(n2503), .Y(n2598) );
  AOI22X1 U2745 ( .A(EX_oprB[62]), .B(n2493), .C(n2596), .D(n2750), .Y(n2597)
         );
  OAI21X1 U2746 ( .A(n2942), .B(n2598), .C(n2003), .Y(EX_alu_B[62]) );
  AOI22X1 U2747 ( .A(dataIn[61]), .B(n2546), .C(WB_alu_result[61]), .D(n2516), 
        .Y(n2943) );
  AOI22X1 U2748 ( .A(EX_oprB[61]), .B(n2493), .C(n2503), .D(n2752), .Y(n2599)
         );
  OAI21X1 U2749 ( .A(n2944), .B(n2480), .C(n2005), .Y(EX_alu_B[61]) );
  AOI22X1 U2750 ( .A(dataIn[60]), .B(n2546), .C(WB_alu_result[60]), .D(n2516), 
        .Y(n2945) );
  OAI21X1 U2751 ( .A(WB_is_mul32), .B(n2756), .C(n2503), .Y(n2602) );
  AOI22X1 U2752 ( .A(EX_oprB[60]), .B(n2493), .C(n2600), .D(n2756), .Y(n2601)
         );
  OAI21X1 U2753 ( .A(n2946), .B(n2602), .C(n2007), .Y(EX_alu_B[60]) );
  AOI22X1 U2754 ( .A(dataIn[59]), .B(n2546), .C(WB_alu_result[59]), .D(n2542), 
        .Y(n2947) );
  AOI22X1 U2755 ( .A(n2503), .B(n2758), .C(EX_oprB[59]), .D(n2493), .Y(n2603)
         );
  OAI21X1 U2756 ( .A(n2948), .B(n2480), .C(n2008), .Y(EX_alu_B[59]) );
  AOI22X1 U2757 ( .A(dataIn[58]), .B(n2546), .C(WB_alu_result[58]), .D(n2516), 
        .Y(n2949) );
  AOI22X1 U2758 ( .A(n2503), .B(n2762), .C(EX_oprB[58]), .D(n2493), .Y(n2604)
         );
  OAI21X1 U2759 ( .A(n2950), .B(n2480), .C(n2009), .Y(EX_alu_B[58]) );
  AOI22X1 U2760 ( .A(dataIn[57]), .B(n2546), .C(WB_alu_result[57]), .D(n2516), 
        .Y(n2767) );
  OAI21X1 U2761 ( .A(n2565), .B(n2606), .C(n2475), .Y(WB_data[57]) );
  OAI21X1 U2762 ( .A(n2629), .B(n3261), .C(n2042), .Y(EX_alu_B[57]) );
  AOI22X1 U2763 ( .A(dataIn[56]), .B(n2546), .C(WB_alu_result[56]), .D(n2542), 
        .Y(n2771) );
  OAI21X1 U2764 ( .A(n2565), .B(n2774), .C(n2435), .Y(WB_data[56]) );
  OAI21X1 U2765 ( .A(n2629), .B(n3259), .C(n2043), .Y(EX_alu_B[56]) );
  AOI22X1 U2766 ( .A(dataIn[55]), .B(n2546), .C(WB_alu_result[55]), .D(n2496), 
        .Y(n2780) );
  OAI21X1 U2767 ( .A(n2565), .B(n2776), .C(n2118), .Y(WB_data[55]) );
  NAND3X1 U2768 ( .A(n2513), .B(n2483), .C(n2132), .Y(n2610) );
  NAND3X1 U2769 ( .A(n2414), .B(n2131), .C(n2446), .Y(n2775) );
  OAI21X1 U2770 ( .A(n2654), .B(n3257), .C(n1971), .Y(EX_alu_B[55]) );
  AOI22X1 U2771 ( .A(dataIn[54]), .B(n2546), .C(WB_alu_result[54]), .D(n2543), 
        .Y(n2781) );
  OAI21X1 U2772 ( .A(n2565), .B(n2612), .C(n2127), .Y(WB_data[54]) );
  OAI21X1 U2773 ( .A(n2654), .B(n3255), .C(n2044), .Y(EX_alu_B[54]) );
  AOI22X1 U2774 ( .A(dataIn[53]), .B(n2546), .C(WB_alu_result[53]), .D(n2539), 
        .Y(n2788) );
  OAI21X1 U2775 ( .A(n2564), .B(n2785), .C(n1993), .Y(WB_data[53]) );
  OAI21X1 U2776 ( .A(n2654), .B(n3253), .C(n2045), .Y(EX_alu_B[53]) );
  AOI22X1 U2777 ( .A(dataIn[52]), .B(n2546), .C(WB_alu_result[52]), .D(n2134), 
        .Y(n2792) );
  OAI21X1 U2778 ( .A(n2564), .B(n2789), .C(n2120), .Y(WB_data[52]) );
  OAI21X1 U2779 ( .A(n2654), .B(n3251), .C(n2046), .Y(EX_alu_B[52]) );
  AOI22X1 U2780 ( .A(dataIn[51]), .B(n2547), .C(WB_alu_result[51]), .D(n2539), 
        .Y(n2794) );
  OAI21X1 U2781 ( .A(n2565), .B(n2793), .C(n2476), .Y(WB_data[51]) );
  OAI21X1 U2782 ( .A(n2654), .B(n3249), .C(n1972), .Y(EX_alu_B[51]) );
  AOI22X1 U2783 ( .A(dataIn[50]), .B(n2547), .C(WB_alu_result[50]), .D(n2496), 
        .Y(n2800) );
  OAI21X1 U2784 ( .A(n2564), .B(n2797), .C(n2122), .Y(WB_data[50]) );
  OAI21X1 U2785 ( .A(n2654), .B(n3247), .C(n1942), .Y(EX_alu_B[50]) );
  AOI22X1 U2786 ( .A(dataIn[49]), .B(n2547), .C(WB_alu_result[49]), .D(n2539), 
        .Y(n2805) );
  OAI21X1 U2787 ( .A(n2565), .B(n2801), .C(n2124), .Y(WB_data[49]) );
  OAI21X1 U2788 ( .A(n2654), .B(n3245), .C(n1943), .Y(EX_alu_B[49]) );
  AOI22X1 U2789 ( .A(dataIn[48]), .B(n2547), .C(WB_alu_result[48]), .D(n2539), 
        .Y(n2806) );
  OAI21X1 U2790 ( .A(n2565), .B(n2619), .C(n2277), .Y(WB_data[48]) );
  OAI21X1 U2791 ( .A(n2654), .B(n3243), .C(n1944), .Y(EX_alu_B[48]) );
  AOI22X1 U2792 ( .A(dataIn[47]), .B(n2547), .C(WB_alu_result[47]), .D(n2543), 
        .Y(n2810) );
  OAI21X1 U2793 ( .A(n2564), .B(n2814), .C(n2255), .Y(WB_data[47]) );
  OAI21X1 U2794 ( .A(n2629), .B(n3241), .C(n2047), .Y(EX_alu_B[47]) );
  AOI22X1 U2795 ( .A(dataIn[46]), .B(n2547), .C(WB_alu_result[46]), .D(n2542), 
        .Y(n2816) );
  OAI21X1 U2796 ( .A(n2564), .B(n2819), .C(n2300), .Y(WB_data[46]) );
  OAI21X1 U2797 ( .A(n2629), .B(n3239), .C(n2048), .Y(EX_alu_B[46]) );
  AOI22X1 U2798 ( .A(dataIn[45]), .B(n2547), .C(WB_alu_result[45]), .D(n2134), 
        .Y(n2820) );
  OAI21X1 U2799 ( .A(n2564), .B(n2823), .C(n2404), .Y(WB_data[45]) );
  OAI21X1 U2800 ( .A(n2629), .B(n3237), .C(n2049), .Y(EX_alu_B[45]) );
  AOI22X1 U2801 ( .A(dataIn[44]), .B(n2547), .C(WB_alu_result[44]), .D(n2516), 
        .Y(n2824) );
  OAI21X1 U2802 ( .A(n2564), .B(n2525), .C(n2368), .Y(WB_data[44]) );
  OAI21X1 U2803 ( .A(n2629), .B(n3235), .C(n2050), .Y(EX_alu_B[44]) );
  AOI22X1 U2804 ( .A(dataIn[43]), .B(n2547), .C(WB_alu_result[43]), .D(n2542), 
        .Y(n2827) );
  OAI21X1 U2805 ( .A(n2564), .B(n2830), .C(n2326), .Y(WB_data[43]) );
  OAI21X1 U2806 ( .A(n2629), .B(n3233), .C(n1945), .Y(EX_alu_B[43]) );
  AOI22X1 U2807 ( .A(dataIn[42]), .B(n2547), .C(WB_alu_result[42]), .D(n2543), 
        .Y(n2831) );
  OAI21X1 U2808 ( .A(n2564), .B(n2834), .C(n2236), .Y(WB_data[42]) );
  OAI21X1 U2809 ( .A(n2629), .B(n3231), .C(n2051), .Y(EX_alu_B[42]) );
  AOI22X1 U2810 ( .A(dataIn[41]), .B(n2547), .C(WB_alu_result[41]), .D(n2540), 
        .Y(n2835) );
  OAI21X1 U2811 ( .A(n2564), .B(n2838), .C(n2256), .Y(WB_data[41]) );
  OAI21X1 U2812 ( .A(n2629), .B(n3229), .C(n1973), .Y(EX_alu_B[41]) );
  AOI22X1 U2813 ( .A(dataIn[40]), .B(n2547), .C(WB_alu_result[40]), .D(n2539), 
        .Y(n2839) );
  OAI21X1 U2814 ( .A(n2564), .B(n2842), .C(n2235), .Y(WB_data[40]) );
  OAI21X1 U2815 ( .A(n2629), .B(n3227), .C(n1946), .Y(EX_alu_B[40]) );
  AOI22X1 U2816 ( .A(WB_alu_result[39]), .B(n2540), .C(dataIn[39]), .D(n2546), 
        .Y(n2631) );
  OAI21X1 U2817 ( .A(n2654), .B(n3225), .C(n2052), .Y(EX_alu_B[39]) );
  AOI22X1 U2818 ( .A(dataIn[38]), .B(n2547), .C(WB_alu_result[38]), .D(n2539), 
        .Y(n2634) );
  OAI21X1 U2819 ( .A(n2654), .B(n3223), .C(n2053), .Y(EX_alu_B[38]) );
  AOI22X1 U2820 ( .A(dataIn[37]), .B(n2548), .C(WB_alu_result[37]), .D(n2540), 
        .Y(n2637) );
  OAI21X1 U2821 ( .A(n2654), .B(n3221), .C(n2054), .Y(EX_alu_B[37]) );
  AOI22X1 U2822 ( .A(dataIn[36]), .B(n2548), .C(WB_alu_result[36]), .D(n2539), 
        .Y(n2640) );
  OAI21X1 U2823 ( .A(n2654), .B(n3219), .C(n2055), .Y(EX_alu_B[36]) );
  AOI22X1 U2824 ( .A(dataIn[35]), .B(n2548), .C(WB_alu_result[35]), .D(n2134), 
        .Y(n2643) );
  OAI21X1 U2825 ( .A(n2654), .B(n3217), .C(n2056), .Y(EX_alu_B[35]) );
  AOI22X1 U2826 ( .A(dataIn[34]), .B(n2548), .C(WB_alu_result[34]), .D(n2540), 
        .Y(n2646) );
  OAI21X1 U2827 ( .A(n2654), .B(n3215), .C(n2057), .Y(EX_alu_B[34]) );
  AOI22X1 U2828 ( .A(dataIn[33]), .B(n2548), .C(WB_alu_result[33]), .D(n2134), 
        .Y(n2649) );
  OAI21X1 U2829 ( .A(n2654), .B(n3213), .C(n2058), .Y(EX_alu_B[33]) );
  AOI22X1 U2830 ( .A(dataIn[32]), .B(n2548), .C(WB_alu_result[32]), .D(n2540), 
        .Y(n2652) );
  OAI21X1 U2831 ( .A(n2654), .B(n3211), .C(n1947), .Y(EX_alu_B[32]) );
  AOI22X1 U2832 ( .A(dataIn[31]), .B(n2548), .C(WB_alu_result[31]), .D(n2516), 
        .Y(n2951) );
  NAND3X1 U2833 ( .A(n2483), .B(n2131), .C(n2132), .Y(n2853) );
  OAI21X1 U2834 ( .A(n2561), .B(n2856), .C(n1991), .Y(n2656) );
  AOI21X1 U2835 ( .A(EX_oprB[31]), .B(n2484), .C(n2360), .Y(n2657) );
  AOI22X1 U2836 ( .A(n2408), .B(n2529), .C(n2408), .D(n2656), .Y(n3271) );
  AOI22X1 U2837 ( .A(dataIn[30]), .B(n2548), .C(WB_alu_result[30]), .D(n2540), 
        .Y(n2952) );
  OAI21X1 U2838 ( .A(n2561), .B(n2858), .C(n2684), .Y(n2659) );
  OAI21X1 U2839 ( .A(n2409), .B(n2659), .C(n2357), .Y(n2660) );
  AOI21X1 U2840 ( .A(n2661), .B(WB_mult32_result[30]), .C(n2660), .Y(n2662) );
  AOI22X1 U2841 ( .A(dataIn[29]), .B(n2548), .C(WB_alu_result[29]), .D(n2516), 
        .Y(n2954) );
  OAI21X1 U2842 ( .A(n2561), .B(n2860), .C(n2684), .Y(n2664) );
  OAI21X1 U2843 ( .A(n2301), .B(n2664), .C(n2059), .Y(n2665) );
  AOI21X1 U2844 ( .A(n2666), .B(n1926), .C(n2665), .Y(n2667) );
  AOI22X1 U2845 ( .A(dataIn[28]), .B(n2548), .C(WB_alu_result[28]), .D(n2497), 
        .Y(n2956) );
  OAI21X1 U2846 ( .A(n2561), .B(n2862), .C(n2684), .Y(n2669) );
  OAI21X1 U2847 ( .A(n2442), .B(n2669), .C(n2356), .Y(n2670) );
  AOI21X1 U2848 ( .A(n2671), .B(n1923), .C(n2670), .Y(n2672) );
  AOI22X1 U2849 ( .A(dataIn[27]), .B(n2548), .C(WB_alu_result[27]), .D(n2516), 
        .Y(n2958) );
  AOI21X1 U2850 ( .A(n2126), .B(n2565), .C(n2129), .Y(n2673) );
  OAI21X1 U2851 ( .A(n1930), .B(n2125), .C(n2036), .Y(n2674) );
  OAI21X1 U2852 ( .A(n2715), .B(n3201), .C(n2674), .Y(EX_alu_B[27]) );
  AOI22X1 U2853 ( .A(dataIn[26]), .B(n2548), .C(WB_alu_result[26]), .D(n2134), 
        .Y(n2960) );
  OAI21X1 U2854 ( .A(n2372), .B(n2129), .C(n2060), .Y(n2676) );
  AOI21X1 U2855 ( .A(n2677), .B(n2684), .C(n2676), .Y(n2678) );
  AOI22X1 U2856 ( .A(dataIn[25]), .B(n2549), .C(WB_alu_result[25]), .D(n2496), 
        .Y(n2962) );
  NAND3X1 U2857 ( .A(n2684), .B(WB_is_mul32), .C(WB_mult32_result[25]), .Y(
        n2680) );
  OAI21X1 U2858 ( .A(n2715), .B(n2681), .C(n2037), .Y(n2682) );
  AOI22X1 U2859 ( .A(dataIn[24]), .B(n2549), .C(WB_alu_result[24]), .D(n2540), 
        .Y(n2873) );
  OAI21X1 U2860 ( .A(n2564), .B(n2876), .C(n2276), .Y(WB_data[24]) );
  OAI21X1 U2861 ( .A(n2715), .B(n3196), .C(n1948), .Y(EX_alu_B[24]) );
  AOI22X1 U2862 ( .A(dataIn[23]), .B(n2549), .C(WB_alu_result[23]), .D(n2496), 
        .Y(n2688) );
  NAND3X1 U2863 ( .A(n2446), .B(n2131), .C(n2132), .Y(n2878) );
  OAI21X1 U2864 ( .A(n2507), .B(n3194), .C(n2061), .Y(EX_alu_B[23]) );
  AOI22X1 U2865 ( .A(dataIn[22]), .B(n2549), .C(WB_alu_result[22]), .D(n2540), 
        .Y(n2692) );
  OAI21X1 U2866 ( .A(n2507), .B(n3192), .C(n1974), .Y(EX_alu_B[22]) );
  AOI22X1 U2867 ( .A(dataIn[21]), .B(n2549), .C(WB_alu_result[21]), .D(n2496), 
        .Y(n2695) );
  OAI21X1 U2868 ( .A(n2507), .B(n3190), .C(n1975), .Y(EX_alu_B[21]) );
  AOI22X1 U2869 ( .A(dataIn[20]), .B(n2549), .C(WB_alu_result[20]), .D(n2496), 
        .Y(n2885) );
  OAI21X1 U2870 ( .A(n2564), .B(n2883), .C(n2406), .Y(WB_data[20]) );
  OAI21X1 U2871 ( .A(n2507), .B(n3188), .C(n1949), .Y(EX_alu_B[20]) );
  AOI22X1 U2872 ( .A(dataIn[19]), .B(n2549), .C(WB_alu_result[19]), .D(n2496), 
        .Y(n2699) );
  OAI21X1 U2873 ( .A(n2507), .B(n3186), .C(n1976), .Y(EX_alu_B[19]) );
  AOI22X1 U2874 ( .A(dataIn[18]), .B(n2549), .C(WB_alu_result[18]), .D(n2496), 
        .Y(n2890) );
  OAI21X1 U2875 ( .A(n2563), .B(n2887), .C(n2440), .Y(WB_data[18]) );
  OAI21X1 U2876 ( .A(n2507), .B(n3184), .C(n2062), .Y(EX_alu_B[18]) );
  AOI22X1 U2877 ( .A(dataIn[17]), .B(n2549), .C(WB_alu_result[17]), .D(n2496), 
        .Y(n2703) );
  OAI21X1 U2878 ( .A(n2507), .B(n3182), .C(n1977), .Y(EX_alu_B[17]) );
  AOI22X1 U2879 ( .A(dataIn[16]), .B(n2549), .C(WB_alu_result[16]), .D(n2496), 
        .Y(n2894) );
  OAI21X1 U2880 ( .A(n2563), .B(n2705), .C(n2369), .Y(WB_data[16]) );
  OAI21X1 U2881 ( .A(n2507), .B(n3180), .C(n1950), .Y(EX_alu_B[16]) );
  AOI22X1 U2882 ( .A(dataIn[15]), .B(n2549), .C(WB_alu_result[15]), .D(n2496), 
        .Y(n2895) );
  OAI21X1 U2883 ( .A(n2563), .B(n2526), .C(n2237), .Y(WB_data[15]) );
  OAI21X1 U2884 ( .A(n2715), .B(n3178), .C(n1978), .Y(EX_alu_B[15]) );
  AOI22X1 U2885 ( .A(dataIn[14]), .B(n2549), .C(WB_alu_result[14]), .D(n2539), 
        .Y(n2898) );
  OAI21X1 U2886 ( .A(n2563), .B(n2901), .C(n2434), .Y(WB_data[14]) );
  OAI21X1 U2887 ( .A(n2715), .B(n3176), .C(n1951), .Y(EX_alu_B[14]) );
  AOI22X1 U2888 ( .A(dataIn[13]), .B(n2549), .C(WB_alu_result[13]), .D(n2496), 
        .Y(n2902) );
  OAI21X1 U2889 ( .A(n2563), .B(n2521), .C(n2327), .Y(WB_data[13]) );
  OAI21X1 U2890 ( .A(n2715), .B(n3174), .C(n1952), .Y(EX_alu_B[13]) );
  AOI22X1 U2891 ( .A(dataIn[12]), .B(n2550), .C(WB_alu_result[12]), .D(n2496), 
        .Y(n2905) );
  OAI21X1 U2892 ( .A(n2563), .B(n2528), .C(n2175), .Y(WB_data[12]) );
  OAI21X1 U2893 ( .A(n2715), .B(n3172), .C(n2063), .Y(EX_alu_B[12]) );
  AOI22X1 U2894 ( .A(dataIn[11]), .B(n2550), .C(WB_alu_result[11]), .D(n2496), 
        .Y(n2908) );
  OAI21X1 U2895 ( .A(n2563), .B(n2530), .C(n2299), .Y(WB_data[11]) );
  OAI21X1 U2896 ( .A(n2715), .B(n3170), .C(n1979), .Y(EX_alu_B[11]) );
  AOI22X1 U2897 ( .A(dataIn[10]), .B(n2550), .C(WB_alu_result[10]), .D(n2134), 
        .Y(n2911) );
  OAI21X1 U2898 ( .A(n2563), .B(n2914), .C(n2257), .Y(WB_data[10]) );
  OAI21X1 U2899 ( .A(n2715), .B(n3168), .C(n2064), .Y(EX_alu_B[10]) );
  AOI22X1 U2900 ( .A(dataIn[9]), .B(n2550), .C(WB_alu_result[9]), .D(n2496), 
        .Y(n2915) );
  OAI21X1 U2901 ( .A(n2563), .B(n2524), .C(n2190), .Y(WB_data[9]) );
  OAI21X1 U2902 ( .A(n2715), .B(n3166), .C(n2065), .Y(EX_alu_B[9]) );
  AOI22X1 U2903 ( .A(dataIn[8]), .B(n2550), .C(WB_alu_result[8]), .D(n2496), 
        .Y(n2918) );
  OAI21X1 U2904 ( .A(n2563), .B(n2921), .C(n2204), .Y(WB_data[8]) );
  OAI21X1 U2905 ( .A(n2715), .B(n3164), .C(n2066), .Y(EX_alu_B[8]) );
  AOI22X1 U2906 ( .A(dataIn[7]), .B(n2550), .C(WB_alu_result[7]), .D(n2542), 
        .Y(n2925) );
  OAI21X1 U2907 ( .A(n2563), .B(n2716), .C(n2329), .Y(WB_data[7]) );
  OAI21X1 U2908 ( .A(n2507), .B(n3162), .C(n2067), .Y(EX_alu_B[7]) );
  AOI22X1 U2909 ( .A(dataIn[6]), .B(n2550), .C(WB_alu_result[6]), .D(n2496), 
        .Y(n2719) );
  OAI21X1 U2910 ( .A(n2507), .B(n3160), .C(n1980), .Y(EX_alu_B[6]) );
  AOI22X1 U2911 ( .A(dataIn[5]), .B(n2550), .C(WB_alu_result[5]), .D(n2496), 
        .Y(n2722) );
  OAI21X1 U2912 ( .A(n2507), .B(n3158), .C(n1981), .Y(EX_alu_B[5]) );
  AOI22X1 U2913 ( .A(dataIn[4]), .B(n2550), .C(WB_alu_result[4]), .D(n2496), 
        .Y(n2725) );
  OAI21X1 U2914 ( .A(n2507), .B(n3156), .C(n1982), .Y(EX_alu_B[4]) );
  AOI22X1 U2915 ( .A(dataIn[3]), .B(n2550), .C(WB_alu_result[3]), .D(n2496), 
        .Y(n2728) );
  OAI21X1 U2916 ( .A(n2507), .B(n3154), .C(n1983), .Y(EX_alu_B[3]) );
  AOI22X1 U2917 ( .A(dataIn[2]), .B(n2550), .C(WB_alu_result[2]), .D(n2496), 
        .Y(n2731) );
  OAI21X1 U2918 ( .A(n2507), .B(n3152), .C(n1984), .Y(EX_alu_B[2]) );
  AOI22X1 U2919 ( .A(dataIn[1]), .B(n2550), .C(WB_alu_result[1]), .D(n2134), 
        .Y(n2734) );
  OAI21X1 U2920 ( .A(n2507), .B(n3150), .C(n2068), .Y(EX_alu_B[1]) );
  AOI22X1 U2921 ( .A(dataIn[0]), .B(n2546), .C(WB_alu_result[0]), .D(n2496), 
        .Y(n2935) );
  OAI21X1 U2922 ( .A(n2563), .B(n2736), .C(n2279), .Y(WB_data[0]) );
  OAI21X1 U2923 ( .A(n2507), .B(n3148), .C(n1985), .Y(EX_alu_B[0]) );
  XNOR2X1 U2924 ( .A(EX_regA[3]), .B(WB_dest_reg[3]), .Y(n2740) );
  XNOR2X1 U2925 ( .A(EX_regA[1]), .B(WB_dest_reg[1]), .Y(n2739) );
  XNOR2X1 U2926 ( .A(EX_regA[0]), .B(WB_dest_reg[0]), .Y(n2738) );
  NAND3X1 U2927 ( .A(n2740), .B(n2739), .C(n2738), .Y(n2745) );
  XNOR2X1 U2928 ( .A(WB_dest_reg[4]), .B(EX_regA[4]), .Y(n2743) );
  XNOR2X1 U2929 ( .A(WB_dest_reg[2]), .B(EX_regA[2]), .Y(n2742) );
  NAND3X1 U2930 ( .A(n2743), .B(n2742), .C(n2487), .Y(n2744) );
  AOI22X1 U2931 ( .A(n2499), .B(n2748), .C(EX_oprA[63]), .D(n2532), .Y(n2749)
         );
  OAI21X1 U2932 ( .A(n2940), .B(n2843), .C(n2011), .Y(EX_alu_A[63]) );
  AOI22X1 U2933 ( .A(EX_oprA[62]), .B(n2532), .C(n2499), .D(n2750), .Y(n2751)
         );
  OAI21X1 U2934 ( .A(n2942), .B(n2843), .C(n1958), .Y(EX_alu_A[62]) );
  OAI21X1 U2935 ( .A(n2561), .B(n2752), .C(n2499), .Y(n2755) );
  AOI22X1 U2936 ( .A(EX_oprA[61]), .B(n2532), .C(n2753), .D(n2752), .Y(n2754)
         );
  OAI21X1 U2937 ( .A(n2944), .B(n2755), .C(n1959), .Y(EX_alu_A[61]) );
  AOI22X1 U2938 ( .A(n2499), .B(n2756), .C(EX_oprA[60]), .D(n2532), .Y(n2757)
         );
  OAI21X1 U2939 ( .A(n2946), .B(n2843), .C(n2320), .Y(EX_alu_A[60]) );
  OAI21X1 U2940 ( .A(n2561), .B(n2758), .C(n2499), .Y(n2761) );
  AOI22X1 U2941 ( .A(EX_oprA[59]), .B(n2532), .C(n2759), .D(n2758), .Y(n2760)
         );
  OAI21X1 U2942 ( .A(n2948), .B(n2761), .C(n1960), .Y(EX_alu_A[59]) );
  OAI21X1 U2943 ( .A(n2561), .B(n2762), .C(n2499), .Y(n2765) );
  AOI22X1 U2944 ( .A(EX_oprA[58]), .B(n2532), .C(n2763), .D(n2762), .Y(n2764)
         );
  OAI21X1 U2945 ( .A(n2950), .B(n2765), .C(n1961), .Y(EX_alu_A[58]) );
  AOI21X1 U2946 ( .A(n2475), .B(n2565), .C(n2498), .Y(n2769) );
  AOI22X1 U2947 ( .A(n1925), .B(EX_oprA[57]), .C(n2078), .D(n2081), .Y(n2770)
         );
  AOI22X1 U2948 ( .A(EX_oprA[56]), .B(n2532), .C(n1929), .D(n2772), .Y(n2773)
         );
  OAI21X1 U2949 ( .A(n2843), .B(n2774), .C(n2012), .Y(EX_alu_A[56]) );
  NAND3X1 U2950 ( .A(n2132), .B(n2483), .C(n2512), .Y(n2851) );
  AOI22X1 U2951 ( .A(n2135), .B(n1939), .C(EX_oprA[55]), .D(n2534), .Y(n2779)
         );
  OAI21X1 U2952 ( .A(n2118), .B(n2133), .C(n2013), .Y(EX_alu_A[55]) );
  AOI21X1 U2953 ( .A(n2127), .B(n2565), .C(n2133), .Y(n2783) );
  AOI22X1 U2954 ( .A(n2534), .B(EX_oprA[54]), .C(n1987), .D(n1954), .Y(n2784)
         );
  OAI21X1 U2955 ( .A(n1993), .B(n2133), .C(n2787), .Y(EX_alu_A[53]) );
  AOI22X1 U2956 ( .A(n1940), .B(n2135), .C(EX_oprA[52]), .D(n2534), .Y(n2791)
         );
  OAI21X1 U2957 ( .A(n2120), .B(n2133), .C(n1962), .Y(EX_alu_A[52]) );
  AOI22X1 U2958 ( .A(n2476), .B(n2563), .C(n2476), .D(n2793), .Y(n2795) );
  AOI22X1 U2959 ( .A(EX_oprA[51]), .B(n2534), .C(n2077), .D(n2135), .Y(n2796)
         );
  AOI22X1 U2960 ( .A(n1941), .B(n2135), .C(EX_oprA[50]), .D(n2534), .Y(n2799)
         );
  OAI21X1 U2961 ( .A(n2122), .B(n2133), .C(n2014), .Y(EX_alu_A[50]) );
  AOI22X1 U2962 ( .A(n2075), .B(n2135), .C(EX_oprA[49]), .D(n2534), .Y(n2803)
         );
  OAI21X1 U2963 ( .A(n2124), .B(n2133), .C(n2016), .Y(EX_alu_A[49]) );
  NAND3X1 U2964 ( .A(WB_is_mul32), .B(n2135), .C(WB_mult32_result[48]), .Y(
        n2809) );
  AOI22X1 U2965 ( .A(EX_oprA[48]), .B(n2534), .C(n2135), .D(n2807), .Y(n2808)
         );
  OAI21X1 U2966 ( .A(n2561), .B(n2811), .C(n1929), .Y(n2815) );
  AOI22X1 U2967 ( .A(n2812), .B(n2811), .C(EX_oprA[47]), .D(n1925), .Y(n2813)
         );
  OAI21X1 U2968 ( .A(n2815), .B(n2814), .C(n1963), .Y(EX_alu_A[47]) );
  AOI22X1 U2969 ( .A(EX_oprA[46]), .B(n2532), .C(n2499), .D(n2817), .Y(n2818)
         );
  OAI21X1 U2970 ( .A(n2843), .B(n2819), .C(n2018), .Y(EX_alu_A[46]) );
  AOI22X1 U2971 ( .A(EX_oprA[45]), .B(n1925), .C(n1929), .D(n2821), .Y(n2822)
         );
  OAI21X1 U2972 ( .A(n2843), .B(n2823), .C(n1964), .Y(EX_alu_A[45]) );
  AOI22X1 U2973 ( .A(n1929), .B(n2825), .C(EX_oprA[44]), .D(n2532), .Y(n2826)
         );
  OAI21X1 U2974 ( .A(n2843), .B(n2525), .C(n1965), .Y(EX_alu_A[44]) );
  AOI22X1 U2975 ( .A(n1929), .B(n2828), .C(EX_oprA[43]), .D(n1925), .Y(n2829)
         );
  OAI21X1 U2976 ( .A(n2843), .B(n2830), .C(n1966), .Y(EX_alu_A[43]) );
  AOI22X1 U2977 ( .A(EX_oprA[42]), .B(n2532), .C(n2499), .D(n2832), .Y(n2833)
         );
  AOI22X1 U2978 ( .A(n1929), .B(n2836), .C(EX_oprA[41]), .D(n1925), .Y(n2837)
         );
  OAI21X1 U2979 ( .A(n2843), .B(n2838), .C(n1967), .Y(EX_alu_A[41]) );
  AOI22X1 U2980 ( .A(n2499), .B(n2840), .C(EX_oprA[40]), .D(n1925), .Y(n2841)
         );
  OAI21X1 U2981 ( .A(n2843), .B(n2842), .C(n1968), .Y(EX_alu_A[40]) );
  AOI22X1 U2982 ( .A(EX_oprA[39]), .B(n2534), .C(n2135), .D(n2149), .Y(n2844)
         );
  AOI22X1 U2983 ( .A(EX_oprA[38]), .B(n2534), .C(n2135), .D(n2437), .Y(n2845)
         );
  AOI22X1 U2984 ( .A(EX_oprA[37]), .B(n2534), .C(n2135), .D(n2258), .Y(n2846)
         );
  AOI22X1 U2985 ( .A(EX_oprA[36]), .B(n2534), .C(n2135), .D(n2191), .Y(n2847)
         );
  AOI22X1 U2986 ( .A(EX_oprA[35]), .B(n2534), .C(n2135), .D(n2162), .Y(n2848)
         );
  AOI22X1 U2987 ( .A(EX_oprA[34]), .B(n2534), .C(n2135), .D(n2238), .Y(n2849)
         );
  AOI22X1 U2988 ( .A(EX_oprA[33]), .B(n2534), .C(n2135), .D(n2205), .Y(n2850)
         );
  AOI22X1 U2989 ( .A(EX_oprA[32]), .B(n2534), .C(n2135), .D(n2330), .Y(n2852)
         );
  AOI22X1 U2990 ( .A(EX_oprA[31]), .B(n2536), .C(n2490), .D(n2856), .Y(n2857)
         );
  OAI21X1 U2991 ( .A(n2922), .B(n2529), .C(n2019), .Y(EX_alu_A[31]) );
  AOI22X1 U2992 ( .A(EX_oprA[30]), .B(n2536), .C(n2490), .D(n2858), .Y(n2859)
         );
  OAI21X1 U2993 ( .A(n2953), .B(n2922), .C(n1969), .Y(EX_alu_A[30]) );
  AOI22X1 U2994 ( .A(EX_oprA[29]), .B(n1917), .C(n2490), .D(n2860), .Y(n2861)
         );
  OAI21X1 U2995 ( .A(n2922), .B(n2955), .C(n2021), .Y(EX_alu_A[29]) );
  AOI22X1 U2996 ( .A(EX_oprA[28]), .B(n2536), .C(n2108), .D(n2862), .Y(n2863)
         );
  OAI21X1 U2997 ( .A(n2922), .B(n2527), .C(n2022), .Y(EX_alu_A[28]) );
  AOI22X1 U2998 ( .A(EX_oprA[27]), .B(n1917), .C(n2490), .D(n2125), .Y(n2864)
         );
  OAI21X1 U2999 ( .A(n2959), .B(n2922), .C(n2023), .Y(EX_alu_A[27]) );
  OAI21X1 U3000 ( .A(WB_is_mul32), .B(n2865), .C(n2869), .Y(n2868) );
  AOI22X1 U3001 ( .A(EX_oprA[26]), .B(n2536), .C(n2866), .D(n2865), .Y(n2867)
         );
  OAI21X1 U3002 ( .A(n2868), .B(n1932), .C(n2024), .Y(EX_alu_A[26]) );
  AOI21X1 U3003 ( .A(n2481), .B(n2565), .C(n2109), .Y(n2871) );
  AOI22X1 U3004 ( .A(n1917), .B(EX_oprA[25]), .C(n2079), .D(n1988), .Y(n2872)
         );
  AOI22X1 U3005 ( .A(n2490), .B(n2874), .C(EX_oprA[24]), .D(n1917), .Y(n2875)
         );
  OAI21X1 U3006 ( .A(n2922), .B(n2876), .C(n2026), .Y(EX_alu_A[24]) );
  AOI22X1 U3007 ( .A(n2537), .B(EX_oprA[23]), .C(n2494), .D(n1928), .Y(n2880)
         );
  AOI22X1 U3008 ( .A(EX_oprA[22]), .B(n2538), .C(n2494), .D(n2377), .Y(n2881)
         );
  AOI22X1 U3009 ( .A(EX_oprA[21]), .B(n2537), .C(n2494), .D(n1938), .Y(n2882)
         );
  OAI21X1 U3010 ( .A(n2406), .B(n2482), .C(n1922), .Y(EX_alu_A[20]) );
  AOI22X1 U3011 ( .A(EX_oprA[19]), .B(n2538), .C(n2494), .D(n2176), .Y(n2886)
         );
  AOI22X1 U3012 ( .A(n1955), .B(n2494), .C(EX_oprA[18]), .D(n2538), .Y(n2889)
         );
  OAI21X1 U3013 ( .A(n2440), .B(n2482), .C(n1970), .Y(EX_alu_A[18]) );
  AOI22X1 U3014 ( .A(EX_oprA[17]), .B(n2537), .C(n2494), .D(n2302), .Y(n2891)
         );
  AOI22X1 U3015 ( .A(n2275), .B(WB_mult32_result[16]), .C(EX_oprA[16]), .D(
        n2537), .Y(n2893) );
  OAI21X1 U3016 ( .A(n2369), .B(n2482), .C(n2274), .Y(EX_alu_A[16]) );
  AOI22X1 U3017 ( .A(n2490), .B(n2896), .C(EX_oprA[15]), .D(n1917), .Y(n2897)
         );
  OAI21X1 U3018 ( .A(n2922), .B(n2526), .C(n2027), .Y(EX_alu_A[15]) );
  AOI22X1 U3019 ( .A(EX_oprA[14]), .B(n1917), .C(n2490), .D(n2899), .Y(n2900)
         );
  OAI21X1 U3020 ( .A(n2922), .B(n2901), .C(n2029), .Y(EX_alu_A[14]) );
  AOI22X1 U3021 ( .A(EX_oprA[13]), .B(n1917), .C(n2490), .D(n2903), .Y(n2904)
         );
  OAI21X1 U3022 ( .A(n2922), .B(n2521), .C(n2030), .Y(EX_alu_A[13]) );
  AOI22X1 U3023 ( .A(n2490), .B(n2906), .C(EX_oprA[12]), .D(n1917), .Y(n2907)
         );
  OAI21X1 U3024 ( .A(n2922), .B(n2528), .C(n2031), .Y(EX_alu_A[12]) );
  AOI22X1 U3025 ( .A(EX_oprA[11]), .B(n1917), .C(n2490), .D(n2909), .Y(n2910)
         );
  OAI21X1 U3026 ( .A(n2922), .B(n2530), .C(n2032), .Y(EX_alu_A[11]) );
  AOI22X1 U3027 ( .A(EX_oprA[10]), .B(n1917), .C(n2490), .D(n2912), .Y(n2913)
         );
  OAI21X1 U3028 ( .A(n2922), .B(n2914), .C(n2033), .Y(EX_alu_A[10]) );
  AOI22X1 U3029 ( .A(n2490), .B(n2916), .C(EX_oprA[9]), .D(n1917), .Y(n2917)
         );
  OAI21X1 U3030 ( .A(n2922), .B(n2524), .C(n2034), .Y(EX_alu_A[9]) );
  AOI22X1 U3031 ( .A(n2490), .B(n2919), .C(EX_oprA[8]), .D(n1917), .Y(n2920)
         );
  OAI21X1 U3032 ( .A(n2922), .B(n2921), .C(n2035), .Y(EX_alu_A[8]) );
  AOI21X1 U3033 ( .A(n2329), .B(n2565), .C(n2482), .Y(n2927) );
  AOI22X1 U3034 ( .A(EX_oprA[7]), .B(n2538), .C(n2080), .D(n2082), .Y(n2928)
         );
  AOI22X1 U3035 ( .A(EX_oprA[6]), .B(n2537), .C(n2494), .D(n2410), .Y(n2929)
         );
  AOI22X1 U3036 ( .A(EX_oprA[5]), .B(n2538), .C(n2494), .D(n2280), .Y(n2930)
         );
  AOI22X1 U3037 ( .A(EX_oprA[4]), .B(n2537), .C(n2494), .D(n2219), .Y(n2931)
         );
  AOI22X1 U3038 ( .A(EX_oprA[3]), .B(n2538), .C(n2494), .D(n2443), .Y(n2932)
         );
  AOI22X1 U3039 ( .A(EX_oprA[2]), .B(n2537), .C(n2494), .D(n2373), .Y(n2933)
         );
  AOI22X1 U3040 ( .A(EX_oprA[1]), .B(n2538), .C(n2494), .D(n2477), .Y(n2934)
         );
  AOI22X1 U3041 ( .A(n2923), .B(n2936), .C(EX_oprA[0]), .D(n2538), .Y(n2938)
         );
  NAND3X1 U3042 ( .A(n2923), .B(WB_mult32_result[0]), .C(n2560), .Y(n2937) );
  OAI21X1 U3043 ( .A(n2563), .B(n2940), .C(n2278), .Y(WB_data[63]) );
  OAI21X1 U3044 ( .A(n2563), .B(n2942), .C(n2367), .Y(WB_data[62]) );
  OAI21X1 U3045 ( .A(n2563), .B(n2944), .C(n2433), .Y(WB_data[61]) );
  OAI21X1 U3046 ( .A(n2563), .B(n2946), .C(n2403), .Y(WB_data[60]) );
  OAI21X1 U3047 ( .A(n2563), .B(n2948), .C(n2402), .Y(WB_data[59]) );
  OAI21X1 U3048 ( .A(n2563), .B(n2950), .C(n2328), .Y(WB_data[58]) );
  OAI21X1 U3049 ( .A(n2563), .B(n2529), .C(n2474), .Y(WB_data[31]) );
  OAI21X1 U3050 ( .A(n2563), .B(n2953), .C(n2409), .Y(WB_data[30]) );
  OAI21X1 U3051 ( .A(n2563), .B(n2955), .C(n2301), .Y(WB_data[29]) );
  OAI21X1 U3052 ( .A(n2564), .B(n2957), .C(n2442), .Y(WB_data[28]) );
  OAI21X1 U3053 ( .A(n2563), .B(n2959), .C(n2126), .Y(WB_data[27]) );
  OAI21X1 U3054 ( .A(n2563), .B(n2961), .C(n2372), .Y(WB_data[26]) );
  OAI21X1 U3055 ( .A(n2563), .B(n2963), .C(n2481), .Y(WB_data[25]) );
  NOR3X1 U3056 ( .A(n2362), .B(n2095), .C(n2400), .Y(n2965) );
  OAI21X1 U3057 ( .A(n2965), .B(n3013), .C(n2964), .Y(n3282) );
  NAND3X1 U3058 ( .A(ID_instruction[4]), .B(ID_instruction[5]), .C(n2517), .Y(
        n3010) );
  NAND3X1 U3059 ( .A(n2517), .B(ID_instruction[4]), .C(n3277), .Y(n3011) );
  NAND3X1 U3060 ( .A(n3072), .B(n3070), .C(n2083), .Y(n2969) );
  NOR3X1 U3061 ( .A(n2089), .B(n2096), .C(n2101), .Y(n2985) );
  NAND3X1 U3062 ( .A(n3056), .B(n3054), .C(n2084), .Y(n2973) );
  NOR3X1 U3063 ( .A(n2090), .B(n2097), .C(n2102), .Y(n2984) );
  NOR3X1 U3064 ( .A(n2432), .B(dataOut[57]), .C(dataOut[56]), .Y(n2977) );
  NOR3X1 U3065 ( .A(n2467), .B(dataOut[61]), .C(dataOut[60]), .Y(n2976) );
  NAND3X1 U3066 ( .A(n3040), .B(n3038), .C(n2085), .Y(n2981) );
  NAND3X1 U3067 ( .A(n3048), .B(n3046), .C(n2086), .Y(n2980) );
  NOR3X1 U3068 ( .A(n2431), .B(n2093), .C(n2099), .Y(n2983) );
  NAND3X1 U3069 ( .A(n2985), .B(n2984), .C(n2983), .Y(n3006) );
  NOR3X1 U3070 ( .A(n2430), .B(dataOut[17]), .C(dataOut[16]), .Y(n2994) );
  NOR3X1 U3071 ( .A(n2466), .B(dataOut[21]), .C(dataOut[20]), .Y(n2993) );
  NAND3X1 U3072 ( .A(n3088), .B(n3086), .C(n2087), .Y(n2991) );
  NOR3X1 U3073 ( .A(n2092), .B(n2098), .C(n2103), .Y(n2992) );
  NAND3X1 U3074 ( .A(n2994), .B(n2993), .C(n2992), .Y(n3005) );
  NOR3X1 U3075 ( .A(n2324), .B(dataOut[1]), .C(dataOut[0]), .Y(n3003) );
  NOR3X1 U3076 ( .A(n2468), .B(dataOut[5]), .C(dataOut[4]), .Y(n3002) );
  NAND3X1 U3077 ( .A(n3120), .B(n3118), .C(n2464), .Y(n3000) );
  NOR3X1 U3078 ( .A(n2366), .B(n2365), .C(n2364), .Y(n3001) );
  NAND3X1 U3079 ( .A(n3003), .B(n3002), .C(n3001), .Y(n3004) );
  NOR3X1 U3080 ( .A(n2091), .B(n2094), .C(n2100), .Y(n3007) );
  MUX2X1 U3081 ( .B(n2405), .A(n2436), .S(n3007), .Y(n3008) );
  NAND3X1 U3082 ( .A(n2371), .B(n1360), .C(n3016), .Y(n3012) );
  NAND3X1 U3083 ( .A(n1391), .B(ID_instruction[5]), .C(n3275), .Y(n3009) );
  OAI21X1 U3084 ( .A(n2555), .B(n3015), .C(n2462), .Y(n1720) );
  OAI21X1 U3085 ( .A(n2559), .B(n3018), .C(n2267), .Y(n1783) );
  OAI21X1 U3086 ( .A(n2556), .B(n3020), .C(n2420), .Y(n1782) );
  OAI21X1 U3087 ( .A(n2555), .B(n3022), .C(n2460), .Y(n1781) );
  OAI21X1 U3088 ( .A(n2556), .B(n3024), .C(n2391), .Y(n1780) );
  OAI21X1 U3089 ( .A(n2555), .B(n3026), .C(n2347), .Y(n1779) );
  OAI21X1 U3090 ( .A(n2556), .B(n3028), .C(n2311), .Y(n1778) );
  OAI21X1 U3091 ( .A(n2555), .B(n3030), .C(n2289), .Y(n1777) );
  OAI21X1 U3092 ( .A(n2556), .B(n3032), .C(n2459), .Y(n1776) );
  OAI21X1 U3093 ( .A(n2559), .B(n3034), .C(n2266), .Y(n1775) );
  OAI21X1 U3094 ( .A(n2556), .B(n3036), .C(n2248), .Y(n1774) );
  OAI21X1 U3095 ( .A(n2556), .B(n3038), .C(n2419), .Y(n1773) );
  OAI21X1 U3096 ( .A(n2556), .B(n3040), .C(n2390), .Y(n1772) );
  OAI21X1 U3097 ( .A(n2556), .B(n3042), .C(n2228), .Y(n1771) );
  OAI21X1 U3098 ( .A(n2556), .B(n3044), .C(n2214), .Y(n1770) );
  OAI21X1 U3099 ( .A(n2556), .B(n3046), .C(n2200), .Y(n1769) );
  OAI21X1 U3100 ( .A(n2556), .B(n3048), .C(n2186), .Y(n1768) );
  OAI21X1 U3101 ( .A(n2556), .B(n3050), .C(n2171), .Y(n1767) );
  OAI21X1 U3102 ( .A(n2556), .B(n3052), .C(n2158), .Y(n1766) );
  OAI21X1 U3103 ( .A(n2556), .B(n3054), .C(n2145), .Y(n1765) );
  OAI21X1 U3104 ( .A(n2556), .B(n3056), .C(n2346), .Y(n1764) );
  OAI21X1 U3105 ( .A(n2556), .B(n3058), .C(n2310), .Y(n1763) );
  OAI21X1 U3106 ( .A(n2556), .B(n3060), .C(n2288), .Y(n1762) );
  OAI21X1 U3107 ( .A(n2556), .B(n3062), .C(n2458), .Y(n1761) );
  OAI21X1 U3108 ( .A(n2556), .B(n3064), .C(n2418), .Y(n1760) );
  OAI21X1 U3109 ( .A(n2555), .B(n3066), .C(n2389), .Y(n1759) );
  OAI21X1 U3110 ( .A(n2559), .B(n3068), .C(n2265), .Y(n1758) );
  OAI21X1 U3111 ( .A(n2556), .B(n3070), .C(n2247), .Y(n1757) );
  OAI21X1 U3112 ( .A(n2555), .B(n3072), .C(n2227), .Y(n1756) );
  OAI21X1 U3113 ( .A(n2555), .B(n3074), .C(n2213), .Y(n1755) );
  OAI21X1 U3114 ( .A(n2556), .B(n3076), .C(n2199), .Y(n1754) );
  OAI21X1 U3115 ( .A(n2555), .B(n3078), .C(n2185), .Y(n1753) );
  OAI21X1 U3116 ( .A(n2556), .B(n3080), .C(n2170), .Y(n1752) );
  OAI21X1 U3117 ( .A(n2556), .B(n3082), .C(n2157), .Y(n1751) );
  OAI21X1 U3118 ( .A(n2555), .B(n3084), .C(n2144), .Y(n1750) );
  OAI21X1 U3119 ( .A(n2559), .B(n3086), .C(n2345), .Y(n1749) );
  OAI21X1 U3120 ( .A(n2555), .B(n3088), .C(n2388), .Y(n1748) );
  OAI21X1 U3121 ( .A(n2555), .B(n3090), .C(n2309), .Y(n1747) );
  OAI21X1 U3122 ( .A(n2555), .B(n3092), .C(n2287), .Y(n1746) );
  OAI21X1 U3123 ( .A(n2555), .B(n3094), .C(n2264), .Y(n1745) );
  OAI21X1 U3124 ( .A(n2555), .B(n3096), .C(n2246), .Y(n1744) );
  OAI21X1 U3125 ( .A(n2555), .B(n3098), .C(n2226), .Y(n1743) );
  OAI21X1 U3126 ( .A(n2555), .B(n3100), .C(n2212), .Y(n1742) );
  OAI21X1 U3127 ( .A(n2555), .B(n3102), .C(n2198), .Y(n1741) );
  OAI21X1 U3128 ( .A(n2555), .B(n3104), .C(n2184), .Y(n1740) );
  OAI21X1 U3129 ( .A(n2555), .B(n3106), .C(n2169), .Y(n1739) );
  OAI21X1 U3130 ( .A(n2555), .B(n3108), .C(n2156), .Y(n1738) );
  OAI21X1 U3131 ( .A(n2555), .B(n3110), .C(n2143), .Y(n1737) );
  OAI21X1 U3132 ( .A(n2556), .B(n3112), .C(n2457), .Y(n1736) );
  OAI21X1 U3133 ( .A(n2555), .B(n3114), .C(n2417), .Y(n1735) );
  OAI21X1 U3134 ( .A(n2555), .B(n3116), .C(n2387), .Y(n1734) );
  OAI21X1 U3135 ( .A(n2555), .B(n3118), .C(n2308), .Y(n1733) );
  OAI21X1 U3136 ( .A(n2556), .B(n3120), .C(n2286), .Y(n1732) );
  OAI21X1 U3137 ( .A(n2555), .B(n3122), .C(n2263), .Y(n1731) );
  OAI21X1 U3138 ( .A(n2556), .B(n3124), .C(n2245), .Y(n1730) );
  OAI21X1 U3139 ( .A(n2556), .B(n3126), .C(n2225), .Y(n1729) );
  OAI21X1 U3140 ( .A(n2556), .B(n3128), .C(n2211), .Y(n1728) );
  OAI21X1 U3141 ( .A(n2555), .B(n3130), .C(n2344), .Y(n1727) );
  OAI21X1 U3142 ( .A(n2555), .B(n3132), .C(n2197), .Y(n1726) );
  OAI21X1 U3143 ( .A(n2559), .B(n3134), .C(n2183), .Y(n1725) );
  OAI21X1 U3144 ( .A(n2556), .B(n3136), .C(n2168), .Y(n1724) );
  OAI21X1 U3145 ( .A(n2555), .B(n3138), .C(n2155), .Y(n1723) );
  OAI21X1 U3146 ( .A(n2556), .B(n3140), .C(n2142), .Y(n1722) );
  OAI21X1 U3147 ( .A(n2559), .B(n3142), .C(n2137), .Y(n1721) );
  OAI21X1 U3148 ( .A(n2554), .B(n3144), .C(n2456), .Y(n1784) );
  OAI21X1 U3149 ( .A(n1920), .B(n3146), .C(n2244), .Y(n1785) );
  OAI21X1 U3150 ( .A(n2554), .B(n3148), .C(n2427), .Y(n1851) );
  OAI21X1 U3151 ( .A(n1920), .B(n3150), .C(n2398), .Y(n1852) );
  OAI21X1 U3152 ( .A(n2554), .B(n3152), .C(n2295), .Y(n1853) );
  OAI21X1 U3153 ( .A(n1920), .B(n3154), .C(n2273), .Y(n1854) );
  OAI21X1 U3154 ( .A(n2554), .B(n3156), .C(n2354), .Y(n1855) );
  OAI21X1 U3155 ( .A(n1920), .B(n3158), .C(n2318), .Y(n1856) );
  OAI21X1 U3156 ( .A(n2554), .B(n3160), .C(n2426), .Y(n1857) );
  OAI21X1 U3157 ( .A(n1920), .B(n3162), .C(n2397), .Y(n1858) );
  OAI21X1 U3158 ( .A(n2554), .B(n3164), .C(n2294), .Y(n1859) );
  OAI21X1 U3159 ( .A(n1920), .B(n3166), .C(n2272), .Y(n1860) );
  OAI21X1 U3160 ( .A(n2554), .B(n3168), .C(n2254), .Y(n1861) );
  OAI21X1 U3161 ( .A(n1920), .B(n3170), .C(n2234), .Y(n1862) );
  OAI21X1 U3162 ( .A(n2554), .B(n3172), .C(n2218), .Y(n1863) );
  OAI21X1 U3163 ( .A(n1920), .B(n3174), .C(n2203), .Y(n1864) );
  OAI21X1 U3164 ( .A(n2554), .B(n3176), .C(n2189), .Y(n1865) );
  OAI21X1 U3165 ( .A(n1920), .B(n3178), .C(n2174), .Y(n1866) );
  OAI21X1 U3166 ( .A(n2554), .B(n3180), .C(n2161), .Y(n1867) );
  OAI21X1 U3167 ( .A(n2554), .B(n3182), .C(n2353), .Y(n1868) );
  OAI21X1 U3168 ( .A(n1920), .B(n3184), .C(n2317), .Y(n1869) );
  OAI21X1 U3169 ( .A(n2554), .B(n3186), .C(n2148), .Y(n1870) );
  OAI21X1 U3170 ( .A(n1920), .B(n3188), .C(n2138), .Y(n1871) );
  OAI21X1 U3171 ( .A(n2554), .B(n3190), .C(n2425), .Y(n1872) );
  OAI21X1 U3172 ( .A(n1920), .B(n3192), .C(n2396), .Y(n1873) );
  OAI21X1 U3173 ( .A(n2554), .B(n3194), .C(n2293), .Y(n1874) );
  OAI21X1 U3174 ( .A(n1920), .B(n3196), .C(n2271), .Y(n1875) );
  OAI21X1 U3175 ( .A(n2554), .B(n2681), .C(n2194), .Y(n1876) );
  OAI21X1 U3176 ( .A(n1920), .B(n3199), .C(n2453), .Y(n1877) );
  OAI21X1 U3177 ( .A(n2554), .B(n3201), .C(n2253), .Y(n1878) );
  OAI21X1 U3178 ( .A(n1920), .B(n3203), .C(n2181), .Y(n1879) );
  OAI21X1 U3179 ( .A(n2554), .B(n3205), .C(n2166), .Y(n1880) );
  OAI21X1 U3180 ( .A(n2554), .B(n3207), .C(n2153), .Y(n1881) );
  OAI21X1 U3181 ( .A(n1920), .B(n3209), .C(n2140), .Y(n1882) );
  OAI21X1 U3182 ( .A(n2554), .B(n3211), .C(n2352), .Y(n1883) );
  OAI21X1 U3183 ( .A(n1920), .B(n3213), .C(n2316), .Y(n1884) );
  OAI21X1 U3184 ( .A(n2554), .B(n3215), .C(n2233), .Y(n1885) );
  OAI21X1 U3185 ( .A(n1920), .B(n3217), .C(n2217), .Y(n1886) );
  OAI21X1 U3186 ( .A(n2554), .B(n3219), .C(n2424), .Y(n1887) );
  OAI21X1 U3187 ( .A(n1920), .B(n3221), .C(n2395), .Y(n1888) );
  OAI21X1 U3188 ( .A(n2554), .B(n3223), .C(n2292), .Y(n1889) );
  OAI21X1 U3189 ( .A(n1920), .B(n3225), .C(n2270), .Y(n1890) );
  OAI21X1 U3190 ( .A(n2554), .B(n3227), .C(n2252), .Y(n1891) );
  OAI21X1 U3191 ( .A(n1920), .B(n3229), .C(n2202), .Y(n1892) );
  OAI21X1 U3192 ( .A(n2554), .B(n3231), .C(n2188), .Y(n1893) );
  OAI21X1 U3193 ( .A(n1920), .B(n3233), .C(n2351), .Y(n1894) );
  OAI21X1 U3194 ( .A(n1920), .B(n3235), .C(n2315), .Y(n1895) );
  OAI21X1 U3195 ( .A(n1920), .B(n3237), .C(n2232), .Y(n1896) );
  OAI21X1 U3196 ( .A(n1920), .B(n3239), .C(n2216), .Y(n1897) );
  OAI21X1 U3197 ( .A(n2554), .B(n3241), .C(n2173), .Y(n1898) );
  OAI21X1 U3198 ( .A(n1920), .B(n3243), .C(n2160), .Y(n1899) );
  OAI21X1 U3199 ( .A(n2554), .B(n3245), .C(n2147), .Y(n1900) );
  OAI21X1 U3200 ( .A(n1920), .B(n3247), .C(n2423), .Y(n1901) );
  OAI21X1 U3201 ( .A(n2554), .B(n3249), .C(n2394), .Y(n1902) );
  OAI21X1 U3202 ( .A(n1920), .B(n3251), .C(n2291), .Y(n1903) );
  OAI21X1 U3203 ( .A(n2554), .B(n3253), .C(n2269), .Y(n1904) );
  OAI21X1 U3204 ( .A(n1920), .B(n3255), .C(n2251), .Y(n1905) );
  OAI21X1 U3205 ( .A(n2554), .B(n3257), .C(n2350), .Y(n1906) );
  OAI21X1 U3206 ( .A(n1920), .B(n3259), .C(n2314), .Y(n1907) );
  OAI21X1 U3207 ( .A(n2554), .B(n3261), .C(n2231), .Y(n1908) );
  OAI21X1 U3208 ( .A(n1920), .B(n3263), .C(n2180), .Y(n1909) );
  OAI21X1 U3209 ( .A(n2554), .B(n3265), .C(n2165), .Y(n1910) );
  OAI21X1 U3210 ( .A(n1920), .B(n3267), .C(n2152), .Y(n1911) );
  OAI21X1 U3211 ( .A(n2554), .B(n3269), .C(n2139), .Y(n1912) );
  AOI21X1 U3212 ( .A(memAddr[30]), .B(memAddr[31]), .C(memAddr[29]), .Y(n3279)
         );
  AOI22X1 U3213 ( .A(n2074), .B(n2401), .C(n3280), .D(n3293), .Y(n299) );
endmodule

